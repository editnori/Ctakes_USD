CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Dyes|Drug|false|false||Dyenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Contrast Media|Drug|false|false||Contrast Medianull|Contrast Media|Drug|false|false||Contrastnull|Contrast|Modifier|false|false||Contrastnull|Communications Media|Finding|false|false||Media
null|PAMS Media|Finding|false|false||Medianull|Tunica Media|Anatomy|false|false||Media
null|Media layer|Anatomy|false|false||Medianull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|cilostazol|Drug|false|false||cilostazol
null|cilostazol|Drug|false|false||cilostazolnull|varenicline|Drug|false|false||Varenicline
null|varenicline|Drug|false|false||Vareniclinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Melena|Finding|false|false||Melenanull|Dyspnea|Finding|false|false||SOBnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Xarelto|Drug|false|false||Xarelto
null|Xarelto|Drug|false|false||Xareltonull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Hypertensive disease|Disorder|false|false||HTNnull|Pad Dosage Form|Drug|false|false||PADnull|Pad Mass|Disorder|false|false||PAD
null|Peripheral Arterial Diseases|Disorder|false|false||PADnull|PADI4 wt Allele|Finding|false|false||PAD
null|PADI4 gene|Finding|false|false||PAD
null|DHX40 gene|Finding|false|false||PADnull|PAD Regimen|Procedure|false|false||PADnull|Strucure of thick cushion of skin|Anatomy|false|false||PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Laboratory test finding|Lab|false|false||labsnull|Dark color|Modifier|false|false||darknull|Tarry|Finding|false|false||tarrynull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|null|Time|false|false||priornull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|DC Red No. 8|Drug|false|false||bright red
null|DC Red No. 8|Drug|false|false||bright rednull|Bright red color (finding)|Finding|false|false||bright rednull|Above average intellect|Finding|false|false||bright
null|ARID1B wt Allele|Finding|false|false||bright
null|ARID3A gene|Finding|false|false||brightnull|Bright|Modifier|false|false||brightnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Towelettes|Device|false|false||wipingnull|Hemorrhoids|Disorder|false|false||hemorrhoidsnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Benign|Modifier|false|false||benignnull|polyps|Disorder|false|false||polypnull|Internal hemorrhoids|Disorder|false|false||internal hemorrhoidsnull|Code System Type - Internal|Modifier|false|false||internal
null|Internal Surface|Modifier|false|false||internal
null|Internal|Modifier|false|false||internalnull|Hemorrhoids|Disorder|false|false||hemorrhoidsnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Last|Modifier|false|false||lastnull|Regular|Modifier|false|false||regularnull|Current (present time)|Time|false|false||currentlynull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Exertional fatigue|Finding|false|false||exertional fatiguenull|exercise induced|Finding|false|false||exertionalnull|Fatigue|Finding|false|false||fatiguenull|More|LabModifier|false|false||morenull|Dyspnea|Finding|false|false||SOBnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Last|Modifier|false|false||lastnull|6 months|Time|false|false||6 monthsnull|month|Time|false|false||monthsnull|out (of) breath|Finding|false|false||out of breathnull|Breath|Finding|false|false||breathnull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Climbing stairs|Finding|false|false||climbing stairsnull|climbing (history)|Finding|false|false||climbing
null|Climbing|Finding|false|false||climbing
null|Does climb|Finding|false|false||climbingnull|Prior functioning.stairs|Finding|false|false||stairsnull|Dyspnea|Finding|false|false||SOBnull|Prior functioning.stairs|Finding|false|false||stairsnull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Block Dosage Form|Drug|false|false||blocknull|Fixed Block|Finding|false|false||block
null|Obstruction|Finding|false|false||block
null|Blocking|Finding|false|false||blocknull|Geographic Block|Entity|false|false||blocknull|Block (unit of presentation)|LabModifier|false|false||block
null|Block Dosing Unit|LabModifier|false|false||block
null|Block (unit of measure)|LabModifier|false|false||blocknull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Vomiting|Finding|true|false||vomit
null|Vomitus|Finding|true|false||vomitnull|rectal discharge diarrhea (physical finding)|Finding|true|false||diarrhea
null|Diarrhea|Finding|true|false||diarrheanull|Dysuria|Finding|true|false||dysurianull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Unintentional weight loss|Finding|false|false||unintentional weight lossnull|Unintentional|Finding|false|false||unintentionalnull|Weight Loss|Finding|false|false||weight loss
null|Losing Weight (question)|Finding|false|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|false|false||weight lossnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Laboratory test finding|Lab|false|false||Labsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Leukocytes|Anatomy|false|false||WBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Last|Modifier|false|false||Lastnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Basic metabolic panel|Procedure|false|false||Chem 7null|chemical aspects|Finding|false|false||Chemnull|Chemical procedure|Procedure|false|false||Chemnull|Science of Chemistry|Subject|false|false||Chemnull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Nebulizer solution|Drug|false|false||nebsnull|On IV|Finding|false|false||on IVnull|Saline Solution|Drug|false|false||saline
null|Saline Solution|Drug|false|false||salinenull|Saline method|Procedure|false|false||salinenull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Happiness|Finding|false|false||in good spiritsnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|distilled alcoholic beverage|Drug|false|false||spiritsnull|Rectal hemorrhage|Finding|false|false||blood per rectumnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Per rectum|Finding|false|false||per rectum
null|Rectal Route of Administration|Finding|false|false||per rectumnull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false||rectum
null|Rectal Diseases|Disorder|false|false||rectum
null|Benign neoplasm of rectum|Disorder|false|false||rectum
null|Carcinoma in situ of rectum|Disorder|false|false||rectumnull|Procedure on rectum|Procedure|false|false||rectumnull|Pelvis>Rectum|Anatomy|false|false||rectum
null|Rectum|Anatomy|false|false||rectumnull|Undergarment|Device|false|false||underwearnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Asthma|Disorder|false|false||ASTHMAnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Encounter due to tobacco use|Finding|false|false||Tobacco use
null|Tobacco user|Finding|false|false||Tobacco use
null|History of tobacco use|Finding|false|false||Tobacco use
null|Tobacco use|Finding|false|false||Tobacco usenull|null|Attribute|false|false||Tobacco usenull|tobacco leaf allergenic extract|Drug|false|false||Tobacco
null|Tobacco|Drug|false|false||Tobacco
null|Tobacco|Drug|false|false||Tobacco
null|tobacco leaf allergenic extract|Drug|false|false||Tobacconull|Nicotiana tabacum|Entity|false|false||Tobacconull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Peripheral Arterial Diseases|Disorder|false|false||Peripheral Arterial disease
null|Peripheral Vascular Diseases|Disorder|false|false||Peripheral Arterial diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Arteriopathic disease|Disorder|false|false||Arterial diseasenull|Arteries|Anatomy|false|false||Arterialnull|Arterial|Modifier|false|false||Arterialnull|Disease|Disorder|false|false||diseasenull|Recent|Time|false|false||recentnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|iliac stents|Procedure|false|false||iliac stentingnull|Bone structure of ilium|Anatomy|false|false||iliacnull|Stenting|Procedure|false|false||stentingnull|null|Device|false|false||stentingnull|Atrial tachycardia|Disorder|false|false||ATRIAL TACHYCARDIAnull|continuous electrocardiogram atrial tachycardia|Finding|false|false||ATRIAL TACHYCARDIAnull|Heart Atrium|Anatomy|false|false||ATRIALnull|Tachycardia by ECG Finding|Finding|false|false||TACHYCARDIA
null|Tachycardia|Finding|false|false||TACHYCARDIAnull|Atypical chest pain|Finding|false|false||ATYPICAL CHEST PAINnull|atypia morphology|Finding|false|false||ATYPICALnull|Atypical|Modifier|false|false||ATYPICALnull|Chest Pain|Finding|false|false||CHEST PAINnull|null|Attribute|false|false||CHEST PAINnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Cervical radiculitis|Disorder|false|false||CERVICAL RADICULITISnull|Neck|Anatomy|false|false||CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Radiculitis|Disorder|false|false||RADICULITISnull|Cervical spondylosis without myelopathy|Disorder|false|false||CERVICAL SPONDYLOSIS
null|Cervical spondylosis|Disorder|false|false||CERVICAL SPONDYLOSISnull|Neck|Anatomy|false|false||CERVICALnull|Cervical|Modifier|false|false||CERVICALnull|Spondylosis|Disorder|false|false||SPONDYLOSISnull|Coronary artery|Anatomy|false|false||CORONARY ARTERYnull|Heart|Anatomy|false|false||CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Arterial system|Anatomy|false|false||ARTERY
null|Arteries|Anatomy|false|false||ARTERYnull|Disease|Disorder|false|false||DISEASEnull|Headache|Finding|false|false||HEADACHEnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false||HIP REPLACEMENTnull|heme iron polypeptide|Drug|false|false||HIP
null|ST13 protein, human|Drug|false|false||HIP
null|ST13 protein, human|Drug|false|false||HIP
null|RPL29 protein, human|Drug|false|false||HIP
null|RPL29 protein, human|Drug|false|false||HIP
null|HHIP protein, human|Drug|false|false||HIP
null|HHIP protein, human|Drug|false|false||HIP
null|heme iron polypeptide|Drug|false|false||HIPnull|RPL29 wt Allele|Finding|false|false||HIP
null|REG3A gene|Finding|false|false||HIP
null|RPL29 gene|Finding|false|false||HIP
null|ST13 wt Allele|Finding|false|false||HIP
null|ST13 gene|Finding|false|false||HIP
null|HHIP gene|Finding|false|false||HIP
null|HHIP wt Allele|Finding|false|false||HIP
null|REG3A wt Allele|Finding|false|false||HIPnull|Procedure on hip|Procedure|false|false||HIPnull|Lower extremity>Hip|Anatomy|false|false||HIP
null|Hip structure|Anatomy|false|false||HIP
null|Structure of habenulopeduncular tract|Anatomy|false|false||HIP
null|Bone structure of ischium|Anatomy|false|false||HIPnull|Replacement|Finding|false|false||REPLACEMENTnull|Replacement - supply|Procedure|false|false||REPLACEMENT
null|Surgical Replantation|Procedure|false|false||REPLACEMENTnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Herpes zoster (disorder)|Disorder|false|false||HERPES ZOSTER
null|herpesvirus 3, human|Disorder|false|false||HERPES ZOSTERnull|Herpes simplex dermatitis|Disorder|false|false||HERPES
null|null|Disorder|false|false||HERPESnull|Herpes <Hyperinae>|Entity|false|false||HERPESnull|Herpes zoster (disorder)|Disorder|false|false||ZOSTERnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Heart Atrium|Anatomy|false|false||ATRIALnull|Fibrillation|Disorder|false|false||FIBRILLATIONnull|Anxiety Disorders|Disorder|false|false||ANXIETY
null|Anxiety|Disorder|false|false||ANXIETYnull|Anxiety symptoms|Finding|false|false||ANXIETYnull|Gastrointestinal Hemorrhage|Finding|false|false||GASTROINTESTINAL BLEEDINGnull|Gastrointestinal attachment|Finding|false|false||GASTROINTESTINALnull|gastrointestinal|Modifier|false|false||GASTROINTESTINALnull|Hemorrhage|Finding|false|false||BLEEDINGnull|Degenerative polyarthritis|Disorder|false|false||OSTEOARTHRITISnull|Atherosclerosis|Disorder|false|false||ATHEROSCLEROTIC CARDIOVASCULAR DISEASEnull|atherosclerotic|Finding|false|false||ATHEROSCLEROTICnull|Cardiovascular Diseases|Disorder|false|false||CARDIOVASCULAR DISEASEnull|Cardiovascular system|Anatomy|false|false||CARDIOVASCULAR
null|Cardiovascular|Anatomy|false|false||CARDIOVASCULARnull|Peripheral Vascular Diseases|Disorder|false|false||DISEASE, PERIPHERAL VASCULARnull|Disease|Disorder|false|false||DISEASEnull|Peripheral|Modifier|false|false||PERIPHERALnull|Blood Vessel|Anatomy|false|false||VASCULARnull|Vascular|Modifier|false|false||VASCULARnull|Disease|Disorder|false|false||DISEASEnull|reported history of cataract surgery|Finding|false|false||CATARACT SURGERY
null|Consent Type - Cataract Surgery|Finding|false|false||CATARACT SURGERYnull|Cataract surgery|Procedure|false|false||CATARACT SURGERY
null|Cataract Extraction|Procedure|false|false||CATARACT SURGERYnull|Cataract surgery specialty (qualifier value)|Title|false|false||CATARACT SURGERYnull|Cataract|Disorder|false|false||CATARACTnull|cataract on exam (physical finding)|Finding|false|false||CATARACTnull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Bilateral|Modifier|false|false||BILATERALnull|Common iliac artery structure|Anatomy|false|false||COMMON ILIAC ARTERYnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||COMMON
null|shared attribute|Finding|false|false||COMMONnull|Common (qualifier value)|LabModifier|false|false||COMMONnull|Structure of iliac artery|Anatomy|false|false||ILIAC ARTERYnull|Bone structure of ilium|Anatomy|false|false||ILIACnull|Arterial system|Anatomy|false|false||ARTERY
null|Arteries|Anatomy|false|false||ARTERYnull|Stenting|Procedure|false|false||STENTINGnull|null|Device|false|false||STENTINGnull|Silver bunionectomy|Procedure|false|false||BUNIONECTOMYnull|Prosthetic arthroplasty of hip (procedure)|Procedure|false|false||HIP REPLACEMENTnull|heme iron polypeptide|Drug|false|false||HIP
null|ST13 protein, human|Drug|false|false||HIP
null|ST13 protein, human|Drug|false|false||HIP
null|RPL29 protein, human|Drug|false|false||HIP
null|RPL29 protein, human|Drug|false|false||HIP
null|HHIP protein, human|Drug|false|false||HIP
null|HHIP protein, human|Drug|false|false||HIP
null|heme iron polypeptide|Drug|false|false||HIPnull|RPL29 wt Allele|Finding|false|false||HIP
null|REG3A gene|Finding|false|false||HIP
null|RPL29 gene|Finding|false|false||HIP
null|ST13 wt Allele|Finding|false|false||HIP
null|ST13 gene|Finding|false|false||HIP
null|HHIP gene|Finding|false|false||HIP
null|HHIP wt Allele|Finding|false|false||HIP
null|REG3A wt Allele|Finding|false|false||HIPnull|Procedure on hip|Procedure|false|false||HIPnull|Lower extremity>Hip|Anatomy|false|false||HIP
null|Hip structure|Anatomy|false|false||HIP
null|Structure of habenulopeduncular tract|Anatomy|false|false||HIP
null|Bone structure of ischium|Anatomy|false|false||HIPnull|Replacement|Finding|false|false||REPLACEMENTnull|Replacement - supply|Procedure|false|false||REPLACEMENT
null|Surgical Replantation|Procedure|false|false||REPLACEMENTnull|null|Time|false|false||PRIORnull|Cesarean section|Procedure|false|false||CESAREAN SECTIONnull|Cesarean|Procedure|false|false||CESAREANnull|section sample|Drug|false|false||SECTIONnull|Html Link Type - section|Finding|false|false||SECTION
null|Act Class - Section|Finding|false|false||SECTIONnull|Sectioning technique|Procedure|false|false||SECTIONnull|Section - Geographic Area|Entity|false|false||SECTION
null|Section (object)|Entity|false|false||SECTIONnull|Square Mile|LabModifier|false|false||SECTIONnull|Synovial Cyst|Disorder|false|false||GANGLION CYST
null|Myxoid cyst|Disorder|false|false||GANGLION CYSTnull|Synovial Cyst|Disorder|false|false||GANGLION
null|Myxoid cyst|Disorder|false|false||GANGLIONnull|Ganglia|Anatomy|false|false||GANGLIONnull|Cyst|Disorder|false|false||CYSTnull|SpecimenType - Cyst|Finding|false|false||CYST
null|null|Finding|false|false||CYSTnull|Cyst form of protozoa|Entity|false|false||CYSTnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|BORNHOLM EYE DISEASE|Disorder|true|false||bednull|Bachelor of Education|Finding|true|false||bednull|Beds|Device|true|false||bednull|Patient Location - Bed|Modifier|true|false||bednull|Alert brand of caffeine|Drug|true|false||Alert
null|Alert brand of caffeine|Drug|true|false||Alertnull|Mentally alert|Finding|true|false||Alert
null|Consciousness clear|Finding|true|false||Alert
null|Alert note|Finding|true|false||Alert
null|Alert|Finding|true|false||Alertnull|null|Attribute|true|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|true|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|true|false||supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Elevated|Modifier|true|false||elevated
null|High|Modifier|true|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|true|false||LUNGSnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||rales
null|Rales|Finding|true|false||ralesnull|Rhonchi|Finding|true|false||rhonchinull|Irregular|Modifier|false|false||irregularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Systolic Murmurs|Finding|true|false||systolic murmurnull|Systole|Finding|true|false||systolicnull|Heart murmur|Finding|true|false||murmurnull|Pericardial friction rub|Finding|true|false||rubsnull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||ABDnull|ABD (body structure)|Anatomy|true|false||ABD
null|Abdomen|Anatomy|true|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|true|false||bowel soundsnull|Intestines|Anatomy|true|false||bowelnull|null|Device|true|false||soundsnull|null|Phenomenon|true|false||soundsnull|Present|Finding|true|false||present
null|Presentation|Finding|true|false||presentnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Organomegaly|Finding|true|false||organomegalynull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|true|false||Rectum
null|Rectal Diseases|Disorder|true|false||Rectum
null|Benign neoplasm of rectum|Disorder|true|false||Rectum
null|Carcinoma in situ of rectum|Disorder|true|false||Rectumnull|Procedure on rectum|Procedure|true|false||Rectumnull|Pelvis>Rectum|Anatomy|true|false||Rectum
null|Rectum|Anatomy|true|false||Rectumnull|Obvious|Modifier|true|false||obviousnull|Hemorrhoids|Disorder|true|false||hemorrhoidsnull|Hereditary Multiple Exostoses|Disorder|true|false||EXTnull|EXT1 wt Allele|Finding|true|false||EXT
null|EXT1 gene|Finding|true|false||EXTnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|null|Drug|true|false||pulsesnull|Physiologic pulse|Finding|true|false||pulsesnull|Pulse taking|Procedure|true|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gross (qualifier value)|Modifier|true|false||grossnull|Deficit|Modifier|true|false||deficitsnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|true|false||supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Elevated|Modifier|true|false||elevated
null|High|Modifier|true|false||elevatednull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|true|false||LUNGSnull|Wheezing|Finding|false|false||wheezesnull|Respiratory, thoracic and mediastinal disorders|Disorder|true|false||respnull|Respiratory rate|Attribute|true|false||respnull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Irregular|Modifier|false|false||irregularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Systolic Murmurs|Finding|true|false||systolic murmurnull|Systole|Finding|true|false||systolicnull|Heart murmur|Finding|true|false||murmurnull|Pericardial friction rub|Finding|true|false||rubsnull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||ABDnull|ABD (body structure)|Anatomy|true|false||ABD
null|Abdomen|Anatomy|true|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|true|false||bowel soundsnull|Intestines|Anatomy|true|false||bowelnull|null|Device|true|false||soundsnull|null|Phenomenon|true|false||soundsnull|Present|Finding|true|false||present
null|Presentation|Finding|true|false||presentnull|Rebound tenderness|Finding|true|false||rebound tendernessnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Protective muscle spasm|Finding|true|false||guardingnull|Organomegaly|Finding|true|false||organomegalynull|Hereditary Multiple Exostoses|Disorder|true|false||EXTnull|EXT1 wt Allele|Finding|true|false||EXT
null|EXT1 gene|Finding|true|false||EXTnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|null|Drug|true|false||pulsesnull|Physiologic pulse|Finding|true|false||pulsesnull|Pulse taking|Procedure|true|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gross (qualifier value)|Modifier|true|false||grossnull|Deficit|Modifier|true|false||deficitsnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first premolar mesial prosthesis|Device|false|false||28PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first premolar mesial prosthesis|Device|false|false||28PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first premolar mesial prosthesis|Device|false|false||28PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|Esophagogastroduodenoscopy|Procedure|true|false||EGDnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Body Substance Discharge|Finding|true|false||DISCHARGE
null|Discharge Body Fluid|Finding|true|false||DISCHARGE
null|Body Fluid Discharge|Finding|true|false||DISCHARGE
null|null|Finding|true|false||DISCHARGEnull|Patient Discharge|Procedure|true|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|MCOLN1 protein, human|Drug|false|false||Mg-2
null|MCOLN1 protein, human|Drug|false|false||Mg-2null|MCOLN1 wt Allele|Finding|false|false||Mg-2null|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Drops - Drug Form|Drug|false|false||dropnull|Dropping|Event|false|false||dropnull|Drop (unit of presentation)|LabModifier|false|false||drop
null|Drop British|LabModifier|false|false||drop
null|Drop Dosing Unit|LabModifier|false|false||drop
null|Medical Drop|LabModifier|false|false||drop
null|Drop Unit of Volume|LabModifier|false|false||dropnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Progressive|Finding|false|false||progressivenull|Dyspnea|Finding|false|false||SOBnull|Problems - What subject filter|Finding|false|false||PROBLEMSnull|Gastrointestinal Hemorrhage|Finding|false|false||GI Bleednull|Hemorrhage|Finding|false|false||Bleednull|Presentation|Finding|false|false||Presentednull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Melena|Finding|false|false||melenanull|Hematochezia|Disorder|false|false||BRBPRnull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Bore (qualifier value)|LabModifier|false|false||borenull|On IV|Finding|false|false||on IVnull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|rivaroxaban|Drug|false|false||rivaroxaban
null|rivaroxaban|Drug|false|false||rivaroxabannull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Xarelto|Drug|false|false||Xarelto
null|Xarelto|Drug|false|false||Xareltonull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Dyspnea|Finding|false|false||SOBnull|Long Variable|Modifier|false|false||Long
null|Long|Modifier|false|false||Longnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Location characteristic ID - Smoking|Finding|false|false||smoking
null|Smoking|Finding|false|false||smoking
null|Tobacco smoking behavior|Finding|false|false||smokingnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Progressive|Finding|false|false||Progressivenull|Dyspnea on exertion|Finding|false|false||exertional dyspneanull|exercise induced|Finding|false|false||exertionalnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Use of|Finding|false|false||use ofnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Spiriva|Drug|false|false||Spiriva
null|Spiriva|Drug|false|false||Spirivanull|Advair|Drug|false|false||advair
null|Advair|Drug|false|false||advairnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|Nasal Spray brand of phenylephrine|Drug|false|false||nasal spraynull|Nasal spray (device)|Device|false|false||nasal spray
null|Nasal Sprays|Device|false|false||nasal spray
null|Nasal Spray|Device|false|false||nasal spraynull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Spray Dosage Form|Drug|false|false||spraynull|Spray (administration method)|Finding|false|false||spraynull|Spray (action)|Event|false|false||spraynull|Spray Dosing Unit|LabModifier|false|false||spraynull|theophylline|Drug|false|false||theophylline
null|theophylline|Drug|false|false||theophyllinenull|Assay of theophylline|Procedure|false|false||theophyllinenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Science of Etiology|Finding|true|false||Etiology
null|Etiology aspects|Finding|true|false||Etiology
null|Etiology|Finding|true|false||Etiologynull|Communicable Diseases|Disorder|true|false||infectiousnull|infectious - Entity Risk|Modifier|true|false||infectiousnull|Chronicity|Time|true|false||chronicitynull|most likely|Finding|false|false||Most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|bentiromide|Drug|false|false||PFT
null|bentiromide|Drug|false|false||PFTnull|fluorouracil/melphalan/tamoxifen|Procedure|false|false||PFT
null|Pulmonary function tests|Procedure|false|false||PFTnull|area PFt|Anatomy|false|false||PFTnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Location characteristic ID - Smoking|Finding|false|false||Smoking
null|Smoking|Finding|false|false||Smoking
null|Tobacco smoking behavior|Finding|false|false||Smokingnull|Cessation|Event|false|false||cessationnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Problems - What subject filter|Finding|false|false||PROBLEMSnull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|amiodarone|Drug|false|false||amiodarone
null|amiodarone|Drug|false|false||amiodaronenull|Drug assay amiodarone|Procedure|false|false||amiodaronenull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|rivaroxaban|Drug|false|false||rivaroxaban
null|rivaroxaban|Drug|false|false||rivaroxabannull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Hypertensive disease|Disorder|false|false||HTNnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|diltiazem|Drug|false|false||diltiazem
null|diltiazem|Drug|false|false||diltiazemnull|Imdur|Drug|false|false||Imdur
null|Imdur|Drug|false|false||Imdurnull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|Anxiety Disorders|Disorder|false|false||Anxiety
null|Anxiety|Disorder|false|false||Anxietynull|Anxiety symptoms|Finding|false|false||Anxietynull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|lorazepam|Drug|false|false||lorazepam
null|lorazepam|Drug|false|false||lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Dry Eyes brand of ocular lubricant|Drug|false|false||Dry eyesnull|Dry Eye Syndromes|Disorder|false|false||Dry eyes
null|Keratoconjunctivitis Sicca|Disorder|false|false||Dry eyesnull|Dryness of eye|Finding|false|false||Dry eyesnull|Eye|Anatomy|false|false||eyesnull|null|Attribute|false|false||eyesnull|null|Finding|false|false||History of glaucomanull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Glaucoma|Disorder|false|false||glaucomanull|Glaucoma <Glaucomidae>|Entity|false|false||glaucomanull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|latanoprost|Drug|false|false||latanoprost
null|latanoprost|Drug|false|false||latanoprostnull|Eye Drops|Drug|false|false||ophthalmic dropsnull|Ophthalmic Dosage Form|Drug|false|false||ophthalmicnull|Ophthalmic Route of Administration|Finding|false|false||ophthalmicnull|Eye|Anatomy|false|false||ophthalmicnull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|Pad Dosage Form|Drug|false|false||PADnull|Pad Mass|Disorder|false|false||PAD
null|Peripheral Arterial Diseases|Disorder|false|false||PADnull|PADI4 wt Allele|Finding|false|false||PAD
null|PADI4 gene|Finding|false|false||PAD
null|DHX40 gene|Finding|false|false||PADnull|PAD Regimen|Procedure|false|false||PADnull|Strucure of thick cushion of skin|Anatomy|false|false||PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|iliac stents|Procedure|false|false||iliac stentnull|Bone structure of ilium|Anatomy|false|false||iliacnull|null|Device|false|false||stentnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Referral category - Outpatient|Finding|true|false||outpatient
null|Patient Class - Outpatient|Finding|true|false||outpatientnull|Outpatients|Subject|true|false||outpatientnull|Consent Type - Colonoscopy|Procedure|true|false||colonoscopy
null|colonoscopy|Procedure|true|false||colonoscopynull|Source (property) (qualifier value)|Finding|true|false||source
null|Term Source|Finding|true|false||source
null|Source|Finding|true|false||sourcenull|Lower gastrointestinal hemorrhage|Finding|true|false||lower GI Bleednull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Gastrointestinal Hemorrhage|Finding|true|false||GI Bleednull|Hemorrhage|Finding|true|false||Bleednull|Hemoglobin.stable|Finding|false|false||stable hemoglobinnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|Referral category - Inpatient|Finding|true|false||inpatient
null|Patient Class - Inpatient|Finding|true|false||inpatientnull|inpatient encounter|Procedure|true|false||inpatientnull|inpatient|Subject|true|false||inpatientnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Esophagogastroduodenoscopy|Procedure|true|false||EGDnull|Xarelto|Drug|false|false||Xarelto
null|Xarelto|Drug|false|false||Xareltonull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||dailynull|Continuous|Finding|false|false||Continuenull|Encourage smoking cessation|Procedure|false|false||encourage smoking cessationnull|Cessation of smoking|Finding|false|false||smoking cessationnull|Smoking cessation therapy|Procedure|false|false||smoking cessationnull|Cessation|Event|false|false||cessationnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal dosage form|Drug|false|false||NASALnull|Nasal Route of Administration|Finding|false|false||NASAL
null|Nasal (intended site)|Finding|false|false||NASALnull|null|Anatomy|false|false||NASALnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Nasal congestion (finding)|Finding|false|false||nasal congestionnull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Congestion|Finding|false|false||congestionnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false||LEFT EYEnull|Left eye structure|Anatomy|false|false||LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false||LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false||EYE
null|Disorder of eye|Disorder|false|false||EYEnull|Eye - Specimen Source Code|Finding|false|false||EYE
null|Eye problem|Finding|false|false||EYE
null|Eye Specimen|Finding|false|false||EYEnull|Head>Eye|Anatomy|false|false||EYE
null|Eye|Anatomy|false|false||EYE
null|Orbital region|Anatomy|false|false||EYEnull|Once a day, at bedtime|Time|false|false||QHSnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|Theophylline ER|Drug|false|false||Theophylline ER
null|Theophylline ER|Drug|false|false||Theophylline ERnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Preserving|Finding|false|false||Preservnull|Biologic Preservation|Procedure|false|false||Preservnull|Free of (attribute)|Finding|false|false||Freenull|Empty (qualifier)|Modifier|false|false||Freenull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Preserving|Finding|false|false||Preservnull|Biologic Preservation|Procedure|false|false||Preservnull|Free of (attribute)|Finding|false|false||Freenull|Empty (qualifier)|Modifier|false|false||Freenull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|diltiazem|Drug|false|false||Diltiazem
null|diltiazem|Drug|false|false||Diltiazemnull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal brand of oxymetazoline|Drug|false|false||NASAL
null|Nasal dosage form|Drug|false|false||NASALnull|Nasal Route of Administration|Finding|false|false||NASAL
null|Nasal (intended site)|Finding|false|false||NASALnull|null|Anatomy|false|false||NASALnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Nasal congestion (finding)|Finding|false|false||nasal congestionnull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Congestion|Finding|false|false||congestionnull|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskus
null|Fluticasone-Salmeterol Diskus|Drug|false|false||Fluticasone-Salmeterol Diskusnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|Diskus|Device|false|false||Diskusnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazide
null|hydrochlorothiazide|Drug|false|false||Hydrochlorothiazidenull|Daily|Time|false|false||DAILYnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|latanoprost|Drug|false|false||Latanoprost
null|latanoprost|Drug|false|false||Latanoprostnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|examination of left eye|Procedure|false|false||LEFT EYEnull|Left eye structure|Anatomy|false|false||LEFT EYEnull|Table Cell Horizontal Align - left|Finding|false|false||LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Carcinoma in situ of eye|Disorder|false|false||EYE
null|Disorder of eye|Disorder|false|false||EYEnull|Eye - Specimen Source Code|Finding|false|false||EYE
null|Eye problem|Finding|false|false||EYE
null|Eye Specimen|Finding|false|false||EYEnull|Head>Eye|Anatomy|false|false||EYE
null|Eye|Anatomy|false|false||EYE
null|Orbital region|Anatomy|false|false||EYEnull|Once a day, at bedtime|Time|false|false||QHSnull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|rivaroxaban|Drug|false|false||Rivaroxaban
null|rivaroxaban|Drug|false|false||Rivaroxabannull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Theophylline ER|Drug|false|false||Theophylline ER
null|Theophylline ER|Drug|false|false||Theophylline ERnull|theophylline|Drug|false|false||Theophylline
null|theophylline|Drug|false|false||Theophyllinenull|Assay of theophylline|Procedure|false|false||Theophyllinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|tiotropium bromide|Drug|false|false||Tiotropium Bromide
null|tiotropium bromide|Drug|false|false||Tiotropium Bromidenull|tiotropium|Drug|false|false||Tiotropium
null|tiotropium|Drug|false|false||Tiotropiumnull|Bromides|Drug|false|false||Bromidenull|Bromides measurement|Procedure|false|false||Bromidenull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Minerals|Drug|false|false||mineralsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Reduced|Finding|false|false||decreasenull|Decrease|LabModifier|false|false||decreasenull|In Blood|Finding|false|false||in bloodnull|Blood Cell Count|Procedure|false|false||blood countnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Laboratory Procedures|Procedure|false|false||laboratory testingnull|Diagnostic Service Section ID - Laboratory|Finding|false|false||laboratory
null|Laboratory domain|Finding|false|false||laboratory
null|Referral type - Laboratory|Finding|false|false||laboratorynull|null|Attribute|false|false||laboratorynull|Laboratory|Device|false|false||laboratorynull|Laboratory observation|Lab|false|false||laboratorynull|Laboratory|Entity|false|false||laboratorynull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|Hemorrhage|Finding|false|false||bleednull|Gastrointestinal tract structure|Anatomy|false|false||GI tractnull|Tract|Anatomy|false|false||tractnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Endoscopy, Gastrointestinal|Procedure|false|false||endoscopy
null|Endoscopy (procedure)|Procedure|false|false||endoscopynull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|counts|LabModifier|false|false||countsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Future|Time|false|false||futurenull|Diagnostic Service Section ID - Pulmonary Function|Finding|false|false||Pulmonary function
null|Pulmonary function|Finding|false|false||Pulmonary function
null|Pulmonary function (finding)|Finding|false|false||Pulmonary functionnull|Pulmonary (intended site)|Finding|false|false||Pulmonarynull|Lung|Anatomy|false|false||Pulmonarynull|null|Attribute|false|false||Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|In care (finding)|Finding|true|false||care
null|Continuity Assessment Record and Evaluation|Finding|true|false||carenull|care activity|Event|true|false||carenull|Referral category - Inpatient|Finding|false|false||Inpatient
null|Patient Class - Inpatient|Finding|false|false||Inpatientnull|inpatient encounter|Procedure|false|false||Inpatientnull|inpatient|Subject|false|false||Inpatientnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions