CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|INJECTION, MEROPENEM, 100 MG ADMINISTERED|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenem
null|meropenem|Drug|false|false||meropenemnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Hematochezia|Disorder|false|false||BRBPRnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|aborted - QueryStatusCode|Finding|false|false||aborted
null|aborted - ActStatus|Finding|false|false||aborted
null|Order aborted|Finding|false|false||abortednull|Flexible fiberoptic sigmoidoscopy|Procedure|false|false|C1550319|flexible sigmoidoscopynull|Flexible|Modifier|false|false||flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false|C1550319|sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false|C1550319|sigmoidoscopynull|Attempt|Event|false|false|C1550319|attemptnull|Feces|Finding|false|false|C1550319|stoolnull|Stool seat|Device|false|false||stoolnull|Vault|Anatomy|false|false|C1516084;C0016234;C1548917;C0037075;C0015733|vaultnull|Flexible fiberoptic sigmoidoscopy|Procedure|false|false||Flexible sigmoidoscopynull|Flexible|Modifier|false|false||Flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||sigmoidoscopynull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|PMH - past medical history|Finding|false|false||past medical history
null|Medical History|Finding|false|false||past medical historynull|Medical History|Finding|false|false||medical history ofnull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hypothyroidism|Disorder|false|false||hypothyroidismnull|Recent|Time|false|false||recentnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|null|Time|false|false||priornull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|DC Red No. 8|Drug|false|false||bright red
null|DC Red No. 8|Drug|false|false||bright rednull|Bright red color (finding)|Finding|false|false||bright rednull|Above average intellect|Finding|false|false||bright
null|ARID1B wt Allele|Finding|false|false||bright
null|ARID3A gene|Finding|false|false||brightnull|Bright|Modifier|false|false||brightnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Per rectum|Finding|false|false|C0034896;C4482211|per rectum
null|Rectal Route of Administration|Finding|false|false|C0034896;C4482211|per rectumnull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Rectal Diseases|Disorder|false|false|C0034896;C4482211|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Carcinoma in situ of rectum|Disorder|false|false|C0034896;C4482211|rectumnull|Procedure on rectum|Procedure|false|false|C0034896;C4482211|rectumnull|Pelvis>Rectum|Anatomy|false|false|C1527425;C4048189;C0869814;C0154062;C0034882;C0496867;C0496908|rectum
null|Rectum|Anatomy|false|false|C1527425;C4048189;C0869814;C0154062;C0034882;C0496867;C0496908|rectumnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Morning|Time|false|false||morningnull|Presentation|Finding|false|false||presentationnull|personal health|Finding|false|false||state of healthnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Health|Finding|false|false||healthnull|Home Health Aid|Subject|false|false||home health aidnull|home health encounter|Procedure|false|false||home healthnull|Home health care specialty|Title|false|false||home healthnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Health|Finding|false|false||healthnull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Helped|Finding|false|false||helpednull|Commodes|Device|false|false||commodenull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Per rectum|Finding|false|false|C0034896;C4482211|per rectum
null|Rectal Route of Administration|Finding|false|false|C0034896;C4482211|per rectumnull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Rectal Diseases|Disorder|false|false|C0034896;C4482211|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Carcinoma in situ of rectum|Disorder|false|false|C0034896;C4482211|rectumnull|Procedure on rectum|Procedure|false|false|C0034896;C4482211|rectumnull|Pelvis>Rectum|Anatomy|false|false|C0869814;C0154062;C0034882;C0496867;C0496908;C1527425;C4048189|rectum
null|Rectum|Anatomy|false|false|C0869814;C0154062;C0034882;C0496867;C0496908;C1527425;C4048189|rectumnull|next - HtmlLinkType|Finding|false|false||nextnull|Then|Time|false|false||next
null|Following|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Following|Time|false|false||subsequentnull|Episode of|Time|false|false||episodesnull|Home Health Aid|Subject|false|false||Home health aidnull|home health encounter|Procedure|false|false||Home healthnull|Home health care specialty|Title|false|false||Home healthnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Health|Finding|false|false||healthnull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Laboratory test finding|Lab|false|false||Labsnull|Leukocytes|Anatomy|false|false||WBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Primed lymphocyte test|Procedure|false|false||Pltnull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Neg - answer|Finding|false|false||negnull|Negative - qualifier|Modifier|false|false||negnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Blood and lymphatic system disorders|Disorder|false|false|C0034896;C4482211|bloodnull|peripheral blood|Finding|false|false|C0034896;C4482211|blood
null|Blood|Finding|false|false|C0034896;C4482211|blood
null|In Blood|Finding|false|false|C0034896;C4482211|bloodnull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Rectal Diseases|Disorder|false|false|C0034896;C4482211|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0034896;C4482211|rectum
null|Carcinoma in situ of rectum|Disorder|false|false|C0034896;C4482211|rectumnull|Procedure on rectum|Procedure|false|false|C0034896;C4482211|rectumnull|Pelvis>Rectum|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767;C0869814;C5890938;C1416798;C0154062;C0034882;C0496867;C0496908;C0019112|rectum
null|Rectum|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767;C0869814;C5890938;C1416798;C0154062;C0034882;C0496867;C0496908;C0019112|rectumnull|LARGE1 wt Allele|Finding|false|false|C0034896;C4482211|large
null|LARGE1 gene|Finding|false|false|C0034896;C4482211|largenull|Large|LabModifier|false|false||largenull|Hemorrhoids|Disorder|true|false|C0034896;C4482211|hemorrhoidsnull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|null|Finding|false|false||lavagenull|Irrigation|Procedure|false|false||lavagenull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|Maroon|Modifier|false|false||maroonnull|DHDDS gene|Finding|false|false||HDSnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Blood coagulation tests|Procedure|false|false||Coagnull|Supportive care|Procedure|false|false||supportive care
null|Palliative Care|Procedure|false|false||supportive carenull|Supportive assistance|Finding|false|false||supportivenull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|null|Finding|false|false||transfusionnull|Transfusion (procedure)|Procedure|false|false||transfusion
null|Blood Transfusion|Procedure|false|false||transfusionnull|Hemorrhage|Finding|false|false||bleedingnull|Hemodynamics|Finding|false|false||hemodynamicnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Concern|Finding|false|false||concernnull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleedingnull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleedingnull|Hemorrhage|Finding|false|false||bleedingnull|null|Finding|false|false||lavagenull|Irrigation|Procedure|false|false||lavagenull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Saline Solution|Drug|false|false||saline
null|Saline Solution|Drug|false|false||salinenull|Saline method|Procedure|false|false||salinenull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|arrival - ActRelationshipType|Finding|false|false|C3714591|arrivalnull|null|Event|false|false|C3714591|arrivalnull|Floor (anatomic)|Anatomy|false|false|C1552828;C1555577;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485;C1706079|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false|C3714591|patient
null|Specimen Type - Patient|Finding|false|false|C3714591|patient
null|Mail Claim Party - Patient|Finding|false|false|C3714591|patient
null|Report source - Patient|Finding|false|false|C3714591|patient
null|null|Finding|false|false|C3714591|patient
null|Disabled Person Code - Patient|Finding|false|false|C3714591|patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Table Frame - above|Finding|false|false|C3714591|abovenull|Upper|Modifier|false|false||abovenull|Recent|Time|false|false||recentnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|Intermittent|Time|false|false||intermittentnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Full|Modifier|false|false||Fullnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Hypothyroidism|Disorder|false|false||Hypothyroidismnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Protein-Energy Malnutrition|Finding|false|false||Protein calorie malnutritionnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|calorie unit of energy|LabModifier|false|false||calorie
null|Nutrition, Calories|LabModifier|false|false||calorie
null|kilocalorie|LabModifier|false|false||calorienull|Malnutrition|Disorder|false|false||malnutritionnull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Hemorrhoids|Disorder|false|false||Hemorrhoidsnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Bronchiectasis|Disorder|false|false||Bronchiectasisnull|Herpes zoster (disorder)|Disorder|false|false||Shinglesnull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Mitral Valve Insufficiency|Disorder|false|false||Mitral regurgitationnull|mitral|Modifier|false|false||Mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Offspring|Subject|false|false||children
null|Child|Subject|false|false||childrennull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Hemorrhoids|Disorder|false|false||hemorrhoidsnull|History of malignant neoplasm|Finding|true|false||history of cancernull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleedingnull|Hemorrhage|Finding|false|false||bleedingnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Supine Position|Modifier|false|false||supinenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Feeling comfortable|Finding|false|false||comfortablenull|Acute limbic encephalitis following transplant|Disorder|false|false||palenull|Body pale (finding)|Finding|false|false||pale
null|Pallor of skin|Finding|false|false||palenull|Pale color saturation|Modifier|false|false||pale
null|Pale color|Modifier|false|false||palenull|Eye|Anatomy|false|false|C5848506|Eyesnull|null|Attribute|false|false|C0015392|Eyesnull|ENT problem|Finding|false|false|C0150934;C0175196|ENT
null|NT5E gene|Finding|false|false|C0150934;C0175196|ENT
null|NT5E wt Allele|Finding|false|false|C0150934;C0175196|ENTnull|Structure of entorhinal cortex|Anatomy|false|false|C0262471;C3889152;C1417861|ENT
null|Ear, nose and throat|Anatomy|false|false|C0262471;C3889152;C1417861|ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|Heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|Heartnull|Systolic Murmurs|Finding|false|false||systolic murmurnull|Systole|Finding|false|false||systolicnull|Heart murmur|Finding|false|false||murmurnull|Axilla|Anatomy|false|false||axillanull|Lung|Anatomy|false|false|C3272310;C3540513;C4554671|Lungsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false|C0024109|CTA
null|CERNA3 gene|Finding|false|false|C0024109|CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false|C0024109|CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Carcinoma in situ of rectum|Disorder|false|false|C1550319;C0034896;C4482211|Rectum
null|Rectal Diseases|Disorder|false|false|C1550319;C0034896;C4482211|Rectum
null|Benign neoplasm of rectum|Disorder|false|false|C1550319;C0034896;C4482211|Rectum
null|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C1550319;C0034896;C4482211|Rectumnull|Procedure on rectum|Procedure|false|false|C1550319;C0034896;C4482211|Rectumnull|Pelvis>Rectum|Anatomy|false|false|C0005768;C0229664;C0005767;C0154062;C0034882;C0496867;C0496908;C0851353;C0869814|Rectum
null|Rectum|Anatomy|false|false|C0005768;C0229664;C0005767;C0154062;C0034882;C0496867;C0496908;C0851353;C0869814|Rectumnull|Dark color|Modifier|false|false||darknull|Maroon|Modifier|false|false||maroonnull|Blood and lymphatic system disorders|Disorder|false|false|C1550319;C0034896;C4482211|bloodnull|In Blood|Finding|false|false|C0034896;C4482211;C1550319|blood
null|peripheral blood|Finding|false|false|C0034896;C4482211;C1550319|blood
null|Blood|Finding|false|false|C0034896;C4482211;C1550319|bloodnull|Vault|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C0869814;C0005768;C0229664;C0005767;C0851353|vaultnull|LARGE1 wt Allele|Finding|true|false||large
null|LARGE1 gene|Finding|true|false||largenull|Large|LabModifier|false|false||largenull|Hemorrhoids|Disorder|true|false||hemorrhoidsnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C0678215;C0241137;C1546781;C0444099;C4750744;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C0678215;C0241137;C1546781;C0444099;C4750744;C0178298;C0496955|Skinnull|Acute limbic encephalitis following transplant|Disorder|false|false|C1123023;C4520765|palenull|Body pale (finding)|Finding|false|false|C1123023;C4520765|pale
null|Pallor of skin|Finding|false|false|C1123023;C4520765|palenull|Pale color saturation|Modifier|false|false||pale
null|Pale color|Modifier|false|false||palenull|Skin rash|Finding|true|false||rashes
null|Exanthema|Finding|true|false||rashesnull|Vascular Diseases|Disorder|false|false||Vascnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|AOX2P gene|Finding|false|false||AOx2null|Full|Modifier|false|false||fullnull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|Appropriate|Modifier|false|false||appropriatenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Supine Position|Modifier|false|false||supinenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Feeling comfortable|Finding|false|false||comfortablenull|Eye|Anatomy|false|false|C5848506|Eyesnull|null|Attribute|false|false|C0015392|Eyesnull|ENT problem|Finding|false|false|C0150934;C0175196|ENT
null|NT5E gene|Finding|false|false|C0150934;C0175196|ENT
null|NT5E wt Allele|Finding|false|false|C0150934;C0175196|ENTnull|Structure of entorhinal cortex|Anatomy|false|false|C0262471;C3889152;C1417861|ENT
null|Ear, nose and throat|Anatomy|false|false|C0262471;C3889152;C1417861|ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0039155;C0232257;C0153957;C0153500;C0795691;C0018808|Heart
null|Heart|Anatomy|false|false|C0039155;C0232257;C0153957;C0153500;C0795691;C0018808|Heartnull|Systolic Murmurs|Finding|false|false|C4037974;C0018787|systolic murmurnull|Systole|Finding|false|false|C4037974;C0018787|systolicnull|Heart murmur|Finding|false|false|C0004454;C4037974;C0018787|murmurnull|Axilla|Anatomy|false|false|C0018808|axillanull|Lung|Anatomy|false|false|C3540513;C4554671;C3272310;C0442739|Lungsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false|C0024109|CTA
null|CERNA3 gene|Finding|false|false|C0024109|CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false|C0024109|CTAnull|null|Finding|false|false|C0024109|unchangednull|About The Same|Modifier|false|false||unchangednull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Time|false|false||priornull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C5779628;C0015230;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C5779628;C0015230;C0178298;C0496955|Skinnull|Skin rash|Finding|true|false|C1123023;C4520765|rashes
null|Exanthema|Finding|true|false|C1123023;C4520765|rashesnull|Vascular Diseases|Disorder|false|false||Vascnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Full|Modifier|false|false||fullnull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|All extremities|Anatomy|false|false||all extremitiesnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|Appropriate|Modifier|false|false||appropriatenull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C1420113;C5960784;C4522245;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Flexible fiberoptic sigmoidoscopy|Procedure|false|false||Flexible Sigmoidoscopynull|Flexible|Modifier|false|false||Flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||Sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||Sigmoidoscopynull|null|Finding|false|false|C0026724|Mucosanull|Mucous Membrane|Anatomy|false|false|C1561514|Mucosanull|null|Finding|false|false|C0034896;C4482211;C0026724;C0227391;C0521377|mucosanull|Mucous Membrane|Anatomy|false|false|C1561514;C0154062;C0034882;C0496867;C0496908|mucosanull|Rectum and sigmoid colon|Anatomy|false|false|C0750873;C0869814;C0154062;C0034882;C0496867;C0496908;C0496864;C0153436;C1561514;C0154061;C0009373;C0496907|rectum and sigmoid colonnull|Carcinoma in situ of rectum|Disorder|false|false|C0034896;C4482211;C0521377;C0026724;C0227391|rectum
null|Rectal Diseases|Disorder|false|false|C0034896;C4482211;C0521377;C0026724;C0227391|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0034896;C4482211;C0521377;C0026724;C0227391|rectum
null|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0034896;C4482211;C0521377;C0026724;C0227391|rectumnull|Procedure on rectum|Procedure|false|false|C0034896;C4482211;C0521377|rectumnull|Pelvis>Rectum|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C1561514;C0869814;C0496864;C0153436;C0750873;C0154061;C0009373;C0496907|rectum
null|Rectum|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C1561514;C0869814;C0496864;C0153436;C0750873;C0154061;C0009373;C0496907|rectumnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0034896;C4482211;C0227391;C0521377|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0034896;C4482211;C0227391;C0521377|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C1561514;C0496864;C0153436;C0154061;C0009373;C0496907;C0154062;C0034882;C0496867;C0496908|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436;C0750873;C0154061;C0009373;C0496907|sigmoidnull|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391;C0034896;C4482211;C0521377|colon
null|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391;C0034896;C4482211;C0521377|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0227391;C0227391;C0034896;C4482211;C0521377|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0521377;C0227391;C0009368;C4071907;C0034896;C4482211|colonnull|Colon structure (body structure)|Anatomy|false|false|C0496864;C0153436;C0154061;C0009373;C0496907;C0750873|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0496864;C0153436;C0154061;C0009373;C0496907;C0750873|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Hemorrhage|Finding|true|false||bleedingnull|Source|Finding|true|false||sourcesnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Extent|Modifier|false|false||extent ofnull|Extent|Modifier|false|false||extentnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C5400798;C1418885;C1425030;C4319962;C0496864;C0153436;C4723750;C1547310;C0750873;C1521827;C0009373;C0154061;C0496907|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C0496864;C0153436;C0009373;C0154061;C0496907|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0009368;C4071907;C0227391|colonnull|Colon structure (body structure)|Anatomy|false|false|C1418885;C1425030;C4319962;C0496864;C0153436;C0009373;C0154061;C0496907;C5400798;C0750873;C4723750;C1547310|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C1418885;C1425030;C4319962;C0496864;C0153436;C0009373;C0154061;C0496907;C5400798;C0750873;C4723750;C1547310|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false|C0227391;C0009368;C4071907|poor
null|Patient Condition Code - Poor|Finding|false|false|C0227391;C0009368;C4071907|poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|PREP gene|Finding|false|false|C0009368;C4071907;C0227391|prep
null|PITRM1 gene|Finding|false|false|C0009368;C4071907;C0227391|prep
null|PITRM1 wt Allele|Finding|false|false|C0009368;C4071907;C0227391|prepnull|null|Procedure|false|false|C0227391;C0009368;C4071907|prepnull|Preparation|Event|false|false|C0227391|prepnull|impression (attitude)|Finding|false|false||Impression
null|EKG impression|Finding|false|false||Impressionnull|null|Finding|false|false|C0026724;C0034896;C4482211;C0521377|mucosanull|Mucous Membrane|Anatomy|false|false|C1561514;C0154062;C0034882;C0496867;C0496908|mucosanull|Rectum and sigmoid colon|Anatomy|false|false|C0154061;C0009373;C0496907;C0496864;C0153436;C1561514;C0154062;C0034882;C0496867;C0496908;C0869814;C0750873|rectum and sigmoid colonnull|Carcinoma in situ of rectum|Disorder|false|false|C0227391;C0034896;C4482211;C0026724;C0521377;C0227391|rectum
null|Rectal Diseases|Disorder|false|false|C0227391;C0034896;C4482211;C0026724;C0521377;C0227391|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0227391;C0034896;C4482211;C0026724;C0521377;C0227391|rectum
null|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0227391;C0034896;C4482211;C0026724;C0521377;C0227391|rectumnull|Procedure on rectum|Procedure|false|false|C0034896;C4482211;C0521377|rectumnull|Pelvis>Rectum|Anatomy|false|false|C0869814;C0496864;C0153436;C1561514;C0154062;C0034882;C0496867;C0496908|rectum
null|Rectum|Anatomy|false|false|C0869814;C0496864;C0153436;C1561514;C0154062;C0034882;C0496867;C0496908|rectumnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0034896;C4482211;C0521377;C0227391;C0009368;C4071907|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0034896;C4482211;C0521377;C0227391;C0009368;C4071907|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C0496864;C0153436;C0154061;C0009373;C0496907;C0750873|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436;C0154061;C0009373;C0496907;C0750873;C0154062;C0034882;C0496867;C0496908|sigmoidnull|Carcinoma in situ of colon|Disorder|false|false|C0227391;C0521377;C0227391;C0009368;C4071907|colon
null|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0227391;C0521377;C0227391;C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0227391;C0521377;C0227391;C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0009368;C4071907;C0227391;C0227391;C0521377|colonnull|Colon structure (body structure)|Anatomy|false|false|C0750873;C0496864;C0153436;C0154061;C0009373;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0750873;C0496864;C0153436;C0154061;C0009373;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Hemorrhage|Finding|true|false||bleedingnull|Source|Finding|true|false||sourcesnull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||blood
null|In Blood|Finding|true|false||bloodnull|Extent|Modifier|false|false||extent ofnull|Extent|Modifier|false|false||extentnull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0227391;C0009368;C4071907|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0227391;C0009368;C4071907|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C1418885;C1425030;C4319962;C0496864;C0153436;C1521827;C0750873;C5400798;C0009373;C0154061;C0496907;C4723750;C1547310|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C0009373;C0154061;C0496907;C0496864;C0153436|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0227391;C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C5400798;C4723750;C1547310;C0750873;C1418885;C1425030;C4319962;C0496864;C0153436|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C5400798;C4723750;C1547310;C0750873;C1418885;C1425030;C4319962;C0496864;C0153436|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false|C0009368;C4071907;C0227391|poor
null|Patient Condition Code - Poor|Finding|false|false|C0009368;C4071907;C0227391|poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|PREP gene|Finding|false|false|C0227391;C0009368;C4071907|prep
null|PITRM1 gene|Finding|false|false|C0227391;C0009368;C4071907|prep
null|PITRM1 wt Allele|Finding|false|false|C0227391;C0009368;C4071907|prepnull|null|Procedure|false|false|C0009368;C4071907;C0227391|prepnull|Preparation|Event|false|false|C0227391|prepnull|Consent Type - Sigmoidoscopy|Procedure|false|false|C0227391;C0227391|sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false|C0227391;C0227391|sigmoidoscopynull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436;C0750873;C1548917;C0037075;C0009373;C0154061;C0496907|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C1548917;C0037075;C0009373;C0154061;C0496907;C0496864;C0153436|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0227391;C0009368;C4071907;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0009368;C4071907;C0227391|colonnull|Colon structure (body structure)|Anatomy|false|false|C0750873;C0496864;C0153436;C0009373;C0154061;C0496907|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0750873;C0496864;C0153436;C0009373;C0154061;C0496907|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Recommendation|Finding|false|false||Recommendationsnull|Hemorrhage|Finding|false|false||bleedingnull|Full|Modifier|false|false||fullnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|PREP gene|Finding|false|false||prep
null|PITRM1 gene|Finding|false|false||prep
null|PITRM1 wt Allele|Finding|false|false||prepnull|null|Procedure|false|false||prepnull|Preparation|Event|false|false||prepnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|PMH - past medical history|Finding|false|false||past medical history
null|Medical History|Finding|false|false||past medical historynull|Medical History|Finding|false|false||medical history ofnull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Hemorrhoids|Disorder|false|false||hemorrhoidsnull|null|Time|false|false||priornull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Hematochezia|Disorder|false|false|C0034896;C4482211|bright red blood per rectumnull|DC Red No. 8|Drug|false|false||bright red
null|DC Red No. 8|Drug|false|false||bright rednull|Bright red color (finding)|Finding|false|false||bright rednull|Above average intellect|Finding|false|false||bright
null|ARID1B wt Allele|Finding|false|false||bright
null|ARID3A gene|Finding|false|false||brightnull|Bright|Modifier|false|false||brightnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Rectal hemorrhage|Finding|false|false|C0034896;C4482211|blood per rectumnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Per rectum|Finding|false|false|C0034896;C4482211|per rectum
null|Rectal Route of Administration|Finding|false|false|C0034896;C4482211|per rectumnull|Neoplasm of uncertain or unknown behavior of rectum|Disorder|false|false|C0034896;C4482211;C1548802|rectum
null|Rectal Diseases|Disorder|false|false|C0034896;C4482211;C1548802|rectum
null|Benign neoplasm of rectum|Disorder|false|false|C0034896;C4482211;C1548802|rectum
null|Carcinoma in situ of rectum|Disorder|false|false|C0034896;C4482211;C1548802|rectumnull|Procedure on rectum|Procedure|false|false|C1548802;C0034896;C4482211|rectumnull|Pelvis>Rectum|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C1527425;C4048189;C0267596;C4319827;C0039869;C0869814;C1547295;C1547229;C0018932|rectum
null|Rectum|Anatomy|false|false|C0154062;C0034882;C0496867;C0496908;C1527425;C4048189;C0267596;C4319827;C0039869;C0869814;C1547295;C1547229;C0018932|rectumnull|Thought|Finding|false|false|C0034896;C4482211|thought
null|null|Finding|false|false|C0034896;C4482211|thoughtnull|Admission Level of Care Code - Acute|Finding|false|false|C1548802;C0034896;C4482211|acute
null|Acute - Triage Code|Finding|false|false|C1548802;C0034896;C4482211|acutenull|acute|Time|false|false||acutenull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C0869814;C0154062;C0034882;C0496867;C0496908;C1547295;C1547229|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Hemorrhage|Finding|false|false||bleednull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Flexible fiberoptic sigmoidoscopy|Procedure|false|false||flexible sigmoidoscopynull|Flexible|Modifier|false|false||flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||sigmoidoscopynull|Identifiable Class|Finding|false|false||identifiablenull|Identified|Modifier|false|false||identifiablenull|Source (property) (qualifier value)|Finding|true|false||source
null|Term Source|Finding|true|false||source
null|Source|Finding|true|false||sourcenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|4 Days|Time|false|false||4 daysnull|day|Time|false|false||daysnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Acute gastrointestinal hemorrhage|Disorder|false|false||Acute GI Bleednull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Gastrointestinal Hemorrhage|Finding|false|false||GI Bleednull|Hemorrhage|Finding|false|false||Bleednull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Hematochezia|Disorder|false|false|C1548802|BRBPRnull|Body Site Modifier - Lower|Anatomy|false|false|C0449416;C1705919;C4521696;C2003888;C0018932|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Source (property) (qualifier value)|Finding|false|false|C1548802|source
null|Term Source|Finding|false|false|C1548802|source
null|Source|Finding|false|false|C1548802|sourcenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|Anemia|Disorder|true|false||anemianull|Anemia <Anemiaceae>|Entity|true|false||anemianull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Further|Modifier|false|false||furthernull|Flexible fiberoptic sigmoidoscopy|Procedure|false|false||flexible sigmoidoscopynull|Flexible|Modifier|false|false||flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||sigmoidoscopynull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Invasive|Modifier|false|false||invasivenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|aborted - QueryStatusCode|Finding|false|false||aborted
null|aborted - ActStatus|Finding|false|false||aborted
null|Order aborted|Finding|false|false||abortednull|Flexible|Modifier|false|false||flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||sigmoidoscopynull|Copious|Finding|false|false||copiousnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Rectal Dosage Form|Drug|false|false||rectalnull|Rectal Route of Administration|Finding|false|false|C1550319|rectal
null|Rectal (intended site)|Finding|false|false|C1550319|rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||rectalnull|rectal|Modifier|false|false||rectalnull|Vault|Anatomy|false|false|C1527425;C4521903;C1720594|vaultnull|Then - dosing instruction fragment|Finding|false|false|C1550319|thennull|Then|Time|false|false||thennull|Success|Finding|false|false||successfulnull|Successful|Modifier|false|false||successfulnull|Flexible|Modifier|false|false||flexiblenull|Consent Type - Sigmoidoscopy|Procedure|false|false||sigmoidoscopy
null|Sigmoidoscopy (procedure)|Procedure|false|false||sigmoidoscopynull|Identifiable Class|Finding|false|false||identifiablenull|Identified|Modifier|false|false||identifiablenull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Hemorrhage|Finding|false|false||bleedingnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Hemoglobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|chrysarobin|Drug|false|false||hemoglobin
null|Hemoglobin|Drug|false|false||hemoglobinnull|Hemoglobin finding|Finding|false|false||hemoglobinnull|Hemoglobin measurement|Procedure|false|false||hemoglobinnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recent|Time|false|false||recentnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Activity of daily living (function)|Finding|false|false||ADLsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Vitamin D Drug Class|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|D Vitamin|Drug|false|false||vitamin D
null|Vitamin D [EPC]|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|Vitamin D Drug Class|Drug|false|false||vitamin Dnull|Vitamin D measurement|Procedure|false|false||vitamin Dnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Calcitonin Precursor, human|Drug|false|false||calcitonin
null|human calcitonin|Drug|false|false||calcitonin
null|human calcitonin|Drug|false|false||calcitonin
null|human calcitonin|Drug|false|false||calcitonin
null|Calcitonin Precursor, human|Drug|false|false||calcitonin
null|Calcitonin [EPC]|Drug|false|false||calcitonin
null|Recombinant Calcitonin|Drug|false|false||calcitonin
null|Recombinant Calcitonin|Drug|false|false||calcitonin
null|Recombinant Calcitonin|Drug|false|false||calcitonin
null|calcitonin|Drug|false|false||calcitonin
null|calcitonin|Drug|false|false||calcitonin
null|calcitonin|Drug|false|false||calcitoninnull|CALCA gene|Finding|false|false||calcitoninnull|Calcitonin measurement|Procedure|false|false||calcitoninnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|good effect|Finding|false|false||good effectnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|null|Disorder|false|false||Severe Protein Calorie Malnutritionnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Protein-Energy Malnutrition|Finding|false|false||Protein Calorie Malnutritionnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|calorie unit of energy|LabModifier|false|false||Calorie
null|Nutrition, Calories|LabModifier|false|false||Calorie
null|kilocalorie|LabModifier|false|false||Calorienull|Malnutrition|Disorder|false|false||Malnutritionnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Charts (publication)|Finding|false|false||chartnull|chart [medical device]|Device|false|false||chartnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Response Modality - Bolus|Finding|false|false||bolus
null|Bolus of ingested food|Finding|false|false||bolusnull|bolus infusion|Procedure|false|false||bolusnull|Bolus Dosing Unit|LabModifier|false|false||bolusnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Feeds|Finding|false|false||feedsnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|At home|Finding|false|false||At homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Full|Modifier|false|false||fullnull|NUTREN|Drug|false|false||Nutrennull|monoclonal antibody CAL|Drug|false|false|C0228225|Cal
null|monoclonal antibody CAL|Drug|false|false|C0228225|Calnull|FBLIM1 wt Allele|Finding|false|false|C0228225|Cal
null|GOPC gene|Finding|false|false|C0228225|Cal
null|FBLP1 gene|Finding|false|false|C0228225|Cal
null|GOPC wt Allele|Finding|false|false|C0228225|Calnull|Structure of calcar avis|Anatomy|false|false|C1425021;C1825283;C5890925;C3273482;C1530795;C1135160;C4546282;C1332410|Calnull|calorie unit of energy|LabModifier|false|false||Cal
null|Nutrition, Calories|LabModifier|false|false||Cal
null|kilocalorie|LabModifier|false|false||Calnull|BID protein, human|Drug|false|false|C0228225|BID
null|BID protein, human|Drug|false|false|C0228225|BIDnull|Body integrity dysphoria|Disorder|false|false|C0228225|BIDnull|BID gene|Finding|false|false|C0228225|BIDnull|Twice a day|Time|false|false||BIDnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Nutrition (function)|Finding|false|false||nutrition
null|Nutritional status|Finding|false|false||nutrition
null|Nutrition outcomes|Finding|false|false||nutritionnull|Feeding and dietary regimes|Procedure|false|false||nutrition
null|Nutritional Study|Procedure|false|false||nutritionnull|Science of nutrition|Title|false|false||nutritionnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C0242297;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Dietary Supplementation|Procedure|false|false|C0226896|supplementationnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|mirtazapine|Drug|false|false||mirtazapine
null|mirtazapine|Drug|false|false||mirtazapinenull|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxine
null|levothyroxine|Drug|false|false||levothyroxinenull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|CODE STATUS|Procedure|false|false||Code statusnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|daunorubicin|Drug|false|false||DNR
null|daunorubicin|Drug|false|false||DNRnull|Do not resuscitate status|Finding|false|false||DNR
null|Do-Not-Resuscitate Orders|Finding|false|false||DNRnull|null|Attribute|false|false||DNRnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Source (property) (qualifier value)|Finding|true|false||source
null|Term Source|Finding|true|false||source
null|Source|Finding|true|false||sourcenull|Hemorrhage|Finding|true|false||bleedingnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|consider|Finding|false|false||considernull|Future|Time|false|false||futurenull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Hemorrhage|Finding|false|false||bleedingnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Goals of Care|Procedure|false|false||goals of carenull|What subject filter - Goals|Finding|false|false||goals
null|objective (goal)|Finding|false|false||goals
null|treatment goals|Finding|false|false||goalsnull|null|Attribute|false|false||goalsnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|encouragement|Finding|false|false||encouragementnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|polyethylene glycol 400|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycols|Drug|false|false||PEG
null|polyethylene glycol 400|Drug|false|false||PEGnull|PEG Study|Procedure|false|false||PEG
null|Percutaneous endoscopic gastrostomy|Procedure|false|false||PEGnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Dietary Supplementation|Procedure|false|false||supplementationnull|Malnutrition|Disorder|false|false||malnutritionnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||Dailynull|Daily|Time|false|false||DAILYnull|Calcium 500+D|Drug|false|false||Calcium 500 + D
null|Calcium 500+D|Drug|false|false||Calcium 500 + Dnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|calcium carbonate|Drug|false|false||calcium carbonate
null|calcium carbonate|Drug|false|false||calcium carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|carbonate ion|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonatenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|mirtazapine|Drug|false|false||Mirtazapine
null|mirtazapine|Drug|false|false||Mirtazapinenull|Once a day, at bedtime|Time|false|false||QHSnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|alendronate sodium|Drug|false|false||Alendronate Sodium
null|alendronate sodium|Drug|false|false||Alendronate Sodiumnull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|salmon calcitonin|Drug|false|false||Calcitonin Salmon
null|salmon calcitonin|Drug|false|false||Calcitonin Salmon
null|salmon calcitonin|Drug|false|false||Calcitonin Salmonnull|Calcitonin Precursor, human|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|Calcitonin Precursor, human|Drug|false|false||Calcitonin
null|Calcitonin [EPC]|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitoninnull|CALCA gene|Finding|false|false||Calcitoninnull|Calcitonin measurement|Procedure|false|false||Calcitoninnull|salmon allergenic extract|Drug|false|false||Salmon
null|salmon allergenic extract|Drug|false|false||Salmon
null|Salmon (substance)|Drug|false|false||Salmon
null|null|Drug|false|false||Salmonnull|Salmon|Entity|false|false||Salmon
null|Salmo salar|Entity|false|false||Salmonnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Tobacco containing mixture|Drug|false|false||NAS
null|N-acetylserotonin|Drug|false|false||NASnull|Neonatal Abstinence Syndrome|Disorder|false|false||NASnull|null|Finding|false|false||NASnull|National Academy of Sciences (U.S.)|Entity|false|false||NASnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|Four times daily|Time|false|false||QIDnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||Dailynull|Daily|Time|false|false||DAILYnull|salmon calcitonin|Drug|false|false||Calcitonin Salmon
null|salmon calcitonin|Drug|false|false||Calcitonin Salmon
null|salmon calcitonin|Drug|false|false||Calcitonin Salmonnull|Calcitonin Precursor, human|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|human calcitonin|Drug|false|false||Calcitonin
null|Calcitonin Precursor, human|Drug|false|false||Calcitonin
null|Calcitonin [EPC]|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|Recombinant Calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitonin
null|calcitonin|Drug|false|false||Calcitoninnull|CALCA gene|Finding|false|false||Calcitoninnull|Calcitonin measurement|Procedure|false|false||Calcitoninnull|salmon allergenic extract|Drug|false|false||Salmon
null|salmon allergenic extract|Drug|false|false||Salmon
null|Salmon (substance)|Drug|false|false||Salmon
null|null|Drug|false|false||Salmonnull|Salmon|Entity|false|false||Salmon
null|Salmo salar|Entity|false|false||Salmonnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Tobacco containing mixture|Drug|false|false||NAS
null|N-acetylserotonin|Drug|false|false||NASnull|Neonatal Abstinence Syndrome|Disorder|false|false||NASnull|null|Finding|false|false||NASnull|National Academy of Sciences (U.S.)|Entity|false|false||NASnull|Daily|Time|false|false||DAILYnull|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodium
null|levothyroxine sodium|Drug|false|false||Levothyroxine Sodiumnull|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|Synthetic Levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxine
null|levothyroxine|Drug|false|false||Levothyroxinenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|microgram|LabModifier|false|false||mcgnull|Daily|Time|false|false||DAILYnull|mirtazapine|Drug|false|false||Mirtazapine
null|mirtazapine|Drug|false|false||Mirtazapinenull|Once a day, at bedtime|Time|false|false||QHSnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|alendronate sodium|Drug|false|false||Alendronate Sodium
null|alendronate sodium|Drug|false|false||Alendronate Sodiumnull|alendronate|Drug|false|false||Alendronate
null|alendronate|Drug|false|false||Alendronatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Calcium 500+D|Drug|false|false||Calcium 500 + D
null|Calcium 500+D|Drug|false|false||Calcium 500 + Dnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|calcium carbonate|Drug|false|false||calcium carbonate
null|calcium carbonate|Drug|false|false||calcium carbonatenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|carbonate ion|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonate
null|Carbonates|Drug|false|false||carbonatenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|artificial tears (medication)|Drug|false|false||Artificial Tears
null|Lubricant Eye Drops|Drug|false|false||Artificial Tears
null|Artificial Tears|Drug|false|false||Artificial Tearsnull|Artificial (qualifier value)|Modifier|false|false||Artificialnull|Tears (substance)|Finding|false|false||Tears
null|null|Finding|false|false||Tears
null|Tears specimen|Finding|false|false||Tearsnull|Drops - Drug Form|Drug|false|false||DROPnull|Dropping|Event|false|false||DROPnull|Drop (unit of presentation)|LabModifier|false|false||DROP
null|Drop British|LabModifier|false|false||DROP
null|Drop Dosing Unit|LabModifier|false|false||DROP
null|Medical Drop|LabModifier|false|false||DROP
null|Drop Unit of Volume|LabModifier|false|false||DROPnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false|C5848506|EYESnull|null|Attribute|false|false|C0015392|EYESnull|Four times daily|Time|false|false||QIDnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Acute gastrointestinal hemorrhage|Disorder|false|false||Acute GI Bleednull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Gastrointestinal Hemorrhage|Finding|false|false||GI Bleednull|Hemorrhage|Finding|false|false||Bleednull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Compression fracture|Finding|false|false||compression fracturenull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Fracture|Disorder|false|false||fracturenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|null|Disorder|false|false||Severe Protein Calorie Malnutritionnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Protein-Energy Malnutrition|Finding|false|false||Protein Calorie Malnutritionnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|calorie unit of energy|LabModifier|false|false||Calorie
null|Nutrition, Calories|LabModifier|false|false||Calorie
null|kilocalorie|LabModifier|false|false||Calorienull|Malnutrition|Disorder|false|false||Malnutritionnull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Confusion|Disorder|false|false||Confusednull|Precaution Code - Confused|Finding|false|false||Confused
null|Clouded consciousness|Finding|false|false||Confusednull|Sometimes|Time|false|false||sometimesnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Gastrointestinal Hemorrhage|Finding|false|false||gastrointestinal bleedingnull|Gastrointestinal attachment|Finding|false|false||gastrointestinalnull|gastrointestinal|Modifier|false|false||gastrointestinalnull|Hemorrhage|Finding|false|false||bleedingnull|Hospital specialist|Subject|false|false||specialistsnull|Flexible|Modifier|false|false||flexiblenull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Hemorrhage|Finding|false|false||bleedingnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Levels (qualifier value)|Modifier|false|false||levelsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Ready for discharge|Finding|false|false||ready for dischargenull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Future|Time|false|false||futurenull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|Hemorrhage|Finding|false|false||bleedingnull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|true||doctornull|Physicians|Subject|false|false||doctornull|Goals of Care|Procedure|false|false||goals of carenull|What subject filter - Goals|Finding|false|false||goals
null|objective (goal)|Finding|false|false||goals
null|treatment goals|Finding|false|false||goalsnull|null|Attribute|false|false||goalsnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions