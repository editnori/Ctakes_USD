 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|true|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|true|false|false|C1717415||Allergies
Event|Event|Allergies|181,190|true|false|false|||Allergies
Finding|Pathologic Function|Allergies|181,190|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|206,215|true|false|false|||Reactions
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|252,261|false|false|false|||Shortness
Attribute|Clinical Attribute|Chief Complaint|252,271|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|Chief Complaint|252,271|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|Chief Complaint|265,271|false|false|false|C0225386|Breath|breath
Finding|Classification|Chief Complaint|274,279|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|280,288|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|280,288|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|292,310|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|301,310|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|301,310|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|301,310|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|301,310|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|301,310|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|369,381|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|369,381|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|383,397|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|History of Present Illness|383,397|false|false|false|||hyperlipidemia
Finding|Finding|History of Present Illness|383,397|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Disorder|Disease or Syndrome|History of Present Illness|399,407|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|History of Present Illness|399,407|false|false|false|||diabetes
Event|Event|History of Present Illness|409,417|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|421,428|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|History of Present Illness|421,428|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|History of Present Illness|421,428|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|History of Present Illness|421,428|false|false|false|||insulin
Finding|Gene or Genome|History of Present Illness|421,428|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|History of Present Illness|421,428|false|false|false|C0202098|Insulin measurement|insulin
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|421,436|false|false|false|C5442411|Insulin therapy|insulin therapy
Event|Event|History of Present Illness|429,436|false|false|false|||therapy
Finding|Finding|History of Present Illness|429,436|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|History of Present Illness|429,436|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|429,436|false|false|false|C0087111|Therapeutic procedure|therapy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|442,452|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|453,462|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|History of Present Illness|463,469|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|History of Present Illness|463,469|false|false|false|||stroke
Finding|Finding|History of Present Illness|463,469|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|History of Present Illness|479,482|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|History of Present Illness|483,488|false|false|false|C1300072|Tumor stage|stage
Event|Event|History of Present Illness|496,506|false|false|false|||presenting
Finding|Idea or Concept|History of Present Illness|496,506|false|false|false|C0449450|Presentation|presenting
Event|Event|History of Present Illness|512,519|false|false|false|||fatigue
Finding|Sign or Symptom|History of Present Illness|512,519|false|false|false|C0015672|Fatigue|fatigue
Event|Event|History of Present Illness|524,531|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|524,531|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|524,531|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|536,544|false|false|false|||exertion
Finding|Organism Function|History of Present Illness|536,544|false|false|false|C0015264|Exertion|exertion
Event|Event|History of Present Illness|546,549|false|false|false|||DOE
Finding|Sign or Symptom|History of Present Illness|546,549|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|History of Present Illness|577,582|false|false|false|||worse
Finding|Finding|History of Present Illness|577,582|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|577,582|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Body Substance|History of Present Illness|627,634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|627,634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|627,634|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|635,640|false|false|false|||noted
Event|Event|History of Present Illness|641,644|false|false|false|||DOE
Event|Event|History of Present Illness|649,658|false|false|false|||shortness
Finding|Body Substance|History of Present Illness|663,669|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|671,674|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|671,674|false|false|false|C0013404|Dyspnea|SOB
Finding|Functional Concept|History of Present Illness|681,688|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|684,688|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|684,688|false|false|false|C1742913|REST protein, human|rest
Finding|Daily or Recreational Activity|History of Present Illness|684,688|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|684,688|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|684,688|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Event|Event|History of Present Illness|703,707|false|false|false|||felt
Event|Event|History of Present Illness|713,718|false|false|false|||tired
Finding|Finding|History of Present Illness|713,718|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|History of Present Illness|713,718|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|History of Present Illness|713,718|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|History of Present Illness|736,741|true|false|false|||notes
Attribute|Clinical Attribute|History of Present Illness|745,756|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|History of Present Illness|745,756|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|History of Present Illness|745,756|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|History of Present Illness|745,756|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|History of Present Illness|757,763|true|false|false|||issues
Event|Event|History of Present Illness|794,798|true|false|false|||walk
Event|Event|History of Present Illness|815,818|true|false|false|||DOE
Finding|Sign or Symptom|History of Present Illness|815,818|true|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|History of Present Illness|824,829|false|false|false|||feels
Event|Event|History of Present Illness|830,833|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|830,833|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|854,862|false|false|false|||distance
Event|Event|History of Present Illness|871,877|false|false|false|||unsure
Finding|Finding|History of Present Illness|871,877|false|false|false|C0087130|Uncertainty|unsure
Event|Event|History of Present Illness|911,917|false|false|false|||states
Attribute|Clinical Attribute|History of Present Illness|927,936|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|927,936|false|false|false|||breathing
Finding|Finding|History of Present Illness|927,936|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|927,936|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|927,936|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|927,936|false|false|false|C1160636|respiratory system process|breathing
Event|Event|History of Present Illness|937,945|false|false|false|||improves
Drug|Organic Chemical|History of Present Illness|951,960|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|History of Present Illness|951,960|false|false|false|C0001927|albuterol|albuterol
Event|Event|History of Present Illness|951,960|false|false|false|||albuterol
Event|Event|History of Present Illness|971,975|false|false|false|||gets
Disorder|Disease or Syndrome|History of Present Illness|1005,1008|false|false|false|C4522181|Brachial Amyotrophic Diplegia|bad
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1005,1008|false|false|false|C1530798|BAD protein, human|bad
Drug|Biologically Active Substance|History of Present Illness|1005,1008|false|false|false|C1530798|BAD protein, human|bad
Finding|Gene or Genome|History of Present Illness|1005,1008|false|false|false|C1366450|BAD gene|bad
Drug|Organic Chemical|History of Present Illness|1009,1014|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1009,1014|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1009,1014|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1009,1014|false|false|false|C0010200|Coughing|cough
Finding|Idea or Concept|History of Present Illness|1024,1029|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|1024,1029|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|History of Present Illness|1030,1033|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1040,1046|true|false|false|||denies
Event|Event|History of Present Illness|1058,1064|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1058,1064|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1066,1072|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1066,1072|true|false|false|C0085593|Chills|chills
Finding|Sign or Symptom|History of Present Illness|1077,1089|true|false|false|C0028081|Night sweats|night sweats
Event|Event|History of Present Illness|1083,1089|false|false|false|||sweats
Finding|Body Substance|History of Present Illness|1083,1089|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|1083,1089|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Anatomy|Body Location or Region|History of Present Illness|1094,1099|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1094,1099|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1101,1105|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1101,1105|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1101,1105|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1101,1105|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1107,1113|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|1107,1113|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1107,1113|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1118,1127|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|1118,1127|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Disorder|Disease or Syndrome|Past Medical History|1156,1159|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1156,1159|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|1156,1159|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|1156,1159|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|1156,1159|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|1156,1159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|1156,1159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1156,1159|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Past Medical History|1160,1164|false|false|false|||RISK
Finding|Idea or Concept|Past Medical History|1160,1164|false|false|false|C0035647|Risk|RISK
Attribute|Clinical Attribute|Past Medical History|1160,1172|false|false|false|C1830376||RISK FACTORS
Finding|Finding|Past Medical History|1160,1172|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Finding|Intellectual Product|Past Medical History|1160,1172|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|RISK FACTORS
Event|Event|Past Medical History|1165,1172|false|false|false|||FACTORS
Disorder|Disease or Syndrome|Past Medical History|1175,1183|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Event|Event|Past Medical History|1175,1183|false|false|false|||Diabetes
Disorder|Disease or Syndrome|Past Medical History|1186,1198|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|1201,1213|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|1201,1213|false|false|false|||Hypertension
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1217,1224|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Past Medical History|1217,1224|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|Patient History|1259,1266|false|false|false|||MEDICAL
Finding|Functional Concept|Patient History|1259,1266|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Idea or Concept|Patient History|1259,1266|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Finding|Intellectual Product|Patient History|1259,1266|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|MEDICAL
Procedure|Health Care Activity|Patient History|1259,1266|false|false|false|C0199168|Medical service|MEDICAL
Disorder|Disease or Syndrome|Patient History|1278,1290|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Patient History|1278,1290|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Patient History|1291,1305|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Patient History|1291,1305|false|false|false|||Hyperlipidemia
Finding|Finding|Patient History|1291,1305|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Disorder|Disease or Syndrome|Patient History|1306,1314|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Patient History|1306,1323|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Event|Event|Patient History|1315,1323|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|Patient History|1327,1334|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Patient History|1327,1334|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Patient History|1327,1334|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Patient History|1327,1334|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Patient History|1327,1334|false|false|false|C0202098|Insulin measurement|insulin
Procedure|Therapeutic or Preventive Procedure|Patient History|1327,1342|false|false|false|C5442411|Insulin therapy|insulin therapy
Event|Event|Patient History|1335,1342|false|false|false|||therapy
Finding|Finding|Patient History|1335,1342|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Patient History|1335,1342|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Patient History|1335,1342|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Patient History|1344,1345|false|false|false|||/
Anatomy|Body Part, Organ, or Organ Component|Patient History|1347,1357|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Patient History|1358,1367|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Patient History|1368,1374|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Patient History|1368,1374|false|false|false|||stroke
Finding|Finding|Patient History|1368,1374|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Patient History|1382,1385|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Patient History|1386,1391|false|false|false|C1300072|Tumor stage|stage
Disorder|Disease or Syndrome|Patient History|1399,1402|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|Patient History|1399,1402|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|Patient History|1399,1402|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Event|Event|Family Medical History|1441,1447|false|false|false|||Denies
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1448,1455|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|1448,1455|true|false|false|C1314974|Cardiac attachment|cardiac
Finding|Classification|Family Medical History|1456,1462|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|1456,1462|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|1456,1462|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|1456,1462|true|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|1456,1470|true|false|false|C0241889|Family Medical History|family history
Event|Event|Family Medical History|1463,1470|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|1463,1470|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1463,1470|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1463,1470|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Classification|Family Medical History|1472,1478|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|Family Medical History|1472,1478|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|Family Medical History|1472,1478|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|Family Medical History|1472,1478|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Disorder|Disease or Syndrome|Family Medical History|1492,1495|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|1492,1495|false|false|false|||HTN
Event|Event|Family Medical History|1508,1524|false|false|false|||non-contributory
Procedure|Health Care Activity|General Exam|1543,1552|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|General Exam|1553,1557|false|false|false|||exam
Finding|Functional Concept|General Exam|1553,1557|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|1553,1557|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|1559,1566|false|false|false|||GENERAL
Finding|Classification|General Exam|1559,1566|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|1559,1566|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|1568,1576|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|General Exam|1581,1585|false|false|false|C2713234||Mood
Event|Event|General Exam|1581,1585|false|false|false|||Mood
Finding|Conceptual Entity|General Exam|1581,1585|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|General Exam|1581,1585|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|General Exam|1581,1585|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Event|Event|General Exam|1587,1593|false|false|false|||affect
Event|Event|General Exam|1594,1605|false|false|false|||appropriate
Event|Event|General Exam|1611,1612|false|false|false|||T
Event|Event|General Exam|1619,1621|false|false|false|||BP
Event|Event|General Exam|1648,1651|false|false|false|||sat
Anatomy|Body Location or Region|General Exam|1664,1669|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|1671,1675|false|false|false|||NCAT
Anatomy|Body Part, Organ, or Organ Component|General Exam|1677,1683|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|1677,1683|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|1677,1683|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|1677,1683|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|1684,1693|false|false|false|||anicteric
Finding|Finding|General Exam|1684,1693|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|1695,1700|false|false|false|||PERRL
Finding|Finding|General Exam|1695,1700|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|1702,1706|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|1708,1719|true|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|General Exam|1708,1719|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|General Exam|1708,1719|true|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Event|Event|General Exam|1708,1719|true|false|false|||Conjunctiva
Finding|Body Substance|General Exam|1708,1719|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|General Exam|1708,1719|true|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|General Exam|1708,1719|true|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Event|Event|General Exam|1735,1741|true|false|false|||pallor
Finding|Finding|General Exam|1735,1741|true|false|false|C0241137|Pallor of skin|pallor
Event|Event|General Exam|1745,1753|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|1745,1753|true|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|General Exam|1761,1765|true|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|General Exam|1761,1765|true|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|General Exam|1761,1765|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|General Exam|1761,1765|true|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|General Exam|1761,1772|true|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|General Exam|1766,1772|true|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|General Exam|1766,1772|true|false|false|C1561514||mucosa
Event|Event|General Exam|1777,1788|true|false|false|||xanthalesma
Anatomy|Body Location or Region|General Exam|1790,1794|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|1790,1794|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|1790,1794|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|1796,1799|false|false|false|||JVD
Finding|Finding|General Exam|1796,1799|false|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Space or Junction|General Exam|1803,1820|false|false|false|C0222753|Structure of angle of mandible|angle of mandible
Anatomy|Body Part, Organ, or Organ Component|General Exam|1812,1820|false|false|false|C0024687;C4299125|Head>Mandible;Mandible|mandible
Disorder|Neoplastic Process|General Exam|1812,1820|false|false|false|C0153511|Malignant neoplasm of mandible|mandible
Anatomy|Body Part, Organ, or Organ Component|General Exam|1821,1828|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|1821,1828|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|1852,1859|true|false|false|||murmurs
Finding|Finding|General Exam|1852,1859|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|1861,1865|true|false|false|||rubs
Finding|Finding|General Exam|1861,1865|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|1869,1876|true|false|false|||gallops
Event|Event|General Exam|1882,1889|true|false|false|||thrills
Finding|Finding|General Exam|1882,1889|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Event|Event|General Exam|1891,1896|true|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|General Exam|1898,1903|false|false|false|C0024109|Lung|LUNGS
Disorder|Acquired Abnormality|General Exam|1905,1913|false|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|Kyphosis
Disorder|Anatomical Abnormality|General Exam|1905,1913|false|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|Kyphosis
Disorder|Congenital Abnormality|General Exam|1905,1913|false|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|Kyphosis
Event|Event|General Exam|1905,1913|false|false|false|||Kyphosis
Finding|Finding|General Exam|1905,1913|false|false|false|C2115817|kyphosis|Kyphosis
Attribute|Clinical Attribute|General Exam|1915,1919|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|1915,1919|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|General Exam|1915,1919|false|false|false|||Resp
Event|Event|General Exam|1925,1932|false|false|false|||labored
Finding|Intellectual Product|General Exam|1934,1938|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Gene or Genome|General Exam|1939,1942|false|false|false|C1417055|MBNL1 gene|exp
Event|Event|General Exam|1943,1950|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|1943,1950|false|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|1965,1972|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|1965,1972|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|1965,1972|true|false|false|||ABDOMEN
Finding|Finding|General Exam|1965,1972|true|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|1974,1978|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|1974,1978|true|false|false|||Soft
Event|Event|General Exam|1996,2005|true|false|false|||distended
Finding|Finding|General Exam|1996,2005|true|false|false|C0700124|Dilated|distended
Anatomy|Body Location or Region|General Exam|2007,2010|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|2007,2010|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Part, Organ, or Organ Component|General Exam|2011,2016|true|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|2011,2016|true|false|false|C0869784|Procedure on aorta|aorta
Event|Event|General Exam|2021,2029|true|false|false|||enlarged
Procedure|Therapeutic or Preventive Procedure|General Exam|2021,2029|true|true|false|C1293134|Enlargement procedure|enlarged
Event|Event|General Exam|2034,2043|true|false|false|||palpation
Procedure|Diagnostic Procedure|General Exam|2034,2043|true|false|false|C0030247|Palpation|palpation
Anatomy|Body Location or Region|General Exam|2048,2057|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|General Exam|2048,2064|true|false|false|C0221755|Abdominal bruit|abdominal bruits
Event|Event|General Exam|2058,2064|true|false|false|||bruits
Finding|Finding|General Exam|2058,2064|true|false|false|C0006318|Bruit|bruits
Anatomy|Body Part, Organ, or Organ Component|General Exam|2066,2077|true|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Disorder|Anatomical Abnormality|General Exam|2082,2090|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|2082,2090|true|false|false|||clubbing
Event|Event|General Exam|2092,2100|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|2092,2100|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|2104,2109|true|false|false|C1717255||edema
Event|Event|General Exam|2104,2109|true|false|false|||edema
Finding|Pathologic Function|General Exam|2104,2109|true|false|false|C0013604|Edema|edema
Anatomy|Body Part, Organ, or Organ Component|General Exam|2114,2121|true|false|false|C0015811|Femur|femoral
Event|Event|General Exam|2122,2128|true|false|false|||bruits
Finding|Finding|General Exam|2122,2128|true|false|false|C0006318|Bruit|bruits
Anatomy|Body System|General Exam|2130,2134|true|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|2130,2134|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|2130,2134|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|2130,2134|true|false|false|||SKIN
Finding|Body Substance|General Exam|2130,2134|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|2130,2134|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|General Exam|2139,2145|true|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|General Exam|2139,2156|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|General Exam|2146,2156|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|General Exam|2146,2156|true|false|false|||dermatitis
Event|Event|General Exam|2158,2164|true|false|false|||ulcers
Finding|Pathologic Function|General Exam|2158,2164|true|false|false|C0041582|Ulcer|ulcers
Event|Event|General Exam|2166,2171|true|false|false|||scars
Finding|Finding|General Exam|2166,2171|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|General Exam|2166,2171|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|General Exam|2176,2185|true|false|false|C0302314|Xanthoma|xanthomas
Event|Event|General Exam|2176,2185|false|false|false|||xanthomas
Event|Event|General Exam|2211,2217|false|false|false|||intact
Finding|Finding|General Exam|2211,2217|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Idea or Concept|General Exam|2219,2227|false|false|false|C0808080|Strength (attribute)|Strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|2235,2238|false|false|false|C0227192|Inferior esophageal sphincter structure|LEs
Finding|Classification|General Exam|2235,2238|false|false|false|C0023595|Lewis Blood-Group System|LEs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2243,2246|false|false|false|C1451819|Upper Esophageal Sphincter|UEs
Disorder|Neoplastic Process|General Exam|2243,2246|false|false|false|C2205345|Embryonal sarcoma of liver|UEs
Event|Event|General Exam|2260,2269|false|false|false|||sensation
Finding|Finding|General Exam|2260,2269|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2260,2269|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2260,2269|false|false|false|C2229507|sensory exam|sensation
Finding|Functional Concept|General Exam|2294,2298|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|2294,2302|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Anatomy|Body Part, Organ, or Organ Component|General Exam|2299,2302|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Drug|Amino Acid, Peptide, or Protein|General Exam|2306,2311|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2306,2311|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2306,2311|false|false|false|||light
Finding|Finding|General Exam|2306,2311|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2306,2311|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2306,2311|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2306,2311|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2306,2311|false|false|false|C0031765|Phototherapy|light
Event|Event|General Exam|2313,2318|false|false|false|||touch
Finding|Mental Process|General Exam|2313,2318|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|2313,2318|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|2313,2318|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|2320,2329|false|false|false|||Discharge
Finding|Body Substance|General Exam|2320,2329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|2320,2329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|2320,2329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|2320,2329|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|General Exam|2330,2334|false|false|false|||exam
Finding|Functional Concept|General Exam|2330,2334|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|2330,2334|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|General Exam|2336,2341|false|false|false|C0024109|Lung|Lungs
Drug|Organic Chemical|General Exam|2343,2347|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|2343,2347|false|false|false|||CTAB
Event|Event|General Exam|2358,2367|false|false|false|||unchanged
Finding|Finding|General Exam|2358,2367|false|false|false|C0442739||unchanged
Procedure|Health Care Activity|General Exam|2389,2398|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|General Exam|2399,2403|false|false|false|||Labs
Lab|Laboratory or Test Result|General Exam|2399,2403|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|General Exam|2416,2421|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2416,2421|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2416,2421|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2422,2425|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2431,2434|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2431,2434|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2431,2434|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2441,2444|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2441,2444|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2441,2444|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2441,2444|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2450,2453|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2450,2453|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2461,2464|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2461,2464|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2461,2464|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2461,2464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2461,2464|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2468,2471|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2468,2471|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2468,2471|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2468,2471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2468,2471|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2468,2471|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2477,2481|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2477,2481|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2496,2499|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2516,2521|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2516,2521|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2516,2521|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2516,2529|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2516,2529|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2516,2529|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2522,2529|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2522,2529|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2522,2529|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2522,2529|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2522,2529|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2522,2529|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2578,2582|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2578,2582|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2578,2582|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2608,2613|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2608,2613|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2608,2613|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|2617,2620|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|2617,2620|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|2617,2620|false|false|false|||CPK
Finding|Gene or Genome|General Exam|2617,2620|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|2617,2620|false|false|false|C0201973|Creatine kinase measurement|CPK
Disorder|Disease or Syndrome|General Exam|2639,2644|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2639,2644|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2639,2644|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|2671,2676|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2671,2676|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2671,2676|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|2677,2682|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|2677,2682|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|2677,2682|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|2677,2682|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|2680,2684|false|false|false|C4722362|MB-6|MB-6
Drug|Amino Acid, Peptide, or Protein|General Exam|2685,2691|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|2685,2691|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|2710,2715|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2710,2715|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2710,2715|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2710,2723|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|2716,2723|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|2716,2723|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|2716,2723|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|2716,2723|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|2716,2723|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|2716,2723|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|2716,2723|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|2716,2723|false|false|false|C0201925|Calcium measurement|Calcium
Lab|Laboratory or Test Result|General Exam|2769,2773|false|false|false|C0587081|Laboratory test finding|Labs
Disorder|Disease or Syndrome|General Exam|2786,2791|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2786,2791|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2786,2791|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2792,2795|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2800,2803|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2800,2803|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2800,2803|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2810,2813|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2810,2813|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2810,2813|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2810,2813|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2819,2822|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2819,2822|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|2830,2833|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|2830,2833|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|2830,2833|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|2830,2833|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|2830,2833|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|2837,2840|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|2837,2840|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|2837,2840|false|false|false|||MCH
Finding|Gene or Genome|General Exam|2837,2840|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|2837,2840|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|2837,2840|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|2846,2850|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|2846,2850|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2865,2868|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2885,2890|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2885,2890|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2885,2890|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2885,2898|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2885,2898|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2885,2898|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2891,2898|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2891,2898|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2891,2898|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2891,2898|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2891,2898|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2891,2898|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|2946,2950|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2946,2950|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2946,2950|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2976,2981|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2976,2981|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2976,2981|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2982,2985|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2982,2985|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2982,2985|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|2982,2985|false|false|false|||ALT
Finding|Gene or Genome|General Exam|2982,2985|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2982,2985|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2982,2985|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2982,2985|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|2989,2992|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2989,2992|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2989,2992|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2989,2992|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2989,2992|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|2989,2992|false|false|false|||AST
Finding|Gene or Genome|General Exam|2989,2992|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Disease or Syndrome|General Exam|3008,3013|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3008,3013|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3008,3013|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3025,3028|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|General Exam|3025,3028|false|false|false|C0023821|High Density Lipoproteins|HDL
Event|Event|General Exam|3025,3028|false|false|false|||HDL
Finding|Gene or Genome|General Exam|3025,3028|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|General Exam|3025,3028|false|false|false|C0392885|High density lipoprotein measurement|HDL
Disorder|Disease or Syndrome|General Exam|3070,3075|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3070,3075|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3070,3075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3077,3082|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|General Exam|3077,3082|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|General Exam|3077,3082|false|false|false|||HbA1c
Procedure|Laboratory Procedure|General Exam|3077,3082|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|General Exam|3088,3091|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|General Exam|3110,3115|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3110,3115|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3110,3115|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3119,3122|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|3119,3122|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|3119,3122|false|false|false|||CPK
Finding|Gene or Genome|General Exam|3119,3122|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|3119,3122|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|3129,3134|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3129,3134|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3129,3134|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3129,3134|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Pharmacologic Substance|General Exam|3132,3136|false|false|false|C4722362|MB-6|MB-6
Disorder|Disease or Syndrome|General Exam|3163,3168|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3163,3168|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3163,3168|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3172,3175|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|3172,3175|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|3172,3175|false|false|false|||CPK
Finding|Gene or Genome|General Exam|3172,3175|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|3172,3175|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|3182,3187|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3182,3187|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3182,3187|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3182,3187|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|General Exam|3185,3189|false|false|false|C0602256|MB 5|MB-5
Disorder|Disease or Syndrome|General Exam|3216,3221|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3216,3221|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3216,3221|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3225,3228|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|3225,3228|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|General Exam|3225,3228|false|false|false|||CPK
Finding|Gene or Genome|General Exam|3225,3228|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|3225,3228|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|General Exam|3235,3240|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3235,3240|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3235,3240|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3235,3240|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|General Exam|3238,3242|false|false|false|C0602256|MB 5|MB-5
Disorder|Disease or Syndrome|General Exam|3269,3274|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3269,3274|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3269,3274|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3322,3328|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|3322,3328|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Amino Acid, Peptide, or Protein|General Exam|3336,3339|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Hormone|General Exam|3336,3339|false|false|false|C0018064|Equine Gonadotropins|ECG
Drug|Pharmacologic Substance|General Exam|3336,3339|false|false|false|C0018064|Equine Gonadotropins|ECG
Event|Event|General Exam|3336,3339|false|false|false|||ECG
Finding|Intellectual Product|General Exam|3336,3339|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|ECG
Procedure|Diagnostic Procedure|General Exam|3336,3339|false|false|false|C1623258|Electrocardiography|ECG
Drug|Biomedical or Dental Material|General Exam|3359,3367|false|false|false|C0168634|BaseLine dental cement|Baseline
Event|Event|General Exam|3359,3367|false|false|false|||Baseline
Finding|Idea or Concept|General Exam|3359,3367|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Event|Event|General Exam|3368,3376|false|false|false|||artifact
Phenomenon|Human-caused Phenomenon or Process|General Exam|3368,3376|false|false|false|C0085089|Morphologic artifact|artifact
Anatomy|Body Space or Junction|General Exam|3378,3383|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|General Exam|3378,3383|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|General Exam|3378,3383|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|General Exam|3378,3383|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|General Exam|3378,3390|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|General Exam|3384,3390|false|false|false|||rhythm
Finding|Finding|General Exam|3384,3390|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3384,3390|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Attribute|Clinical Attribute|General Exam|3396,3408|false|false|false|C0429028;C0488414|QT interval feature (observable entity)|Q-T interval
Event|Event|General Exam|3400,3408|false|false|false|||interval
Finding|Intellectual Product|General Exam|3400,3408|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|General Exam|3417,3429|false|false|false|||milliseconds
Event|Event|General Exam|3433,3438|false|false|false|||waves
Finding|Finding|General Exam|3462,3468|false|false|false|C0429103|T wave feature|T wave
Event|Event|General Exam|3464,3468|false|false|false|||wave
Finding|Gene or Genome|General Exam|3464,3468|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|General Exam|3464,3468|false|false|false|C0678544||wave
Disorder|Congenital Abnormality|General Exam|3470,3483|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|3470,3483|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|3470,3483|false|false|false|C0000769|teratologic|abnormalities
Anatomy|Body Location or Region|General Exam|3497,3504|false|false|false|C0449220|Lead site V6|lead V6
Event|Event|General Exam|3506,3514|false|false|false|||Consider
Disorder|Disease or Syndrome|General Exam|3521,3529|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|General Exam|3521,3529|false|false|false|||anterior
Anatomy|Tissue|General Exam|3531,3541|false|false|false|C0027061|Myocardium|myocardial
Attribute|Clinical Attribute|General Exam|3531,3552|false|false|false|C2926063||myocardial infarction
Disorder|Disease or Syndrome|General Exam|3531,3552|false|false|false|C0027051|Myocardial Infarction|myocardial infarction
Event|Event|General Exam|3542,3552|false|false|false|||infarction
Finding|Pathologic Function|General Exam|3542,3552|false|false|false|C0021308|Infarction|infarction
Event|Event|General Exam|3573,3580|false|false|false|||tracing
Anatomy|Body Part, Organ, or Organ Component|General Exam|3589,3595|true|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|General Exam|3589,3611|true|false|false|C0033036|Atrial Premature Complexes|atrial premature beats
Finding|Finding|General Exam|3596,3605|true|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Finding|Pathologic Function|General Exam|3596,3605|true|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Disorder|Disease or Syndrome|General Exam|3596,3611|true|false|false|C0340464|Premature Cardiac Complex|premature beats
Event|Event|General Exam|3606,3611|true|false|false|||beats
Event|Event|General Exam|3620,3624|true|false|false|||seen
Attribute|Clinical Attribute|General Exam|3630,3642|false|false|false|C0429028;C0488414|QT interval feature (observable entity)|Q-T interval
Event|Event|General Exam|3634,3642|false|false|false|||interval
Finding|Intellectual Product|General Exam|3634,3642|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|General Exam|3647,3654|false|false|false|||shorter
Finding|Finding|General Exam|3659,3665|false|false|false|C0429103|T wave feature|T wave
Finding|Gene or Genome|General Exam|3661,3665|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|General Exam|3661,3665|false|false|false|C0678544||wave
Disorder|Congenital Abnormality|General Exam|3666,3679|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|General Exam|3666,3679|false|false|false|||abnormalities
Finding|Functional Concept|General Exam|3666,3679|false|false|false|C0000769|teratologic|abnormalities
Event|Event|General Exam|3689,3698|false|false|false|||prominent
Event|Event|General Exam|3704,3707|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|3704,3707|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|3728,3733|false|false|false|||views
Anatomy|Body Location or Region|General Exam|3741,3746|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|3741,3746|false|false|false|C0741025|Chest problem|chest
Event|Event|General Exam|3747,3758|false|false|false|||demonstrate
Finding|Finding|General Exam|3759,3762|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|3759,3762|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Location or Region|General Exam|3763,3767|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|3763,3767|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|3763,3767|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|3763,3767|false|false|false|C0740941|Lung Problem|lung
Finding|Organ or Tissue Function|General Exam|3763,3775|false|false|false|C0231953|Lung Volumes|lung volumes
Event|Event|General Exam|3768,3775|false|false|false|||volumes
Anatomy|Tissue|General Exam|3793,3800|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|3793,3800|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|3793,3810|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|General Exam|3801,3810|false|false|false|||effusions
Finding|Pathologic Function|General Exam|3801,3810|false|false|false|C0013687|effusion|effusions
Event|Event|General Exam|3815,3818|false|false|false|||new
Finding|Finding|General Exam|3815,3818|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|3815,3818|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|General Exam|3834,3839|true|false|false|||signs
Finding|Finding|General Exam|3834,3839|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|General Exam|3834,3839|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|General Exam|3843,3852|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|General Exam|3843,3852|true|false|false|||pneumonia
Anatomy|Body Part, Organ, or Organ Component|General Exam|3856,3865|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|3856,3865|true|false|false|C2707265||pulmonary
Finding|Finding|General Exam|3856,3865|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|General Exam|3856,3885|true|false|false|C5849517|Pulmonary vascular congestion|pulmonary vascular congestion
Anatomy|Body Part, Organ, or Organ Component|General Exam|3866,3874|true|false|false|C0005847|Blood Vessel|vascular
Event|Event|General Exam|3875,3885|false|false|false|||congestion
Finding|Pathologic Function|General Exam|3875,3885|false|false|false|C0700148|Congestion|congestion
Anatomy|Body Part, Organ, or Organ Component|General Exam|3887,3892|false|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|General Exam|3887,3892|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Event|Event|General Exam|3887,3892|false|false|false|||Heart
Finding|Sign or Symptom|General Exam|3887,3892|false|false|false|C0795691|HEART PROBLEM|Heart
Event|Event|General Exam|3901,3907|false|false|false|||normal
Event|Event|General Exam|3931,3937|false|false|false|||stable
Finding|Intellectual Product|General Exam|3931,3937|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|General Exam|3939,3944|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|Aorta
Procedure|Health Care Activity|General Exam|3939,3944|false|false|false|C0869784|Procedure on aorta|Aorta
Event|Event|General Exam|3958,3966|false|false|false|||tortuous
Finding|Finding|General Exam|3958,3966|false|false|false|C4068863|Tortuous|tortuous
Event|Event|General Exam|3968,3977|false|false|false|||unchanged
Finding|Finding|General Exam|3968,3977|false|false|false|C0442739||unchanged
Anatomy|Body Part, Organ, or Organ Component|General Exam|3979,3985|false|false|false|C0003483|Aorta|Aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|3979,3990|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|Aortic arch
Disorder|Anatomical Abnormality|General Exam|3979,3990|false|false|false|C4759703|Aortic arch malformation|Aortic arch
Finding|Pathologic Function|General Exam|3979,4005|false|false|false|C1969291|Aortic arch calcification|Aortic arch calcifications
Anatomy|Body Location or Region|General Exam|3986,3990|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|3986,3990|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|3986,3990|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|3986,3990|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|3986,3990|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|General Exam|3991,4005|false|false|false|||calcifications
Finding|Finding|General Exam|3991,4005|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|General Exam|3991,4005|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Event|Event|General Exam|4010,4014|false|false|false|||seen
Disorder|Disease or Syndrome|General Exam|4029,4041|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|General Exam|4029,4041|true|false|false|||pneumothorax
Disorder|Disease or Syndrome|General Exam|4052,4065|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|4052,4065|true|false|false|||consolidation
Event|Event|General Exam|4077,4083|false|false|false|||imaged
Anatomy|Body Location or Region|General Exam|4085,4098|false|false|false|C0230165;C2937240|Upper abdomen (surface region);Upper abdomen structure|upper abdomen
Anatomy|Body Part, Organ, or Organ Component|General Exam|4085,4098|false|false|false|C0230165;C2937240|Upper abdomen (surface region);Upper abdomen structure|upper abdomen
Anatomy|Body Location or Region|General Exam|4091,4098|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|4091,4098|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|General Exam|4091,4098|false|false|false|||abdomen
Finding|Finding|General Exam|4091,4098|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|General Exam|4102,4114|false|false|false|||unremarkable
Event|Event|General Exam|4116,4126|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|4116,4126|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|4116,4126|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Anatomy|Tissue|General Exam|4133,4140|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|4133,4140|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|General Exam|4133,4150|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|General Exam|4141,4150|false|false|false|||effusions
Finding|Pathologic Function|General Exam|4141,4150|false|false|false|C0013687|effusion|effusions
Event|Event|General Exam|4152,4155|false|false|false|||new
Finding|Finding|General Exam|4152,4155|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|4152,4155|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|General Exam|4167,4179|false|false|false|||unremarkable
Event|Event|General Exam|4182,4186|false|false|false|||ECHO
Procedure|Health Care Activity|General Exam|4182,4186|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|General Exam|4182,4186|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|General Exam|4196,4200|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4196,4207|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|General Exam|4201,4207|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|General Exam|4218,4225|false|false|false|||dilated
Finding|Functional Concept|General Exam|4241,4246|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4247,4253|false|false|false|C0018792|Heart Atrium|atrial
Event|Event|General Exam|4255,4263|false|false|false|||pressure
Finding|Finding|General Exam|4255,4263|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|4255,4263|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|4255,4263|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|4255,4263|false|false|false|C0033095||pressure
Finding|Functional Concept|General Exam|4277,4281|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4277,4298|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|4282,4293|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|4282,4298|false|false|false|C0507618|Wall of ventricle|ventricular wall
Finding|Finding|General Exam|4282,4308|false|false|false|C2024242|cardiac evaluation of ventricular wall thickness|ventricular wall thickness
Event|Event|General Exam|4299,4308|false|false|false|||thickness
Anatomy|Body Space or Junction|General Exam|4310,4316|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|4310,4316|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|4310,4316|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|General Exam|4318,4322|false|false|false|||size
Finding|Organ or Tissue Function|General Exam|4343,4351|false|false|false|C0039155|Systole|systolic
Event|Event|General Exam|4352,4360|false|false|false|||function
Finding|Finding|General Exam|4352,4360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|4352,4360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|4352,4360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|4352,4360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|General Exam|4365,4371|false|false|false|||normal
Attribute|Clinical Attribute|General Exam|4373,4377|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|General Exam|4373,4377|false|false|false|||LVEF
Procedure|Diagnostic Procedure|General Exam|4373,4377|false|false|false|C3837267|LVEF (procedure)|LVEF
Finding|Functional Concept|General Exam|4386,4391|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|4392,4403|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|4404,4411|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|General Exam|4421,4425|false|false|false|||free
Finding|Functional Concept|General Exam|4421,4425|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|General Exam|4426,4437|false|false|false|C1980023|Wall motion|wall motion
Event|Event|General Exam|4431,4437|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|General Exam|4431,4437|false|false|false|C0026597|Motion|motion
Event|Event|General Exam|4443,4449|false|false|false|||normal
Event|Event|General Exam|4455,4464|false|false|false|||diameters
Anatomy|Body Part, Organ, or Organ Component|General Exam|4468,4473|false|false|false|C0003483;C4037978|Aorta;Chest+Abdomen>Aorta|aorta
Procedure|Health Care Activity|General Exam|4468,4473|false|false|false|C0869784|Procedure on aorta|aorta
Anatomy|Body Space or Junction|General Exam|4481,4486|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|General Exam|4481,4486|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|General Exam|4481,4486|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|General Exam|4481,4486|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|General Exam|4488,4497|false|false|false|||ascending
Finding|Functional Concept|General Exam|4488,4497|false|false|false|C1547175;C1962987|Ascend (action);Sequencing - Ascending|ascending
Anatomy|Body Location or Region|General Exam|4502,4506|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|4502,4506|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|4502,4506|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|4502,4506|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|4502,4506|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|General Exam|4508,4514|false|false|false|||levels
Event|Event|General Exam|4519,4525|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|4531,4537|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4531,4543|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|4538,4543|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|4544,4552|false|false|false|||leaflets
Event|Event|General Exam|4569,4578|false|false|false|||thickened
Anatomy|Body Part, Organ, or Organ Component|General Exam|4583,4589|true|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|General Exam|4583,4598|true|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|General Exam|4590,4598|true|false|false|||stenosis
Finding|Pathologic Function|General Exam|4590,4598|true|false|false|C1261287|Stenosis|stenosis
Event|Event|General Exam|4606,4613|true|false|false|||present
Finding|Finding|General Exam|4606,4613|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|4606,4613|true|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|General Exam|4618,4624|true|false|false|||masses
Disorder|Anatomical Abnormality|General Exam|4629,4640|true|false|false|C1285498|Vegetation|vegetations
Event|Event|General Exam|4629,4640|true|false|false|||vegetations
Event|Event|General Exam|4645,4649|true|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|General Exam|4657,4663|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4657,4669|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|4664,4669|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|4692,4700|true|false|false|||excluded
Finding|Finding|General Exam|4708,4724|true|false|false|C2828075|Suboptimal Image Reason|suboptimal image
Disorder|Disease or Syndrome|General Exam|4719,4724|true|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|General Exam|4719,4724|true|false|false|||image
Finding|Intellectual Product|General Exam|4719,4724|true|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Finding|Functional Concept|General Exam|4734,4739|false|false|false|C1883002|Sequence Chromatogram|Trace
Anatomy|Body Part, Organ, or Organ Component|General Exam|4740,4746|false|false|false|C0003483|Aorta|aortic
Event|Event|General Exam|4748,4761|false|false|false|||regurgitation
Finding|Finding|General Exam|4748,4761|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4748,4761|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4748,4761|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4765,4769|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|General Exam|4775,4787|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|4782,4787|false|false|false|C1186983|Anatomical valve|valve
Event|Event|General Exam|4788,4796|false|false|false|||leaflets
Event|Event|General Exam|4815,4821|false|false|false|||normal
Event|Event|General Exam|4848,4856|false|false|false|||directed
Disorder|Disease or Syndrome|General Exam|4857,4860|false|false|false|C0039235|Tachycardia, Ectopic Junctional|jet
Event|Event|General Exam|4857,4860|false|false|false|||jet
Finding|Gene or Genome|General Exam|4857,4860|false|false|false|C1539482|FBXL15 gene|jet
Event|Event|General Exam|4865,4869|false|false|false|||mild
Finding|Intellectual Product|General Exam|4865,4869|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|General Exam|4873,4881|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4873,4881|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|General Exam|4888,4908|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|4895,4908|false|false|false|||regurgitation
Finding|Finding|General Exam|4895,4908|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4895,4908|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4895,4908|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4912,4916|false|false|false|||seen
Finding|Finding|General Exam|4918,4926|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|4918,4926|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|General Exam|4933,4956|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|General Exam|4943,4956|false|false|false|||regurgitation
Finding|Finding|General Exam|4943,4956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|4943,4956|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|4943,4956|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|4960,4964|false|false|false|||seen
Event|Event|General Exam|4975,4983|false|false|false|||moderate
Finding|Finding|General Exam|4975,4983|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|4975,4983|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Body Part, Organ, or Organ Component|General Exam|4985,4994|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|4985,4994|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|4985,4994|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|4985,5001|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|4995,5001|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|4995,5001|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|5002,5010|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|General Exam|5002,5023|false|false|false|C0221155|Systolic Hypertension|systolic hypertension
Disorder|Disease or Syndrome|General Exam|5011,5023|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|5011,5023|false|false|false|||hypertension
Drug|Amino Acid, Peptide, or Protein|General Exam|5029,5032|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|General Exam|5029,5032|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|General Exam|5029,5032|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|General Exam|5029,5032|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Attribute|Clinical Attribute|General Exam|5029,5042|false|false|false|C0442709|end diastolic|end-diastolic
Attribute|Clinical Attribute|General Exam|5033,5042|false|false|false|C0012000|Diastole|diastolic
Event|Event|General Exam|5033,5042|false|false|false|||diastolic
Finding|Pathologic Function|General Exam|5044,5066|false|false|false|C0034088|Pulmonary Valve Insufficiency|pulmonic regurgitation
Event|Event|General Exam|5053,5066|false|false|false|||regurgitation
Finding|Finding|General Exam|5053,5066|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5053,5066|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5053,5066|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|5079,5088|false|false|false|||increased
Event|Event|General Exam|5089,5099|false|false|false|||suggesting
Anatomy|Body Part, Organ, or Organ Component|General Exam|5101,5110|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|5101,5110|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|5101,5110|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5101,5117|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|5111,5117|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5111,5117|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Attribute|Clinical Attribute|General Exam|5118,5127|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|General Exam|5118,5140|false|false|false|C0235222|Diastolic hypertension|diastolic hypertension
Disorder|Disease or Syndrome|General Exam|5128,5140|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|5128,5140|false|false|false|||hypertension
Disorder|Disease or Syndrome|General Exam|5154,5162|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|General Exam|5154,5162|false|false|false|||anterior
Phenomenon|Natural Phenomenon or Process|General Exam|5164,5169|false|false|false|C0282173|Space (Astronomy)|space
Finding|Idea or Concept|General Exam|5176,5187|false|false|false|C0750501|most likely|most likely
Finding|Finding|General Exam|5181,5187|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5181,5187|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|5188,5198|false|false|false|||represents
Anatomy|Tissue|General Exam|5211,5214|false|false|false|C0001527|Adipose tissue|fat
Drug|Amino Acid, Peptide, or Protein|General Exam|5211,5214|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Biologically Active Substance|General Exam|5211,5214|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Organic Chemical|General Exam|5211,5214|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Drug|Pharmacologic Substance|General Exam|5211,5214|false|false|false|C0015677;C1435181;C3887682|FAT1 protein, human;Fatty acid glycerol esters;Platelet Glycoprotein 4, human|fat
Finding|Gene or Genome|General Exam|5211,5214|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Finding|Receptor|General Exam|5211,5214|false|false|false|C0812278;C1366645;C1705088;C1708004;C3887682|CD36 gene;CD36 wt Allele;FAT1 gene;FAT1 wt Allele;Platelet Glycoprotein 4, human|fat
Procedure|Therapeutic or Preventive Procedure|General Exam|5211,5214|false|false|false|C0279453|doxorubicin/fluorouracil/triazinate protocol|fat
Anatomy|Tissue|General Exam|5211,5218|false|false|false|C0935625|Fat pad|fat pad
Anatomy|Anatomical Structure|General Exam|5215,5218|false|false|false|C3669270|Strucure of thick cushion of skin|pad
Disorder|Disease or Syndrome|General Exam|5215,5218|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Disorder|Neoplastic Process|General Exam|5215,5218|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Drug|Biomedical or Dental Material|General Exam|5215,5218|false|false|false|C2347441|Pad Dosage Form|pad
Event|Event|General Exam|5215,5218|false|false|false|||pad
Finding|Gene or Genome|General Exam|5215,5218|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|pad
Procedure|Therapeutic or Preventive Procedure|General Exam|5215,5218|false|false|false|C3814046|PAD Regimen|pad
Event|Event|General Exam|5220,5230|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|5220,5230|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|5220,5230|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Finding|General Exam|5232,5248|false|false|false|C2828075|Suboptimal Image Reason|Suboptimal image
Disorder|Disease or Syndrome|General Exam|5243,5248|false|false|false|C1846009|Intrauterine growth restriction, metaphyseal dysplasia, adrenal hypoplasia congenita, and genital anomaly syndrome|image
Event|Event|General Exam|5243,5248|false|false|false|||image
Finding|Intellectual Product|General Exam|5243,5248|false|false|false|C1696103;C1704254;C1704922;C3542466|Image;Image (foundation metadata concept);Medical Image;image - dosage form|image
Event|Event|General Exam|5249,5256|false|false|false|||quality
Anatomy|Body Space or Junction|General Exam|5280,5286|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|5280,5286|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5280,5286|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|General Exam|5287,5292|false|false|false|||sizes
Procedure|Laboratory Procedure|General Exam|5298,5307|false|false|false|C0033085|Biologic Preservation|preserved
Finding|Organ or Tissue Function|General Exam|5343,5351|false|false|false|C0039155|Systole|systolic
Event|Event|General Exam|5352,5360|false|false|false|||function
Finding|Finding|General Exam|5352,5360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|5352,5360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|5352,5360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|5352,5360|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Anatomy|Body Part, Organ, or Organ Component|General Exam|5362,5371|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|General Exam|5362,5371|false|false|false|C2707265||Pulmonary
Finding|Finding|General Exam|5362,5371|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5362,5378|false|false|false|C0034052|Pulmonary artery structure|Pulmonary artery
Disorder|Disease or Syndrome|General Exam|5362,5391|false|false|false|C2973725|Pulmonary arterial hypertension|Pulmonary artery hypertension
Anatomy|Body Part, Organ, or Organ Component|General Exam|5372,5378|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5372,5378|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|General Exam|5379,5391|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|5379,5391|false|false|false|||hypertension
Finding|Intellectual Product|General Exam|5393,5397|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|General Exam|5398,5406|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|5398,5406|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|General Exam|5408,5428|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|General Exam|5415,5428|false|false|false|||regurgitation
Finding|Finding|General Exam|5415,5428|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5415,5428|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5415,5428|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Finding|General Exam|5430,5438|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|General Exam|5430,5438|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Finding|General Exam|5430,5462|false|false|false|C3276922|Tricuspid regurgitation, moderate|Moderate tricuspid regurgitation
Disorder|Disease or Syndrome|General Exam|5439,5462|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|General Exam|5449,5462|false|false|false|||regurgitation
Finding|Finding|General Exam|5449,5462|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5449,5462|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5449,5462|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|5489,5494|false|false|false|||study
Finding|Intellectual Product|General Exam|5489,5494|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|General Exam|5489,5494|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Event|Event|General Exam|5503,5511|false|false|false|||reviewed
Event|Event|General Exam|5526,5534|false|false|false|||severity
Disorder|Disease or Syndrome|General Exam|5549,5572|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|General Exam|5559,5572|false|false|false|||regurgitation
Finding|Finding|General Exam|5559,5572|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5559,5572|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5559,5572|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|General Exam|5577,5586|false|false|false|||increased
Finding|Finding|General Exam|5592,5600|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|5592,5600|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|General Exam|5604,5616|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|General Exam|5604,5616|false|false|false|||hypertension
Event|Event|General Exam|5624,5634|false|false|false|||identified
Event|Event|Hospital Course|5665,5670|false|false|false|||woman
Disorder|Disease or Syndrome|Hospital Course|5680,5692|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|5680,5692|false|false|false|||hypertension
Event|Event|Hospital Course|5694,5707|false|false|false|||hypelipidemia
Disorder|Disease or Syndrome|Hospital Course|5709,5717|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|Hospital Course|5709,5717|false|false|false|||diabetes
Event|Event|Hospital Course|5719,5727|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5731,5738|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|5731,5738|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|5731,5738|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|5731,5738|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|5731,5738|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|5731,5738|false|false|false|C0202098|Insulin measurement|insulin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5740,5750|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5751,5760|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Hospital Course|5761,5767|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|5761,5767|false|false|false|||stroke
Finding|Finding|Hospital Course|5761,5767|false|false|false|C5977286|Stroke (heart beat)|stroke
Attribute|Clinical Attribute|Hospital Course|5777,5782|false|false|false|C1300072|Tumor stage|stage
Disorder|Disease or Syndrome|Hospital Course|5787,5790|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|Hospital Course|5787,5790|false|false|false|||CKD
Event|Event|Hospital Course|5810,5820|false|false|false|||presenting
Event|Event|Hospital Course|5826,5833|false|false|false|||fatigue
Finding|Sign or Symptom|Hospital Course|5826,5833|false|false|false|C0015672|Fatigue|fatigue
Event|Event|Hospital Course|5839,5842|false|false|false|||DOE
Finding|Sign or Symptom|Hospital Course|5839,5842|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|Hospital Course|5869,5874|false|false|false|||worse
Finding|Finding|Hospital Course|5869,5874|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Hospital Course|5869,5874|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Event|Hospital Course|5890,5899|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5890,5899|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|5906,5913|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5906,5913|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5906,5913|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|5906,5917|false|false|false|C0332310|Has patient|patient has
Event|Event|Hospital Course|5918,5923|false|false|false|||known
Attribute|Clinical Attribute|Hospital Course|5924,5933|false|false|false|C0012000|Diastole|diastolic
Finding|Pathologic Function|Hospital Course|5924,5945|false|false|false|C0520863|Diastolic dysfunction|diastolic dysfunction
Disorder|Disease or Syndrome|Hospital Course|5934,5945|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|5934,5945|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|5934,5945|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|5934,5945|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|5934,5945|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|Hospital Course|5970,5982|false|false|false|||noncompliant
Attribute|Clinical Attribute|Hospital Course|5992,6003|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5992,6003|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|5992,6003|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|5992,6003|false|false|false|C4284232|Medications|medications
Finding|Finding|Hospital Course|6004,6011|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|6007,6011|false|false|false|||home
Finding|Idea or Concept|Hospital Course|6007,6011|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6007,6011|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6007,6011|false|false|false|C1553498|home health encounter|home
Event|Activity|Hospital Course|6016,6023|false|false|false|C1706079||arrival
Event|Event|Hospital Course|6016,6023|false|false|false|||arrival
Finding|Functional Concept|Hospital Course|6016,6023|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|Hospital Course|6032,6037|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|6043,6051|false|false|false|||required
Drug|Organic Chemical|Hospital Course|6052,6063|false|false|false|C0020223|hydralazine|hydralazine
Drug|Pharmacologic Substance|Hospital Course|6052,6063|false|false|false|C0020223|hydralazine|hydralazine
Event|Event|Hospital Course|6052,6063|false|false|false|||hydralazine
Event|Event|Hospital Course|6073,6078|false|false|false|||bring
Finding|Finding|Hospital Course|6101,6107|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6101,6107|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|6121,6124|false|true|false|C1849718|POPLITEAL PTERYGIUM SYNDROME, LETHAL TYPE|BPs
Drug|Organic Chemical|Hospital Course|6121,6124|false|true|false|C2740858|BPS|BPs
Drug|Pharmacologic Substance|Hospital Course|6121,6124|false|true|false|C2740858|BPS|BPs
Event|Event|Hospital Course|6121,6124|false|false|false|||BPs
Finding|Finding|Hospital Course|6125,6132|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|6128,6132|false|false|false|||home
Finding|Idea or Concept|Hospital Course|6128,6132|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6128,6132|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6128,6132|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|6156,6168|false|false|false|||contributing
Event|Event|Hospital Course|6176,6179|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|6176,6179|false|false|false|C0013404|Dyspnea|SOB
Anatomy|Body Space or Junction|Hospital Course|6181,6184|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|6181,6184|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|6185,6197|false|false|false|||exacerbation
Finding|Finding|Hospital Course|6185,6197|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Neoplastic Process|Hospital Course|6203,6212|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|6203,6212|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|Hospital Course|6213,6219|false|false|false|||demand
Finding|Idea or Concept|Hospital Course|6213,6219|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6213,6219|false|false|false|C0441516|Demand (clinical)|demand
Event|Event|Hospital Course|6221,6232|false|false|false|||myonecrosis
Finding|Pathologic Function|Hospital Course|6221,6232|false|false|false|C0235957|Muscle necrosis|myonecrosis
Finding|Finding|Hospital Course|6234,6246|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Disorder|Disease or Syndrome|Hospital Course|6234,6254|false|false|false|C0745138|Hypertensive Urgency|hypertensive urgency
Event|Event|Hospital Course|6247,6254|false|false|false|||urgency
Event|Event|Hospital Course|6268,6276|false|false|false|||elevated
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6278,6286|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|6278,6286|false|false|false|C0041199|Troponin|troponin
Event|Event|Hospital Course|6278,6286|false|false|false|||troponin
Procedure|Laboratory Procedure|Hospital Course|6278,6286|false|false|false|C0523952|Troponin measurement|troponin
Disorder|Disease or Syndrome|Hospital Course|6291,6294|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6291,6294|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|6291,6294|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|6291,6294|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|6291,6294|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|6291,6294|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|6291,6294|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6291,6294|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|6340,6352|true|false|false|||presentation
Finding|Idea or Concept|Hospital Course|6340,6352|true|false|false|C0449450|Presentation|presentation
Finding|Body Substance|Hospital Course|6355,6362|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6355,6362|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6355,6362|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|6355,6366|false|false|false|C0332310|Has patient|patient has
Finding|Idea or Concept|Hospital Course|6375,6379|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|Hospital Course|6375,6387|false|false|false|C1830376||risk factors
Finding|Finding|Hospital Course|6375,6387|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|Hospital Course|6375,6387|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|Hospital Course|6380,6387|false|false|false|||factors
Finding|Intellectual Product|Hospital Course|6392,6397|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|6392,6415|false|false|false|C0948089|Acute Coronary Syndrome|acute coronary syndrome
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6398,6406|false|false|false|C0018787|Heart|coronary
Disorder|Disease or Syndrome|Hospital Course|6407,6415|false|false|false|C0039082|Syndrome|syndrome
Event|Event|Hospital Course|6407,6415|false|false|false|||syndrome
Attribute|Clinical Attribute|Hospital Course|6427,6434|false|false|false|C3854129||symptom
Event|Event|Hospital Course|6427,6434|false|false|false|||symptom
Finding|Sign or Symptom|Hospital Course|6427,6434|false|false|false|C1457887|Symptoms|symptom
Event|Event|Hospital Course|6439,6442|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|6439,6442|false|false|false|C0013404|Dyspnea|SOB
Finding|Mental Process|Hospital Course|6450,6457|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|6470,6473|false|false|false|C1849718|POPLITEAL PTERYGIUM SYNDROME, LETHAL TYPE|BPs
Drug|Organic Chemical|Hospital Course|6470,6473|false|false|false|C2740858|BPS|BPs
Drug|Pharmacologic Substance|Hospital Course|6470,6473|false|false|false|C2740858|BPS|BPs
Event|Event|Hospital Course|6470,6473|false|false|false|||BPs
Event|Event|Hospital Course|6475,6485|false|false|false|||attributed
Drug|Pharmacologic Substance|Hospital Course|6489,6499|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|6489,6499|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|6489,6499|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Hospital Course|6489,6513|false|false|false|C0746935|Medication Nonadherence|medication noncompliance
Event|Event|Hospital Course|6500,6513|false|false|false|||noncompliance
Finding|Finding|Hospital Course|6514,6521|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|6517,6521|false|false|false|||home
Finding|Idea or Concept|Hospital Course|6517,6521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6517,6521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6517,6521|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6527,6535|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|6527,6535|false|false|false|C0041199|Troponin|troponin
Event|Event|Hospital Course|6527,6535|false|false|false|||troponin
Procedure|Laboratory Procedure|Hospital Course|6527,6535|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|Hospital Course|6537,6541|false|false|false|||fell
Finding|Finding|Hospital Course|6552,6564|false|false|false|C4533677|at admission|at admission
Event|Event|Hospital Course|6555,6564|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|6555,6564|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|6576,6585|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6576,6585|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6576,6585|false|false|false|C0030685|Patient Discharge|discharge
Finding|Mental Process|Hospital Course|6593,6600|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6605,6610|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|6605,6610|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|6605,6622|false|false|false|C1565489|Renal Insufficiency|renal dysfunction
Finding|Finding|Hospital Course|6605,6622|false|false|false|C3279454|Renal dysfunction|renal dysfunction
Disorder|Disease or Syndrome|Hospital Course|6611,6622|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|6611,6622|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|6611,6622|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|6611,6622|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|6611,6622|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Idea or Concept|Hospital Course|6644,6649|true|false|false|C1550016|Remote control command - Clear|clear
Drug|Organic Chemical|Hospital Course|6650,6654|true|false|false|C0246719|risedronate|rise
Drug|Pharmacologic Substance|Hospital Course|6650,6654|true|false|false|C0246719|risedronate|rise
Event|Event|Hospital Course|6650,6654|true|false|false|||rise
Finding|Intellectual Product|Hospital Course|6650,6654|true|false|false|C4321377|Relational and Item-Specific Encoding Task|rise
Event|Event|Hospital Course|6659,6663|true|false|false|||fall
Finding|Finding|Hospital Course|6659,6663|true|false|false|C0085639|Falls|fall
Finding|Intellectual Product|Hospital Course|6679,6684|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Hospital Course|6685,6695|false|false|false|||infarction
Finding|Pathologic Function|Hospital Course|6685,6695|false|false|false|C0021308|Infarction|infarction
Anatomy|Tissue|Hospital Course|6701,6707|false|false|false|C4316797|Plaque Tissue|plaque
Disorder|Acquired Abnormality|Hospital Course|6701,6707|false|false|false|C0011389;C0333463|Dental Plaque;Senile Plaques|plaque
Disorder|Disease or Syndrome|Hospital Course|6701,6707|false|false|false|C0011389;C0333463|Dental Plaque;Senile Plaques|plaque
Finding|Finding|Hospital Course|6701,6707|false|false|false|C0241148;C0332461|Cutaneous plaque;Plaque (lesion)|plaque
Disorder|Injury or Poisoning|Hospital Course|6708,6715|false|false|false|C3203359|Rupture|rupture
Event|Event|Hospital Course|6708,6715|false|false|false|||rupture
Event|Event|Hospital Course|6720,6730|false|false|false|||thrombosis
Finding|Pathologic Function|Hospital Course|6720,6730|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|Hospital Course|6741,6750|false|false|false|||scheduled
Finding|Classification|Hospital Course|6758,6768|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|6758,6768|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Attribute|Clinical Attribute|Hospital Course|6769,6775|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|6769,6775|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|6769,6775|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|6769,6775|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|6769,6780|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Hospital Course|6776,6780|false|false|false|C4318744|Test - temporal region|test
Event|Event|Hospital Course|6776,6780|false|false|false|||test
Finding|Functional Concept|Hospital Course|6776,6780|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|6776,6780|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|6776,6780|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|6776,6780|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Hospital Course|6784,6792|false|false|false|||evaluate
Event|Event|Hospital Course|6798,6806|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|6798,6806|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|6798,6809|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Hospital Course|6810,6818|false|false|false|||ischemia
Finding|Pathologic Function|Hospital Course|6810,6818|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6810,6818|false|false|false|C4321499|Ischemia Procedure|ischemia
Phenomenon|Natural Phenomenon or Process|Hospital Course|6824,6828|false|false|false|C0806140|Flow|flow
Disorder|Disease or Syndrome|Hospital Course|6838,6841|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6838,6841|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|6838,6841|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|6838,6841|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|6838,6841|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|6838,6841|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|6838,6841|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6838,6841|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|6846,6855|false|false|false|||decreased
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6856,6859|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|6856,6859|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|6856,6859|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|6856,6859|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Hospital Course|6856,6859|false|false|false|||ASA
Finding|Gene or Genome|Hospital Course|6856,6859|false|false|false|C1412553|ARSA gene|ASA
Event|Event|Hospital Course|6891,6899|false|false|false|||decrease
Event|Event|Hospital Course|6904,6908|false|false|false|||risk
Finding|Idea or Concept|Hospital Course|6904,6908|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|Hospital Course|6904,6911|false|false|true|C0035647|Risk|risk of
Finding|Finding|Hospital Course|6904,6920|false|false|false|C3251812|Bleeding risk|risk of bleeding
Event|Event|Hospital Course|6912,6920|false|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|6912,6920|false|false|true|C0019080|Hemorrhage|bleeding
Drug|Biologically Active Substance|Hospital Course|6927,6930|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Hospital Course|6927,6930|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Hospital Course|6927,6930|false|false|false|||LDL
Procedure|Laboratory Procedure|Hospital Course|6927,6930|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Event|Event|Hospital Course|6935,6940|false|false|false|||found
Event|Event|Hospital Course|6955,6961|false|false|false|||wanted
Event|Event|Hospital Course|6965,6971|false|false|false|||change
Event|Event|Hospital Course|6976,6980|false|false|false|||from
Drug|Organic Chemical|Hospital Course|6982,6993|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|6982,6993|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Hospital Course|6982,6993|false|false|false|||simvastatin
Drug|Organic Chemical|Hospital Course|7013,7025|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7013,7025|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|7013,7025|false|false|false|||atorvastatin
Event|Event|Hospital Course|7037,7043|false|false|false|||issues
Drug|Pharmacologic Substance|Hospital Course|7050,7054|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Hospital Course|7050,7054|false|false|false|C0740721|Drug problem|drug
Finding|Finding|Hospital Course|7050,7059|false|false|false|C4036061|Drug-drug|drug-drug
Drug|Pharmacologic Substance|Hospital Course|7055,7059|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Hospital Course|7055,7059|false|false|false|C0740721|Drug problem|drug
Finding|Pathologic Function|Hospital Course|7055,7072|false|false|false|C0687133|Drug Interactions|drug interactions
Event|Event|Hospital Course|7060,7072|false|false|false|||interactions
Finding|Pathologic Function|Hospital Course|7060,7072|false|false|false|C0687133|Drug Interactions|interactions
Event|Event|Hospital Course|7083,7092|true|false|false|||insurance
Finding|Idea or Concept|Hospital Course|7083,7092|true|false|false|C0021672|Insurance|insurance
Event|Event|Hospital Course|7103,7108|true|false|false|||cover
Drug|Organic Chemical|Hospital Course|7110,7122|true|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7110,7122|true|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|7110,7122|true|false|false|||atorvastatin
Event|Event|Hospital Course|7142,7150|false|false|false|||switched
Drug|Organic Chemical|Hospital Course|7154,7165|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|Hospital Course|7154,7165|false|false|false|C0085542|pravastatin|pravastatin
Event|Event|Hospital Course|7154,7165|false|false|false|||pravastatin
Event|Event|Hospital Course|7176,7185|false|false|false|||discharge
Finding|Body Substance|Hospital Course|7176,7185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7176,7185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7176,7185|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7176,7185|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7194,7201|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|7194,7201|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Hospital Course|7225,7229|true|false|false|||feel
Drug|Organic Chemical|Hospital Course|7236,7242|true|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|7236,7242|true|false|false|C0633084|Plavix|Plavix
Event|Event|Hospital Course|7236,7242|true|false|false|||Plavix
Event|Event|Hospital Course|7247,7256|true|false|false|||necessary
Disorder|Disease or Syndrome|Hospital Course|7261,7264|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7261,7264|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7261,7264|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7261,7264|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7261,7264|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7261,7264|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7261,7264|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7261,7264|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|7274,7285|false|false|false|||neurologist
Event|Event|Hospital Course|7290,7299|false|false|false|||contacted
Event|Event|Hospital Course|7305,7311|false|false|false|||wanted
Drug|Organic Chemical|Hospital Course|7312,7318|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|7312,7318|false|false|false|C0633084|Plavix|Plavix
Event|Event|Hospital Course|7319,7328|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|7345,7355|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|7345,7355|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|7345,7355|false|false|false|||metoprolol
Event|Event|Hospital Course|7385,7394|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7385,7394|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|7404,7414|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|7404,7414|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|7404,7414|false|false|false|||metoprolol
Finding|Molecular Function|Hospital Course|7421,7425|false|false|false|C1150186|matrix metalloproteinase 7 activity|Pump
Event|Event|Hospital Course|7432,7436|false|false|false|||echo
Procedure|Health Care Activity|Hospital Course|7432,7436|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7432,7436|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|Hospital Course|7444,7450|false|false|false|||showed
Finding|Finding|Hospital Course|7451,7454|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Hospital Course|7451,7454|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Attribute|Clinical Attribute|Hospital Course|7462,7466|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|Hospital Course|7462,7466|false|false|false|||LVEF
Procedure|Diagnostic Procedure|Hospital Course|7462,7466|false|false|false|C3837267|LVEF (procedure)|LVEF
Phenomenon|Natural Phenomenon or Process|Hospital Course|7472,7479|false|false|false|C1705970|Electrical Current|current
Event|Event|Hospital Course|7481,7493|false|false|false|||presentation
Finding|Idea or Concept|Hospital Course|7481,7493|false|false|false|C0449450|Presentation|presentation
Event|Event|Hospital Course|7498,7508|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|7498,7508|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|7498,7513|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Space or Junction|Hospital Course|7514,7517|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|7514,7517|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|7518,7530|false|false|false|||exacerbation
Finding|Finding|Hospital Course|7518,7530|false|false|false|C4086268|Exacerbation|exacerbation
Anatomy|Tissue|Hospital Course|7547,7554|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Hospital Course|7547,7554|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Pathologic Function|Hospital Course|7547,7564|false|false|false|C0032227|Pleural effusion (disorder)|pleural effusions
Event|Event|Hospital Course|7555,7564|false|false|false|||effusions
Finding|Pathologic Function|Hospital Course|7555,7564|false|false|false|C0013687|effusion|effusions
Event|Event|Hospital Course|7566,7573|false|false|false|||dyspnea
Finding|Finding|Hospital Course|7566,7573|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|7566,7573|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7588,7598|false|false|false|C5441781|N-Terminal Fragment Brain Natriuretic Protein, human|NT-Pro-BNP
Drug|Biologically Active Substance|Hospital Course|7588,7598|false|false|false|C5441781|N-Terminal Fragment Brain Natriuretic Protein, human|NT-Pro-BNP
Event|Event|Hospital Course|7591,7598|false|false|false|||Pro-BNP
Event|Event|Hospital Course|7604,7607|false|false|false|||TTE
Procedure|Diagnostic Procedure|Hospital Course|7604,7607|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|Hospital Course|7609,7615|false|false|false|||showed
Finding|Intellectual Product|Hospital Course|7616,7620|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|Hospital Course|7621,7629|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|7621,7629|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|Hospital Course|7630,7636|false|false|false|||mitral
Finding|Finding|Hospital Course|7641,7649|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Hospital Course|7641,7649|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Event|Event|Hospital Course|7650,7659|false|false|false|||tricuspid
Event|Event|Hospital Course|7661,7674|false|false|false|||regurgitation
Finding|Finding|Hospital Course|7661,7674|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Hospital Course|7661,7674|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Hospital Course|7661,7674|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Attribute|Clinical Attribute|Hospital Course|7676,7680|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|Hospital Course|7676,7680|false|false|false|||LVEF
Procedure|Diagnostic Procedure|Hospital Course|7676,7680|false|false|false|C3837267|LVEF (procedure)|LVEF
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7693,7702|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|7693,7702|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|7693,7702|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|7693,7715|false|false|false|C0020542|Pulmonary Hypertension|pulmonary hypertension
Disorder|Disease or Syndrome|Hospital Course|7703,7715|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|7703,7715|false|false|false|||hypertension
Event|Event|Hospital Course|7721,7728|false|false|false|||changed
Drug|Organic Chemical|Hospital Course|7733,7737|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Hospital Course|7733,7737|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|Hospital Course|7733,7737|false|false|false|||HCTZ
Drug|Organic Chemical|Hospital Course|7741,7746|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|7741,7746|false|false|false|C0699992|Lasix|Lasix
Event|Event|Hospital Course|7741,7746|false|false|false|||Lasix
Event|Event|Hospital Course|7759,7768|false|false|false|||discharge
Finding|Body Substance|Hospital Course|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7759,7768|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7759,7768|false|false|false|C0030685|Patient Discharge|discharge
Drug|Pharmacologic Substance|Hospital Course|7775,7785|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|7775,7785|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|7775,7785|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|7794,7804|false|false|false|||uptitrated
Event|Event|Hospital Course|7808,7814|false|false|false|||needed
Disorder|Disease or Syndrome|Hospital Course|7819,7831|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|7819,7831|false|false|false|||Hypertension
Finding|Body Substance|Hospital Course|7837,7844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7837,7844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7837,7844|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7847,7859|false|false|false|||nephrologist
Event|Event|Hospital Course|7870,7876|false|false|false|||agreed
Drug|Pharmacologic Substance|Hospital Course|7896,7906|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Hospital Course|7896,7906|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|7907,7918|false|false|false|||adjustments
Finding|Functional Concept|Hospital Course|7907,7918|false|false|false|C0456081||adjustments
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7907,7918|false|false|false|C2945673|Clinical adjustment|adjustments
Event|Event|Hospital Course|7924,7935|false|false|false|||recommended
Finding|Idea or Concept|Hospital Course|7924,7935|false|false|false|C0034866|Recommendation|recommended
Event|Event|Hospital Course|7937,7944|false|false|false|||staying
Drug|Organic Chemical|Hospital Course|7955,7964|false|false|false|C0009014|clonidine|clonidine
Drug|Pharmacologic Substance|Hospital Course|7955,7964|false|false|false|C0009014|clonidine|clonidine
Event|Event|Hospital Course|7955,7964|false|false|false|||clonidine
Drug|Pharmacologic Substance|Hospital Course|7987,7997|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|7987,7997|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|7987,7997|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|7999,8012|false|false|false|||non-adherence
Finding|Functional Concept|Hospital Course|8014,8020|false|false|false|C0728831|Social|Social
Event|Event|Hospital Course|8021,8025|false|false|false|||work
Event|Occupational Activity|Hospital Course|8021,8025|false|false|false|C0043227|Work|work
Event|Event|Hospital Course|8030,8038|false|false|false|||involved
Event|Event|Hospital Course|8042,8051|false|false|false|||discharge
Finding|Body Substance|Hospital Course|8042,8051|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8042,8051|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8042,8051|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8042,8051|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Health Care Activity|Hospital Course|8042,8060|false|false|false|C0012622|Discharge Planning|discharge planning
Event|Event|Hospital Course|8052,8060|false|false|false|||planning
Finding|Functional Concept|Hospital Course|8052,8060|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|Hospital Course|8052,8060|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|Hospital Course|8079,8088|false|false|false|||assisting
Finding|Body Substance|Hospital Course|8093,8100|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8093,8100|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8093,8100|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|8101,8108|false|false|false|C4534363|At home|at home
Event|Event|Hospital Course|8104,8108|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8104,8108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8104,8108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8104,8108|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8113,8118|false|false|false|||added
Finding|Functional Concept|Hospital Course|8113,8118|false|false|false|C1524062|Additional|added
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8120,8130|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|8120,8130|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|8120,8130|false|false|false|||lisinopril
Drug|Organic Chemical|Hospital Course|8144,8149|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|8144,8149|false|false|false|C0699992|Lasix|Lasix
Event|Event|Hospital Course|8144,8149|false|false|false|||Lasix
Event|Event|Hospital Course|8166,8175|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|8177,8187|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|8177,8187|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|8177,8187|false|false|false|||nifedipine
Drug|Organic Chemical|Hospital Course|8206,8214|false|false|false|C0004147|atenolol|atenolol
Drug|Pharmacologic Substance|Hospital Course|8206,8214|false|false|false|C0004147|atenolol|atenolol
Event|Event|Hospital Course|8206,8214|false|false|false|||atenolol
Event|Event|Hospital Course|8219,8226|false|false|false|||stopped
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8239,8244|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|8239,8244|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|8239,8256|false|false|false|C1565489|Renal Insufficiency|renal dysfunction
Finding|Finding|Hospital Course|8239,8256|false|false|false|C3279454|Renal dysfunction|renal dysfunction
Disorder|Disease or Syndrome|Hospital Course|8245,8256|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|8245,8256|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|8245,8256|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|8245,8256|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|8245,8256|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Drug|Organic Chemical|Hospital Course|8266,8276|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8266,8276|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|8266,8276|false|false|false|||metoprolol
Event|Event|Hospital Course|8287,8294|false|false|false|||stopped
Event|Event|Hospital Course|8303,8314|false|false|false|||bradycardia
Finding|Finding|Hospital Course|8303,8314|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|Hospital Course|8327,8335|false|false|false|||continue
Finding|Intellectual Product|Hospital Course|8339,8343|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|8339,8349|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|8346,8349|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8346,8349|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|Hospital Course|8350,8360|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|8350,8360|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|8350,8360|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|8361,8367|false|false|false|||dosing
Event|Event|Hospital Course|8372,8376|false|false|false|||help
Event|Event|Hospital Course|8382,8392|false|false|false|||compliance
Finding|Finding|Hospital Course|8382,8392|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|Hospital Course|8382,8392|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|Hospital Course|8382,8392|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Disorder|Disease or Syndrome|Hospital Course|8399,8403|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|8399,8403|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|8399,8403|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|8399,8403|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Body Substance|Hospital Course|8409,8416|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8409,8416|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8409,8416|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8428,8437|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|8428,8437|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|8428,8437|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|8428,8437|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|8428,8437|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|8428,8437|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Disease or Syndrome|Hospital Course|8441,8445|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|8441,8445|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|8441,8445|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|8441,8445|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|8458,8466|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|8458,8466|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|8470,8479|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8470,8479|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|8484,8493|false|false|false|||responded
Drug|Organic Chemical|Hospital Course|8497,8506|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|8497,8506|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|8497,8506|false|false|false|||albuterol
Event|Event|Hospital Course|8516,8521|false|false|false|||given
Attribute|Clinical Attribute|Hospital Course|8525,8537|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Hospital Course|8525,8537|false|false|false|||prescription
Finding|Intellectual Product|Hospital Course|8525,8537|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Hospital Course|8525,8537|false|false|false|C0033080|Prescription (procedure)|prescription
Drug|Organic Chemical|Hospital Course|8542,8551|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|8542,8551|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|8542,8551|false|false|false|||albuterol
Finding|Gene or Genome|Hospital Course|8552,8555|false|false|false|C1422467|CIAO3 gene|prn
Finding|Idea or Concept|Hospital Course|8558,8570|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|Hospital Course|8593,8602|false|false|false|||scheduled
Attribute|Clinical Attribute|Hospital Course|8613,8619|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|8613,8619|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|8613,8619|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|8613,8619|false|false|false|C0038435|Stress|stress
Attribute|Clinical Attribute|Hospital Course|8620,8626|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|8620,8626|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|8620,8626|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|8620,8626|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|8620,8631|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Hospital Course|8627,8631|false|false|false|C4318744|Test - temporal region|test
Event|Event|Hospital Course|8627,8631|false|false|false|||test
Finding|Functional Concept|Hospital Course|8627,8631|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|8627,8631|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|8627,8631|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|8627,8631|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Hospital Course|8642,8648|false|false|false|||follow
Event|Activity|Hospital Course|8652,8664|false|false|false|C0003629|Appointments|appointments
Event|Event|Hospital Course|8652,8664|false|false|false|||appointments
Event|Event|Hospital Course|8704,8708|false|false|false|||work
Event|Event|Hospital Course|8712,8723|false|false|false|||uptitrating
Event|Event|Hospital Course|8728,8730|false|false|false|||BP
Disorder|Disease or Syndrome|Hospital Course|8732,8736|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Hospital Course|8732,8736|false|false|false|||meds
Finding|Intellectual Product|Hospital Course|8732,8736|false|false|false|C4284232|Medications|meds
Event|Event|Hospital Course|8740,8746|false|false|false|||needed
Event|Event|Hospital Course|8759,8763|false|false|false|||need
Event|Event|Hospital Course|8767,8771|false|false|false|||work
Finding|Body Substance|Hospital Course|8777,8784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8777,8784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8777,8784|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Pharmacologic Substance|Hospital Course|8788,8798|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|8788,8798|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|8788,8798|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Finding|Hospital Course|8788,8809|false|false|false|C2364172;C3489773|Adherence To Medication Regime;Medication Compliance|medication compliance
Finding|Individual Behavior|Hospital Course|8788,8809|false|false|false|C2364172;C3489773|Adherence To Medication Regime;Medication Compliance|medication compliance
Event|Event|Hospital Course|8799,8809|false|false|false|||compliance
Finding|Finding|Hospital Course|8799,8809|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Idea or Concept|Hospital Course|8799,8809|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Finding|Individual Behavior|Hospital Course|8799,8809|false|false|false|C1321605;C3244300;C4054143|Compliance behavior;Operational Compliance;Pulmonary compliance|compliance
Attribute|Clinical Attribute|Hospital Course|8813,8824|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8813,8824|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8813,8824|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8813,8824|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8813,8837|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8828,8837|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8828,8837|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|8839,8847|false|false|false|C0004147|atenolol|ATENOLOL
Drug|Pharmacologic Substance|Hospital Course|8839,8847|false|false|false|C0004147|atenolol|ATENOLOL
Drug|Biomedical or Dental Material|Hospital Course|8857,8863|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8870,8876|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|8880,8888|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8883,8888|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8883,8888|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|8889,8893|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|8889,8899|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|8896,8899|false|false|false|||day
Finding|Idea or Concept|Hospital Course|8896,8899|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8896,8899|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|8901,8910|false|false|false|C0009014|clonidine|CLONIDINE
Drug|Pharmacologic Substance|Hospital Course|8901,8910|false|false|false|C0009014|clonidine|CLONIDINE
Drug|Biomedical or Dental Material|Hospital Course|8920,8933|false|false|false|C5708820|24 Hour Release Patch Dosage Form|24 hour Patch
Drug|Biomedical or Dental Material|Hospital Course|8928,8933|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|8928,8933|false|false|false|||Patch
Finding|Finding|Hospital Course|8928,8933|false|false|false|C0332461|Plaque (lesion)|Patch
Event|Activity|Hospital Course|8943,8948|false|false|false|C1882509|put - instruction imperative|place
Event|Event|Hospital Course|8943,8948|false|false|false|||place
Finding|Functional Concept|Hospital Course|8943,8948|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|8943,8948|false|false|false|C1533810||place
Anatomy|Body Location or Region|Hospital Course|8952,8960|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|Hospital Course|8952,8960|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8952,8960|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Intellectual Product|Hospital Course|8961,8965|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Intellectual Product|Hospital Course|8969,8973|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|Hospital Course|8974,8985|false|false|false|C0070166|clopidogrel|CLOPIDOGREL
Drug|Pharmacologic Substance|Hospital Course|8974,8985|false|false|false|C0070166|clopidogrel|CLOPIDOGREL
Drug|Organic Chemical|Hospital Course|8987,8993|false|false|false|C0633084|Plavix|PLAVIX
Drug|Pharmacologic Substance|Hospital Course|8987,8993|false|false|false|C0633084|Plavix|PLAVIX
Drug|Biomedical or Dental Material|Hospital Course|9003,9009|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9014,9020|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|9024,9032|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9027,9032|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9027,9032|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9033,9037|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|Hospital Course|9041,9044|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9041,9044|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|Hospital Course|9045,9052|false|false|false|C0085155|Generic Drugs|generic
Event|Event|Hospital Course|9045,9052|false|false|false|||generic
Event|Event|Hospital Course|9056,9065|false|false|false|||available
Finding|Functional Concept|Hospital Course|9056,9065|false|false|false|C0470187|Availability of|available
Event|Event|Hospital Course|9085,9089|false|false|false|||call
Event|Activity|Hospital Course|9101,9112|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|9101,9112|false|false|false|||appointment
Drug|Organic Chemical|Hospital Course|9115,9126|false|false|false|C0033228|fenofibrate|FENOFIBRATE
Drug|Pharmacologic Substance|Hospital Course|9115,9126|false|false|false|C0033228|fenofibrate|FENOFIBRATE
Drug|Organic Chemical|Hospital Course|9115,9137|false|false|false|C0724585|fenofibrate micronized|FENOFIBRATE MICRONIZED
Drug|Pharmacologic Substance|Hospital Course|9115,9137|false|false|false|C0724585|fenofibrate micronized|FENOFIBRATE MICRONIZED
Event|Event|Hospital Course|9127,9137|false|false|false|||MICRONIZED
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9147,9154|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9147,9154|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9147,9154|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9159,9166|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9159,9166|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9159,9166|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|9170,9178|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9173,9178|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9173,9178|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9180,9184|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9180,9190|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9187,9190|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9187,9190|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9187,9190|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|9191,9210|false|false|false|C0020261|hydrochlorothiazide|HYDROCHLOROTHIAZIDE
Drug|Pharmacologic Substance|Hospital Course|9191,9210|false|false|false|C0020261|hydrochlorothiazide|HYDROCHLOROTHIAZIDE
Drug|Biomedical or Dental Material|Hospital Course|9219,9225|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9236,9242|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9236,9242|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|9246,9254|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9249,9254|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9249,9254|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9256,9260|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9256,9266|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9263,9266|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9263,9266|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9263,9266|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|9267,9277|false|false|false|C0028066|nifedipine|NIFEDIPINE
Drug|Pharmacologic Substance|Hospital Course|9267,9277|false|false|false|C0028066|nifedipine|NIFEDIPINE
Event|Event|Hospital Course|9267,9277|false|false|false|||NIFEDIPINE
Drug|Organic Chemical|Hospital Course|9279,9287|false|false|false|C1602464|Nifediac|NIFEDIAC
Drug|Pharmacologic Substance|Hospital Course|9279,9287|false|false|false|C1602464|Nifediac|NIFEDIAC
Drug|Organic Chemical|Hospital Course|9279,9290|false|false|false|C1330421|Nifediac CC|NIFEDIAC CC
Drug|Pharmacologic Substance|Hospital Course|9279,9290|false|false|false|C1330421|Nifediac CC|NIFEDIAC CC
Event|Event|Hospital Course|9288,9290|false|false|false|||CC
Drug|Biomedical or Dental Material|Hospital Course|9300,9306|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Hospital Course|9307,9315|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9307,9315|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|9316,9323|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9316,9323|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9316,9323|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9316,9323|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|9329,9335|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9329,9335|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|9339,9347|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9342,9347|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9342,9347|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9348,9352|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9348,9358|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9355,9358|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9355,9358|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9355,9358|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|9359,9372|false|false|false|C0017887|nitroglycerin|NITROGLYCERIN
Drug|Pharmacologic Substance|Hospital Course|9359,9372|false|false|false|C0017887|nitroglycerin|NITROGLYCERIN
Drug|Organic Chemical|Hospital Course|9374,9383|false|false|false|C0699241|Nitrostat|NITROSTAT
Drug|Pharmacologic Substance|Hospital Course|9374,9383|false|false|false|C0699241|Nitrostat|NITROSTAT
Drug|Biomedical or Dental Material|Hospital Course|9394,9400|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9394,9400|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|9394,9412|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Event|Event|Hospital Course|9402,9412|false|false|false|||Sublingual
Finding|Finding|Hospital Course|9402,9412|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|9402,9412|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Drug|Biomedical or Dental Material|Hospital Course|9418,9424|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9418,9424|false|false|false|||Tablet
Event|Event|Hospital Course|9447,9453|false|false|false|||needed
Finding|Gene or Genome|Hospital Course|9458,9461|false|false|false|C1422467|CIAO3 gene|prn
Anatomy|Body Location or Region|Hospital Course|9462,9467|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9462,9467|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9462,9472|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9462,9472|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9468,9472|false|true|false|C2598155||pain
Event|Event|Hospital Course|9468,9472|false|false|false|||pain
Finding|Functional Concept|Hospital Course|9468,9472|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9468,9472|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9477,9480|false|false|false|||use
Event|Event|Hospital Course|9484,9489|false|false|false|||doses
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9491,9500|false|false|false|C0886384|5 minutes Office visit|5 minutes
Drug|Organic Chemical|Hospital Course|9514,9520|true|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|Hospital Course|9514,9520|true|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|Hospital Course|9514,9520|true|false|false|||relief
Finding|Finding|Hospital Course|9514,9520|true|false|false|C0564405|Feeling relief|relief
Event|Event|Hospital Course|9525,9530|true|false|false|||visit
Finding|Social Behavior|Hospital Course|9525,9530|true|false|false|C0545082|Visit|visit
Drug|Organic Chemical|Hospital Course|9532,9542|true|false|false|C0034665|ranitidine|RANITIDINE
Drug|Pharmacologic Substance|Hospital Course|9532,9542|true|false|false|C0034665|ranitidine|RANITIDINE
Event|Event|Hospital Course|9532,9542|true|false|false|||RANITIDINE
Drug|Organic Chemical|Hospital Course|9532,9546|true|false|false|C0700466|ranitidine hydrochloride|RANITIDINE HCL
Drug|Pharmacologic Substance|Hospital Course|9532,9546|true|false|false|C0700466|ranitidine hydrochloride|RANITIDINE HCL
Disorder|Neoplastic Process|Hospital Course|9543,9546|true|false|false|C0023443|Hairy Cell Leukemia|HCL
Drug|Immunologic Factor|Hospital Course|9543,9546|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Drug|Inorganic Chemical|Hospital Course|9543,9546|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Drug|Pharmacologic Substance|Hospital Course|9543,9546|true|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCL
Event|Event|Hospital Course|9543,9546|true|false|false|||HCL
Drug|Biomedical or Dental Material|Hospital Course|9556,9562|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9567,9573|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|9577,9585|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9580,9585|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9580,9585|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9586,9590|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9586,9596|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9593,9596|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9593,9596|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9593,9596|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|9597,9608|false|false|false|C0074554|simvastatin|SIMVASTATIN
Drug|Pharmacologic Substance|Hospital Course|9597,9608|false|false|false|C0074554|simvastatin|SIMVASTATIN
Drug|Biomedical or Dental Material|Hospital Course|9617,9623|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9628,9634|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|9638,9646|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9641,9646|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9641,9646|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Attribute|Clinical Attribute|Hospital Course|9659,9670|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9659,9670|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9659,9670|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9659,9670|false|false|false|C4284232|Medications|Medications
Drug|Pharmacologic Substance|Hospital Course|9673,9676|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|9673,9676|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|9673,9676|false|false|false|C1418193|OTC gene|OTC
Drug|Organic Chemical|Hospital Course|9679,9686|false|false|false|C0004057|aspirin|ASPIRIN
Drug|Pharmacologic Substance|Hospital Course|9679,9686|false|false|false|C0004057|aspirin|ASPIRIN
Event|Event|Hospital Course|9679,9686|false|false|false|||ASPIRIN
Attribute|Clinical Attribute|Hospital Course|9688,9710|false|false|false|C4554471||ENTERIC COATED ASPIRIN
Drug|Organic Chemical|Hospital Course|9688,9710|false|false|false|C0718690|Aspirin Enteric Coated|ENTERIC COATED ASPIRIN
Drug|Pharmacologic Substance|Hospital Course|9688,9710|false|false|false|C0718690|Aspirin Enteric Coated|ENTERIC COATED ASPIRIN
Drug|Organic Chemical|Hospital Course|9703,9710|false|false|false|C0004057|aspirin|ASPIRIN
Drug|Pharmacologic Substance|Hospital Course|9703,9710|false|false|false|C0004057|aspirin|ASPIRIN
Event|Event|Hospital Course|9703,9710|false|false|false|||ASPIRIN
Drug|Biomedical or Dental Material|Hospital Course|9721,9727|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9721,9727|false|false|false|||Tablet
Attribute|Clinical Attribute|Hospital Course|9729,9736|false|false|false|C1545665|Views delayed|Delayed
Event|Event|Hospital Course|9738,9745|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9738,9745|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9738,9745|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9738,9745|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|9763,9769|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9763,9769|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|9773,9781|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9776,9781|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9776,9781|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9782,9786|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9782,9792|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9789,9792|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9789,9792|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9789,9792|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9793,9800|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Drug|Hormone|Hospital Course|9793,9800|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Drug|Pharmacologic Substance|Hospital Course|9793,9800|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|INSULIN
Event|Event|Hospital Course|9793,9800|false|false|false|||INSULIN
Finding|Gene or Genome|Hospital Course|9793,9800|false|false|false|C1337112|INS gene|INSULIN
Procedure|Laboratory Procedure|Hospital Course|9793,9800|false|false|false|C0202098|Insulin measurement|INSULIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9793,9804|false|false|false|C0021658|insulin isophane|INSULIN NPH
Drug|Hormone|Hospital Course|9793,9804|false|false|false|C0021658|insulin isophane|INSULIN NPH
Drug|Pharmacologic Substance|Hospital Course|9793,9804|false|false|false|C0021658|insulin isophane|INSULIN NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9801,9804|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|9801,9804|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|9801,9804|false|false|false|||NPH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9822,9829|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HUMULIN
Drug|Hormone|Hospital Course|9822,9829|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HUMULIN
Drug|Pharmacologic Substance|Hospital Course|9822,9829|false|false|false|C0020171;C0020172;C3538423|Humulin;Humulin S;Humulin insulin|HUMULIN
Event|Event|Hospital Course|9822,9829|false|false|false|||HUMULIN
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9822,9835|false|false|false|C0306367|HumuLIN 70/30|HUMULIN 70/30
Drug|Hormone|Hospital Course|9822,9835|false|false|false|C0306367|HumuLIN 70/30|HUMULIN 70/30
Drug|Pharmacologic Substance|Hospital Course|9822,9835|false|false|false|C0306367|HumuLIN 70/30|HUMULIN 70/30
Drug|Biomedical or Dental Material|Hospital Course|9860,9870|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|9860,9870|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|Hospital Course|9860,9870|false|false|false|||Suspension
Finding|Functional Concept|Hospital Course|9860,9870|false|false|false|C1705537|Suspension (action)|Suspension
Event|Event|Hospital Course|9876,9881|false|false|false|||units
Event|Event|Hospital Course|9885,9891|false|false|false|||dinner
Finding|Daily or Recreational Activity|Hospital Course|9885,9891|false|false|false|C4048877|Dinner|dinner
Event|Event|Hospital Course|9895,9901|false|false|false|||dinner
Finding|Daily or Recreational Activity|Hospital Course|9895,9901|false|false|false|C4048877|Dinner|dinner
Drug|Organic Chemical|Hospital Course|9902,9914|false|false|false|C0301532|Multivitamin preparation|MULTIVITAMIN
Drug|Pharmacologic Substance|Hospital Course|9902,9914|false|false|false|C0301532|Multivitamin preparation|MULTIVITAMIN
Drug|Vitamin|Hospital Course|9902,9914|false|false|false|C0301532|Multivitamin preparation|MULTIVITAMIN
Drug|Pharmacologic Substance|Hospital Course|9918,9921|false|false|false|C0013231|Drugs, Non-Prescription|OTC
Event|Event|Hospital Course|9918,9921|false|false|false|||OTC
Finding|Gene or Genome|Hospital Course|9918,9921|false|false|false|C1418193|OTC gene|OTC
Drug|Biomedical or Dental Material|Hospital Course|9925,9931|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|9936,9942|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|9946,9954|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9949,9954|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9949,9954|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|9955,9959|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9955,9965|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|9962,9965|false|false|false|||day
Finding|Idea or Concept|Hospital Course|9962,9965|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9962,9965|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|9968,9977|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9968,9977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9968,9977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9968,9977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9968,9977|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9968,9989|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9978,9989|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9978,9989|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9978,9989|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9978,9989|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9994,10005|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|9994,10005|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Biomedical or Dental Material|Hospital Course|10012,10018|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10032,10038|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10032,10038|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10067,10073|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|10078,10085|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10093,10106|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|10093,10106|false|false|false|C0017887|nitroglycerin|nitroglycerin
Drug|Biomedical or Dental Material|Hospital Course|10114,10120|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10114,10132|false|false|false|C0991582|Sublingual Tablet|Tablet, Sublingual
Finding|Finding|Hospital Course|10122,10132|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|10122,10132|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10133,10136|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10133,10136|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|10133,10136|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|10133,10136|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|10146,10152|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10146,10152|false|false|false|||Tablet
Finding|Finding|Hospital Course|10155,10165|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|10155,10165|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Finding|Hospital Course|10166,10176|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|10166,10176|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Event|Event|Hospital Course|10177,10180|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|10177,10180|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|10185,10191|false|false|false|||needed
Event|Event|Hospital Course|10196,10202|false|false|false|||needed
Anatomy|Body Location or Region|Hospital Course|10207,10212|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|10207,10212|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|10207,10217|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|10207,10217|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|10213,10217|false|false|false|C2598155||pain
Event|Event|Hospital Course|10213,10217|false|false|false|||pain
Finding|Functional Concept|Hospital Course|10213,10217|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10213,10217|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|10224,10228|false|false|false|||take
Drug|Biomedical or Dental Material|Hospital Course|10263,10269|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10263,10269|false|false|false|||Tablet
Finding|Finding|Hospital Course|10272,10282|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Functional Concept|Hospital Course|10272,10282|false|false|false|C0001565;C4521982|Sublingual (intended site);Sublingual Route of Administration|Sublingual
Finding|Idea or Concept|Hospital Course|10287,10294|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10302,10314|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|10302,10314|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|10302,10314|false|false|false|C0301532|Multivitamin preparation|multivitamin
Event|Event|Hospital Course|10302,10314|false|false|false|||multivitamin
Drug|Pharmacologic Substance|Hospital Course|10302,10325|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|10319,10325|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10319,10325|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10339,10345|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10339,10345|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10374,10380|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|10385,10392|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10400,10410|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|10400,10410|false|false|false|C0034665|ranitidine|ranitidine
Event|Event|Hospital Course|10400,10410|false|false|false|||ranitidine
Drug|Organic Chemical|Hospital Course|10400,10414|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Drug|Pharmacologic Substance|Hospital Course|10400,10414|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Disorder|Neoplastic Process|Hospital Course|10411,10414|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|10411,10414|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|10411,10414|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|10411,10414|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|10411,10414|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|10422,10428|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10442,10448|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10449,10451|false|false|false|||PO
Drug|Biomedical or Dental Material|Hospital Course|10477,10483|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|10488,10495|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10503,10514|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|Hospital Course|10503,10514|false|false|false|C0085542|pravastatin|pravastatin
Event|Event|Hospital Course|10503,10514|false|false|false|||pravastatin
Drug|Biomedical or Dental Material|Hospital Course|10521,10527|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10528,10531|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|10541,10547|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10541,10547|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10576,10582|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10587,10594|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10587,10594|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10602,10609|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|10602,10609|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|10602,10609|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Hospital Course|10616,10622|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10616,10632|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10633,10636|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10633,10636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|10633,10636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|10633,10636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|10646,10652|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10646,10652|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10646,10662|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Event|Event|Hospital Course|10654,10662|false|false|false|||Chewable
Drug|Biomedical or Dental Material|Hospital Course|10691,10697|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10691,10697|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10691,10707|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Event|Event|Hospital Course|10712,10719|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10712,10719|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10727,10737|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|10727,10737|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|Hospital Course|10727,10737|false|false|false|||lisinopril
Drug|Biomedical or Dental Material|Hospital Course|10744,10750|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10764,10770|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10764,10770|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|10799,10805|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10810,10817|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10810,10817|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10825,10835|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10825,10835|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|Hospital Course|10825,10835|false|false|false|||nifedipine
Drug|Biomedical or Dental Material|Hospital Course|10842,10848|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Hospital Course|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10858,10865|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10858,10865|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10858,10865|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10858,10865|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|10879,10885|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10879,10885|false|false|false|||Tablet
Finding|Finding|Hospital Course|10887,10895|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10887,10895|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10896,10903|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10896,10903|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10896,10903|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10896,10903|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|10931,10937|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|10938,10946|false|false|false|||Extended
Finding|Finding|Hospital Course|10938,10946|false|true|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10938,10946|false|true|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10948,10955|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10948,10955|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10948,10955|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10948,10955|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|10960,10967|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|10960,10967|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|10975,10985|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|10975,10985|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|10975,10985|false|false|false|||furosemide
Drug|Biomedical or Dental Material|Hospital Course|10992,10998|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11012,11018|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11012,11018|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|11047,11053|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|11058,11065|false|false|false|C0807726|refill|Refills
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11074,11081|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|11074,11081|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|11074,11081|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|Hospital Course|11074,11081|false|false|false|||insulin
Finding|Gene or Genome|Hospital Course|11074,11081|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|11074,11081|false|false|false|C0202098|Insulin measurement|insulin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11074,11085|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Hormone|Hospital Course|11074,11085|false|false|false|C0021658|insulin isophane|insulin NPH
Drug|Pharmacologic Substance|Hospital Course|11074,11085|false|false|false|C0021658|insulin isophane|insulin NPH
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11082,11085|false|false|false|C0027442|Nasopharynx|NPH
Disorder|Disease or Syndrome|Hospital Course|11082,11085|false|false|false|C0020258|Hydrocephalus, Normal Pressure|NPH
Event|Event|Hospital Course|11082,11085|false|false|false|||NPH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11122,11129|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Hormone|Hospital Course|11122,11129|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Drug|Pharmacologic Substance|Hospital Course|11122,11129|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|Insulin
Event|Event|Hospital Course|11122,11129|false|false|false|||Insulin
Finding|Gene or Genome|Hospital Course|11122,11129|false|false|false|C1337112|INS gene|Insulin
Procedure|Laboratory Procedure|Hospital Course|11122,11129|false|false|false|C0202098|Insulin measurement|Insulin
Drug|Organic Chemical|Hospital Course|11130,11133|false|false|false|C0070220|penclomedine|Pen
Drug|Pharmacologic Substance|Hospital Course|11130,11133|false|false|false|C0070220|penclomedine|Pen
Finding|Gene or Genome|Hospital Course|11130,11133|false|false|false|C1424886;C1428887;C1823520|PCSK1N gene;PUM3 gene;TSPAN33 gene|Pen
Event|Event|Hospital Course|11135,11138|false|false|false|||Sig
Event|Event|Hospital Course|11158,11170|false|false|false|||Subcutaneous
Finding|Functional Concept|Hospital Course|11158,11170|false|false|false|C1522438|Subcutaneous Route of Administration|Subcutaneous
Event|Event|Hospital Course|11200,11207|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|11200,11207|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11216,11225|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|11216,11225|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|11216,11225|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|11216,11233|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|11216,11233|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|11226,11233|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|11226,11233|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|11226,11233|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|11226,11233|false|false|false|||sulfate
Disorder|Disease or Syndrome|Hospital Course|11251,11254|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|11251,11254|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|11251,11254|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|11255,11262|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|Hospital Course|11263,11270|false|false|false|||Inhaler
Finding|Functional Concept|Hospital Course|11263,11270|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Hospital Course|11287,11297|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|11287,11297|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Hospital Course|11317,11323|false|false|false|||needed
Event|Event|Hospital Course|11328,11337|false|false|false|||shortness
Event|Event|Hospital Course|11342,11348|false|false|false|||breath
Finding|Body Substance|Hospital Course|11342,11348|false|false|false|C0225386|Breath|breath
Event|Event|Hospital Course|11352,11360|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|11352,11360|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|11370,11377|false|false|false|||inhaler
Finding|Functional Concept|Hospital Course|11370,11377|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Finding|Idea or Concept|Hospital Course|11379,11386|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|11393,11402|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11393,11402|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11393,11402|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11393,11402|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11393,11402|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|11393,11414|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|11393,11414|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|11403,11414|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|11403,11414|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|11403,11414|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|11416,11420|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|11416,11420|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|11416,11420|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|11416,11420|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|11426,11433|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|11426,11433|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|11436,11444|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|11436,11444|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|11452,11461|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11452,11461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11452,11461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11452,11461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11452,11461|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11452,11471|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|11462,11471|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|11462,11471|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|11462,11471|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|11462,11471|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|11462,11471|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|11474,11486|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|11474,11486|false|false|false|||Hypertension
Finding|Finding|Hospital Course|11492,11504|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Disorder|Disease or Syndrome|Hospital Course|11492,11512|false|false|false|C0745138|Hypertensive Urgency|hypertensive urgency
Event|Event|Hospital Course|11505,11512|false|false|false|||urgency
Anatomy|Tissue|Hospital Course|11514,11524|false|false|false|C0027061|Myocardium|Myocardial
Attribute|Clinical Attribute|Hospital Course|11514,11535|false|false|false|C2926063||Myocardial infarction
Disorder|Disease or Syndrome|Hospital Course|11514,11535|false|false|false|C0027051|Myocardial Infarction|Myocardial infarction
Event|Event|Hospital Course|11525,11535|false|false|false|||infarction
Finding|Pathologic Function|Hospital Course|11525,11535|false|false|false|C0021308|Infarction|infarction
Event|Event|Hospital Course|11536,11546|false|false|false|||attributed
Finding|Idea or Concept|Hospital Course|11550,11556|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11550,11556|false|false|false|C0441516|Demand (clinical)|demand
Event|Event|Hospital Course|11557,11568|false|false|false|||myonecrosis
Finding|Pathologic Function|Hospital Course|11557,11568|false|false|false|C0235957|Muscle necrosis|myonecrosis
Finding|Intellectual Product|Hospital Course|11570,11575|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Finding|Intellectual Product|Hospital Course|11579,11586|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|11579,11586|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|Hospital Course|11587,11591|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11592,11603|false|false|false|C0018827|Heart Ventricle|ventricular
Attribute|Clinical Attribute|Hospital Course|11604,11613|false|false|false|C0012000|Diastole|diastolic
Disorder|Disease or Syndrome|Hospital Course|11604,11627|false|false|false|C1135196|Heart Failure, Diastolic|diastolic heart failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11614,11619|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Hospital Course|11614,11619|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Hospital Course|11614,11619|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Hospital Course|11614,11627|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Hospital Course|11620,11627|false|false|false|||failure
Finding|Functional Concept|Hospital Course|11620,11627|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|11620,11627|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|11620,11627|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Hospital Course|11629,11636|false|false|false|||Chronic
Finding|Intellectual Product|Hospital Course|11629,11636|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|11629,11636|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|11629,11651|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Finding|Classification|Hospital Course|11629,11658|false|false|false|C2074731|chronic kidney disease stage|Chronic kidney disease, stage
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11637,11643|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|11637,11643|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|11637,11643|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|11637,11643|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11637,11643|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|11637,11651|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|11644,11651|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|11644,11651|false|false|false|||disease
Attribute|Clinical Attribute|Hospital Course|11653,11658|false|false|false|C1300072|Tumor stage|stage
Event|Event|Hospital Course|11653,11658|false|false|false|||stage
Event|Event|Hospital Course|11664,11671|false|false|false|||Chronic
Finding|Intellectual Product|Hospital Course|11664,11671|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|11664,11671|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|11664,11701|false|false|false|C0024117|Chronic Obstructive Airway Disease|Chronic obstructive pulmonary disease
Finding|Functional Concept|Hospital Course|11672,11683|false|false|false|C0549186|Obstructed|obstructive
Disorder|Disease or Syndrome|Hospital Course|11672,11701|false|false|false|C0600260|Lung Diseases, Obstructive|obstructive pulmonary disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11684,11693|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|11684,11693|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|11684,11693|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|Hospital Course|11684,11701|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|Hospital Course|11684,11701|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|Hospital Course|11694,11701|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|11694,11701|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11709,11719|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11720,11729|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Hospital Course|11730,11736|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|11730,11736|false|false|false|||stroke
Finding|Finding|Hospital Course|11730,11736|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Hospital Course|11738,11752|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Hospital Course|11738,11752|false|false|false|||Hyperlipidemia
Finding|Finding|Hospital Course|11738,11752|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Disorder|Disease or Syndrome|Hospital Course|11754,11762|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Hospital Course|11754,11771|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Event|Event|Hospital Course|11763,11771|false|false|false|||mellitus
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11782,11789|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|11782,11789|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|11782,11789|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|11782,11789|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|11782,11789|false|false|false|C0202098|Insulin measurement|insulin
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11782,11797|false|false|false|C5442411|Insulin therapy|insulin therapy
Event|Event|Hospital Course|11790,11797|false|false|false|||therapy
Finding|Finding|Hospital Course|11790,11797|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|11790,11797|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11790,11797|false|false|false|C0087111|Therapeutic procedure|therapy
Drug|Pharmacologic Substance|Hospital Course|11799,11809|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11799,11809|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Finding|Hospital Course|11799,11823|false|false|false|C0746935|Medication Nonadherence|Medication non-adherence
Event|Event|Hospital Course|11810,11823|false|false|false|||non-adherence
Finding|Mental Process|Discharge Condition|11847,11853|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|11847,11860|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|11847,11860|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|11854,11860|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|11854,11860|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11862,11867|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|11862,11867|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|11872,11880|false|false|false|||coherent
Finding|Finding|Discharge Condition|11872,11880|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|11882,11887|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|11882,11904|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|11882,11904|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|11891,11904|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|11891,11904|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|11891,11904|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|11906,11911|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|11906,11911|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|11906,11911|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|11906,11911|false|false|false|||Alert
Finding|Finding|Discharge Condition|11906,11911|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|11906,11911|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|11906,11911|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|11916,11927|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|11916,11927|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|11929,11937|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|11929,11937|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|11929,11937|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11938,11944|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11938,11944|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11938,11944|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|11946,11956|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|11946,11956|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11946,11956|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11946,11956|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11946,11956|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11959,11970|false|false|false|||Independent
Finding|Finding|Discharge Condition|11959,11970|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|11959,11970|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|11998,12002|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|12023,12031|false|false|false|||admitted
Event|Event|Discharge Instructions|12036,12045|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|12036,12055|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|12036,12055|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|12049,12055|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|12066,12071|false|false|false|||found
Disorder|Disease or Syndrome|Discharge Instructions|12090,12095|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|12090,12095|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|12090,12095|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|12090,12104|true|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|12090,12104|true|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|12090,12104|true|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Discharge Instructions|12096,12104|true|false|false|||pressure
Finding|Finding|Discharge Instructions|12096,12104|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|12096,12104|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|12096,12104|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|12096,12104|true|false|false|C0033095||pressure
Event|Event|Discharge Instructions|12108,12117|true|false|false|||admission
Procedure|Health Care Activity|Discharge Instructions|12108,12117|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Mental Process|Discharge Instructions|12125,12132|true|false|false|C0542559|contextual factors|setting
Attribute|Clinical Attribute|Discharge Instructions|12160,12171|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12160,12171|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12160,12171|true|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12160,12171|true|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12186,12194|false|false|false|||obtained
Event|Event|Discharge Instructions|12199,12213|false|false|false|||echocargiogram
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12222,12227|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|12222,12227|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|12222,12227|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Discharge Instructions|12234,12240|false|false|false|||showed
Disorder|Injury or Poisoning|Discharge Instructions|12246,12252|false|false|false|C0080194|Muscle strain|strain
Event|Event|Discharge Instructions|12246,12252|false|false|false|||strain
Finding|Idea or Concept|Discharge Instructions|12246,12252|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|Discharge Instructions|12246,12252|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|Discharge Instructions|12246,12252|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|Discharge Instructions|12246,12252|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12262,12267|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|12262,12267|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|Discharge Instructions|12262,12267|false|false|false|||heart
Finding|Sign or Symptom|Discharge Instructions|12262,12267|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Finding|Discharge Instructions|12268,12276|false|false|false|C0332149|Possible|possibly
Drug|Organic Chemical|Discharge Instructions|12277,12284|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Discharge Instructions|12277,12284|false|false|false|||related
Finding|Finding|Discharge Instructions|12277,12284|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Discharge Instructions|12277,12284|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|Discharge Instructions|12302,12307|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|12302,12307|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|12302,12307|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|12302,12317|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|Discharge Instructions|12308,12317|false|false|false|||pressures
Finding|Finding|Discharge Instructions|12308,12317|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|Discharge Instructions|12308,12317|false|false|false|C0033095||pressures
Event|Event|Discharge Instructions|12332,12341|false|false|false|||contacted
Finding|Classification|Discharge Instructions|12351,12361|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|12351,12361|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Attribute|Clinical Attribute|Discharge Instructions|12362,12368|false|false|true|C1718621|W stress|stress
Drug|Organic Chemical|Discharge Instructions|12362,12368|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Discharge Instructions|12362,12368|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Event|Event|Discharge Instructions|12362,12368|false|false|false|||stress
Finding|Finding|Discharge Instructions|12362,12368|false|false|true|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Discharge Instructions|12362,12373|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Discharge Instructions|12369,12373|false|false|false|C4318744|Test - temporal region|test
Event|Event|Discharge Instructions|12369,12373|false|false|false|||test
Finding|Functional Concept|Discharge Instructions|12369,12373|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|12369,12373|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|12369,12373|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|12369,12373|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Discharge Instructions|12389,12398|false|false|false|||completed
Finding|Idea or Concept|Discharge Instructions|12410,12414|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Idea or Concept|Discharge Instructions|12415,12420|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|Discharge Instructions|12415,12420|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|Discharge Instructions|12435,12445|false|false|false|||prescribed
Finding|Finding|Discharge Instructions|12454,12457|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|12454,12457|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|12454,12469|false|false|false|C1718097|New medications|new medications
Attribute|Clinical Attribute|Discharge Instructions|12458,12469|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12458,12469|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12458,12469|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12458,12469|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12473,12478|false|false|false|||shown
Event|Event|Discharge Instructions|12508,12512|false|false|false|||come
Event|Event|Discharge Instructions|12521,12525|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|12521,12525|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|12521,12525|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|12521,12525|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|12529,12533|false|false|false|||help
Event|Event|Discharge Instructions|12539,12547|false|false|false|||managing
Attribute|Clinical Attribute|Discharge Instructions|12554,12565|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12554,12565|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12554,12565|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12554,12565|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12578,12585|false|false|false|||dispose
Finding|Idea or Concept|Discharge Instructions|12598,12602|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|12598,12602|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|12598,12602|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|12603,12614|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12603,12614|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12603,12614|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12603,12614|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12625,12629|false|false|false|||take
Attribute|Clinical Attribute|Discharge Instructions|12634,12645|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|12634,12645|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|12634,12645|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|12634,12645|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|12646,12651|false|false|false|||shown
Event|Event|Discharge Instructions|12660,12669|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|12660,12669|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|12660,12669|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|12660,12669|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|12660,12669|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Discharge Instructions|12670,12679|false|false|false|||paperwork
Drug|Inorganic Chemical|Medications|12695,12699|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Medications|12695,12699|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Medications|12695,12699|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|Medications|12695,12699|false|false|false|||STOP
Finding|Gene or Genome|Medications|12695,12699|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|Medications|12700,12719|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Medications|12700,12719|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Inorganic Chemical|Medications|12720,12724|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Medications|12720,12724|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Medications|12720,12724|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|Medications|12720,12724|false|false|false|||STOP
Finding|Gene or Genome|Medications|12720,12724|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|Medications|12725,12736|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Medications|12725,12736|false|false|false|C0074554|simvastatin|Simvastatin
Event|Event|Medications|12725,12736|false|false|false|||Simvastatin
Drug|Inorganic Chemical|Medications|12737,12741|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Medications|12737,12741|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Medications|12737,12741|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|Medications|12737,12741|false|false|false|||STOP
Finding|Gene or Genome|Medications|12737,12741|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|Medications|12742,12751|false|false|false|C0009014|clonidine|Clonidine
Drug|Pharmacologic Substance|Medications|12742,12751|false|false|false|C0009014|clonidine|Clonidine
Event|Event|Medications|12742,12751|false|false|false|||Clonidine
Drug|Inorganic Chemical|Medications|12752,12756|false|false|false|C0723457|Stop brand of fluoride|STOP
Drug|Pharmacologic Substance|Medications|12752,12756|false|false|false|C0723457|Stop brand of fluoride|STOP
Event|Activity|Medications|12752,12756|false|false|false|C1947925|Stop (Instruction Imperative)|STOP
Event|Event|Medications|12752,12756|false|false|false|||STOP
Finding|Gene or Genome|Medications|12752,12756|false|false|false|C1417022|MAP6 gene|STOP
Drug|Organic Chemical|Medications|12757,12765|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|Medications|12757,12765|false|false|false|C0004147|atenolol|Atenolol
Finding|Finding|Medications|12773,12776|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Medications|12773,12776|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|Medications|12773,12787|false|false|false|C0428977|Bradycardia|low heart rate
Anatomy|Body Part, Organ, or Organ Component|Medications|12777,12782|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Medications|12777,12782|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Medications|12777,12782|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Medications|12777,12787|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Medications|12777,12787|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Medications|12777,12787|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Medications|12783,12787|false|false|false|C0871208|Rating (action)|rate
Event|Event|Medications|12783,12787|false|false|false|||rate
Finding|Idea or Concept|Medications|12783,12787|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Medications|12788,12794|false|false|false|||CHANGE
Finding|Functional Concept|Medications|12788,12794|false|false|false|C0392747|Changing|CHANGE
Procedure|Therapeutic or Preventive Procedure|Medications|12788,12794|false|false|false|C4319952|Change - procedure|CHANGE
Finding|Intellectual Product|Medications|12809,12813|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Food|Medications|12820,12825|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|Medications|12820,12825|false|false|false|||START
Finding|Intellectual Product|Medications|12820,12825|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Medications|12820,12825|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Amino Acid, Peptide, or Protein|Medications|12826,12836|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Medications|12826,12836|false|false|false|C0065374|lisinopril|Lisinopril
Finding|Intellectual Product|Medications|12842,12846|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Food|Medications|12853,12858|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|Medications|12853,12858|false|false|false|||START
Finding|Intellectual Product|Medications|12853,12858|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Medications|12853,12858|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Drug|Organic Chemical|Medications|12859,12864|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Medications|12859,12864|false|false|false|C0699992|Lasix|Lasix
Finding|Intellectual Product|Medications|12870,12874|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Food|Medications|12881,12886|false|false|false|C0452588|Start brand of breakfast cereal|START
Event|Event|Medications|12881,12886|false|false|false|||START
Finding|Intellectual Product|Medications|12881,12886|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Medications|12881,12886|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Finding|Intellectual Product|Medications|12902,12906|false|false|false|C1720092|Once - dosing instruction fragment|once
Event|Event|Medications|12921,12931|true|false|false|||experience
Anatomy|Body Location or Region|Medications|12936,12941|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Medications|12936,12941|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Medications|12936,12946|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Medications|12936,12946|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Medications|12942,12946|true|false|false|C2598155||pain
Event|Event|Medications|12942,12946|true|false|false|||pain
Finding|Functional Concept|Medications|12942,12946|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|12942,12946|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|12958,12967|true|false|false|||shortness
Attribute|Clinical Attribute|Medications|12958,12977|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Medications|12958,12977|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Medications|12971,12977|true|false|false|C0225386|Breath|breath
Event|Event|Medications|12993,13001|true|false|false|||symptoms
Finding|Functional Concept|Medications|12993,13001|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Medications|12993,13001|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Medications|13028,13032|false|false|false|||call
Event|Event|Medications|13036,13040|false|false|false|||come
Event|Event|Medications|13051,13060|false|false|false|||emergency
Finding|Finding|Medications|13051,13060|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Medications|13051,13060|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Medications|13051,13060|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Medications|13051,13060|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Medications|13051,13060|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Medications|13051,13060|false|false|false|C1553500|emergency encounter|emergency
Finding|Idea or Concept|Medications|13061,13071|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Event|Event|Medications|13084,13094|false|false|false|||evaluation
Finding|Idea or Concept|Medications|13084,13094|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Medications|13084,13094|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|Medications|13111,13119|false|false|false|||allowing
Event|Event|Medications|13137,13148|false|false|false|||participate
Event|Activity|Medications|13157,13161|false|false|false|C1947933|care activity|care
Event|Event|Medications|13157,13161|false|false|false|||care
Finding|Finding|Medications|13157,13161|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Medications|13157,13161|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Health Care Activity|Medications|13165,13173|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|13174,13186|false|false|false|C3263700||Instructions
Event|Event|Medications|13174,13186|false|false|false|||Instructions
Finding|Intellectual Product|Medications|13174,13186|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

