CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Neurosurgical Procedures|Procedure|false|false||NEUROSURGERYnull|Science of neurosurgery|Title|false|false||NEUROSURGERYnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|false|false||Drugsnull|Drugs - dental services|Procedure|false|false||Drugsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Gait, Unsteady|Finding|false|false||Gait instabilitynull|Gait|Finding|false|false||Gaitnull|Instability|Finding|false|false||instabilitynull|multiple falls|Finding|false|false||multiple fallsnull|Numerous|LabModifier|false|false||multiplenull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Pleasant|Finding|false|false|C0230370|pleasantnull|Structure of right hand|Anatomy|false|false|C2987187;C1706180;C1561543;C1561544|right handednull|Right handed|Subject|false|false||right handednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Transaction counts and value totals - year|Finding|false|false|C0230370|year
null|Precision - year|Finding|false|false|C0230370|yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Male Gender|Finding|false|false|C0230370|malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Atrial Fibrillation|Disorder|false|false||Afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||Afibnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Coordination of Benefits - Independent|Finding|false|false||independent
null|Religious Affiliation - Independent|Finding|false|false||independent
null|Independence|Finding|false|false||independent
null|Independently able|Finding|false|false||independentnull|wife|Subject|false|false||wifenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|personal health|Finding|false|false||state of healthnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Health|Finding|false|false||healthnull|Middle|Modifier|false|false||midnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|wife|Subject|false|false||wifenull|Menstruation|Finding|false|false||periodsnull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|Gait, Unsteady|Finding|false|false||gait instabilitynull|Gait|Finding|false|false||gaitnull|Instability|Finding|false|false||instabilitynull|History of fall|Finding|false|false||a fallnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|month|Time|false|false||monthsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Several|LabModifier|false|false||severalnull|Bone structure of rib|Anatomy|false|false||ribsnull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Data Table|Finding|false|false||tablenull|Table - furniture|Device|false|false||tablenull|Craniocerebral Trauma|Disorder|true|false|C0018670;C0152336|head traumanull|Problems with head|Disorder|true|false|C0018670;C0152336|headnull|Procedure on head|Procedure|true|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0548346;C0362076;C0018674;C0876917;C3714660;C3263723;C1368081|head
null|Head|Anatomy|false|false|C0548346;C0362076;C0018674;C0876917;C3714660;C3263723;C1368081|headnull|Head Device|Device|true|false||headnull|Physical trauma|Disorder|true|false|C0018670;C0152336|trauma
null|Traumatic injury|Disorder|true|false|C0018670;C0152336|trauma
null|Trauma|Disorder|true|false|C0018670;C0152336|traumanull|Trauma assessment and care|Procedure|true|false|C0018670;C0152336|traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Speech|Finding|false|false||speechnull|Speech assessment|Procedure|false|false||speechnull|General unsteadiness|Finding|false|false||unsteadinessnull|Past 6 Months|Time|false|false||past 6 monthsnull|6 months|Time|false|false||6 monthsnull|month|Time|false|false||monthsnull|wife|Subject|false|false||wifenull|Much|Finding|false|false||muchnull|Diuretics|Drug|false|false||diureticsnull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Last|Modifier|false|false||Lastnull|Night time|Time|false|false||nightnull|Paper|Device|false|false||papersnull|Dining room|Device|false|false||dining roomnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Data Table|Finding|false|false||tablenull|Table - furniture|Device|false|false||tablenull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Location|Modifier|false|false||LOCnull|Craniocerebral Trauma|Disorder|true|false|C0018670;C0152336|head traumanull|Problems with head|Disorder|true|false|C0018670;C0152336|headnull|Procedure on head|Procedure|true|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0548346;C3714660;C3263723;C1368081;C0362076;C0018674;C0876917|head
null|Head|Anatomy|false|false|C0548346;C3714660;C3263723;C1368081;C0362076;C0018674;C0876917|headnull|Head Device|Device|true|false||headnull|Physical trauma|Disorder|false|false|C0018670;C0152336|trauma
null|Traumatic injury|Disorder|false|false|C0018670;C0152336|trauma
null|Trauma|Disorder|false|false|C0018670;C0152336|traumanull|Trauma assessment and care|Procedure|false|false|C0018670;C0152336|traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Continuous|Finding|false|false||continuenull|Work|Event|false|false||worknull|wife|Subject|false|false||wifenull|Bathroom|Device|false|false||bathroom
null|Toilet Facilities|Device|false|false||bathroomnull|Location|Modifier|false|false||LOCnull|Problems with head|Disorder|true|false|C0018670;C0152336|headnull|Procedure on head|Procedure|true|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076|head
null|Head|Anatomy|false|false|C0876917;C0362076|headnull|Head Device|Device|true|false||headnull|Physical trauma|Disorder|false|false||trauma
null|Traumatic injury|Disorder|false|false||trauma
null|Trauma|Disorder|false|false||traumanull|Trauma assessment and care|Procedure|false|false||traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|Instability|Finding|false|false||instabilitynull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Tongue biting|Disorder|false|false|C0040408|tongue bitingnull|Benign neoplasm of tongue|Disorder|false|false|C0040408|tonguenull|Procedure on tongue|Procedure|false|false|C0040408|tonguenull|Tongue|Anatomy|false|false|C0005658;C0872394;C0496930;C0154017;C0154091;C0872388;C0153933;C2584293;C0241424;C0876938;C4319531|tonguenull|bite injury|Disorder|false|false|C0040408|bitingnull|Biting|Finding|false|false|C0040408|bitingnull|Loss (adaptation)|Finding|false|false|C0021853|lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Intestines|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091;C5890125;C0876938;C4319531|bowelnull|Bladder Continence Question|Finding|false|false|C0021853;C0005682;C0040408|bladder continence
null|Urinary bladder control|Finding|false|false|C0021853;C0005682;C0040408|bladder continencenull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0040408;C0005682;C0021853|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0040408;C0005682;C0021853|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0040408;C0005682;C0021853|bladdernull|Procedures on bladder|Procedure|false|false|C0005682;C0040408;C0021853|bladdernull|Urinary Bladder|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091;C0876938;C4319531|bladdernull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|Morning|Time|false|false||morningnull|Presentation|Finding|false|false||presentationnull|wife|Subject|false|false||wifenull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|elongation factor DmS-II|Drug|false|false||DM IInull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Oral hypoglycemic|Drug|false|false|C0226896|oral hypoglycemicsnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C5203106;C4522223;C1550472;C1272919;C1527415;C4521986;C0359086|oralnull|Oral|Modifier|false|false||oralnull|Hypoglycemic Agents|Drug|false|false||hypoglycemicsnull|IPSS-R Risk Category Low|Finding|false|false|C0226896|low
null|IPSS Risk Category Low|Finding|false|false|C0226896|low
null|low confidentiality|Finding|false|false|C0226896|lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Neurologists|Subject|false|false||neurologistnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|null|Time|false|false||priornull|CAT scan of head|Procedure|false|false|C0018670;C0152336|CT headnull|null|Attribute|false|false|C0018670;C0152336|CT headnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C1561540;C0876917;C0202691;C0362076;C0881943|head
null|Head|Anatomy|false|false|C1561540;C0876917;C0202691;C0362076;C0881943|headnull|Head Device|Device|false|false||headnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Transaction counts and value totals - week|Finding|false|false|C0018670;C0152336|weeknull|week|Time|false|false||weeknull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917;C0019080|head
null|Head|Anatomy|false|false|C0362076;C0876917;C0019080|headnull|Head Device|Device|false|false||headnull|Hemorrhage|Finding|false|false|C0018670;C0152336|bleednull|malignant neoplasm of frontal lobe|Disorder|false|false|C0796494;C0016733|frontal lobenull|frontal lobe|Anatomy|false|false|C3539671;C1428707;C0153635;C4283905;C1546709;C2700045;C0577573;C0577559;C1414542|frontal lobenull|Coronal (qualifier value)|Modifier|false|false||frontalnull|AKT1S1 wt Allele|Finding|false|false|C0016733;C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0016733;C0796494|lobenull|lobe|Anatomy|false|false|C4283905;C1546709;C2700045;C0577573;C0577559;C1414542;C0153635;C3539671;C1428707|lobenull|Mass of body structure|Finding|false|false|C0796494;C0016733|mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false|C0796494;C0016733|mass
null|null|Finding|false|false|C0796494;C0016733|mass
null|FBN1 wt Allele|Finding|false|false|C0796494;C0016733|mass
null|FBN1 gene|Finding|false|false|C0796494;C0016733|mass
null|Mass of body region|Finding|false|false|C0796494;C0016733|massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Midline Shift|Finding|true|false|C1660780|midline shiftnull|midline cell component|Anatomy|false|false|C2347509;C0333051;C4086580|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|shift displacement|Finding|true|false|C1660780|shiftnull|Physical Shift|Phenomenon|true|false|C1660780|shiftnull|Neurosurgical Procedures|Procedure|false|false||Neurosurgerynull|Science of neurosurgery|Title|false|false||Neurosurgerynull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||mass
null|Mass of body structure|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Terminology Role Entity|Finding|false|false||role
null|Role|Finding|false|false||role
null|Security Role Object|Finding|false|false||role
null|Social Role|Finding|false|false||role
null|role - RoleClass|Finding|false|false||role
null|NCI Thesaurus Role|Finding|false|false||rolenull|null|Attribute|false|false||rolenull|Generic Role|Modifier|false|false||rolenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recent|Time|false|false||recentnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|elongation factor DmS-II|Drug|false|false||DM IInull|Hypertensive disease|Disorder|false|false||HTNnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate CAnull|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0376358;C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0376358;C0496923;C0154088;C0033575;C0154009|prostatenull|at admission|Finding|false|false||At Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Feeling comfortable|Finding|false|false||comfortablenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Lung|Anatomy|false|false||Lungsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Pansystolic murmur|Finding|false|false||holosystolic murmurnull|Heart murmur|Finding|false|false||murmurnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Awake (finding)|Finding|false|false||Awakenull|Awakening (time frame)|Time|false|false||Awakenull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Mental Recall|Finding|false|false||Recallnull|Recall (activity)|Event|false|false||Recallnull|Physical object|Entity|false|false||objectsnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|Difficult (qualifier value)|Finding|false|false||Difficulty withnull|Has difficulty doing (qualifier value)|Finding|false|false||Difficultynull|Naming (function)|Finding|false|false||Namingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dysarthria|Disorder|true|false||dysarthrianull|error|Modifier|false|false||errorsnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false|C0027740;C0037303;C0010268|Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false|C0027740;C0037303;C0010268|Cranial Nervesnull|Cranial Nerves|Anatomy|false|false|C0004992;C0496937|Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false|C0004992;C0496937|Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false|C0004992;C0496937|Nervesnull|Pupil|Anatomy|false|false||Pupilsnull|Round shape|Modifier|false|false||roundnull|Reactive to light|Finding|false|false||reactive to lightnull|Reactive Therapy|Procedure|false|false||reactivenull|Reactive|Modifier|false|false||reactivenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Visual Fields|Modifier|false|false||Visual fieldsnull|Visual|Finding|false|false||Visualnull|Full|Modifier|false|false||fullnull|Social confrontation skill|Finding|false|false||confrontationnull|Confrontation visual field test|Procedure|false|false||confrontation
null|Confrontation|Procedure|false|false||confrontationnull|examination of extraocular movements|Procedure|false|false||Extraocular movementsnull|Extraocular|Finding|false|false||Extraocularnull|Movement|Finding|false|false||movementsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Nystagmus|Disorder|false|false||nystagmusnull|Roman numeral VII|Finding|false|false|C2338708;C3496273;C3496274|VIInull|Lamina VII of gray matter of spinal cord|Anatomy|false|false|C0445385|VII
null|lobule VII|Anatomy|false|false|C0445385|VII
null|layer VII (Cajal)|Anatomy|false|false|C0445385|VIInull|Face|Anatomy|false|false|C0808080|Facialnull|Facial|Modifier|false|false||Facialnull|Strength (attribute)|Finding|false|false|C0015450|strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Roman numeral VIII|Finding|false|false|C2327388;C0228488|VIII
null|COX8A gene|Finding|false|false|C2327388;C0228488|VIIInull|Lamina VIII of gray matter of spinal cord|Anatomy|false|false|C0445599;C1413661|VIII
null|Cerebellar pyramis|Anatomy|false|false|C0445599;C1413661|VIIInull|outcomes otolaryngology hearing|Finding|false|false||Hearing
null|Hearing finding|Finding|false|false||Hearing
null|Hearing|Finding|false|false||Hearingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Palate|Anatomy|false|false|C0439775|Palatalnull|Elevation procedure|Procedure|false|false|C0700374|elevationnull|Elevation|Modifier|false|false||elevationnull|Symmetrical|Finding|false|false||symmetricalnull|Structure of sternocleidomastoid muscle|Anatomy|false|false||Sternocleidomastoidnull|Structure of trapezius muscle|Anatomy|false|false||trapeziusnull|tongue midline|Finding|false|false|C0040408;C1660780|Tongue midlinenull|Benign neoplasm of tongue|Disorder|false|false|C1660780;C0040408|Tonguenull|Procedure on tongue|Procedure|false|false|C0040408;C1660780|Tonguenull|Tongue|Anatomy|false|false|C3693372;C0872394;C0015644;C0153933|Tonguenull|midline cell component|Anatomy|false|false|C0153933;C0872394;C3693372;C0015644|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Muscular fasciculation|Finding|true|false|C0040408;C1660780|fasciculationsnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Bulk (conceptual)|Drug|false|false||bulk
null|Dietary Fiber|Drug|false|false||bulknull|Dyskinetic syndrome|Disorder|true|false||abnormal movementsnull|Abnormal movement|Finding|true|false||abnormal movementsnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Movement|Finding|true|false||movementsnull|Tremor|Finding|false|false||tremorsnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Full|Modifier|false|false||fullnull|Power (Psychology)|Finding|false|false||powernull|Power|LabModifier|false|false||powernull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Pronator drift|Finding|false|false||pronator driftnull|Gait, Unsteady|Finding|false|false||Gait unsteadynull|Gait|Finding|false|false|C4318744|Gaitnull|Unsteady|Modifier|false|false||unsteadynull|rhomberg test|Procedure|false|false|C4318744|rhomberg testnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0427108;C0016928;C0456984;C1656968;C0022885;C0039593;C0392366|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|General unsteadiness|Finding|false|false|C4318744|unsteadinessnull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Light touch|Finding|false|false||light touchnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Exposed to vibration|Disorder|false|false||vibrationnull|Vibration - treatment|Procedure|false|false||vibrationnull|null|Phenomenon|false|false||vibrationnull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Lower extremity>Toes|Anatomy|false|false||Toes
null|Toes|Anatomy|false|false||Toesnull|Coordination of Benefits - Coordination|Finding|false|false||Coordination
null|Coordinated|Finding|false|false||Coordination
null|Physiologic Coordination|Finding|false|false||Coordinationnull|Heel|Anatomy|false|false||heelnull|Shin|Anatomy|false|false||shinnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Structure of right hand|Anatomy|false|false|C0741992|R handnull|Hand problem|Finding|false|false|C0230370;C4285005;C0018563|handnull|Upper extremity>Hand|Anatomy|false|false|C0741992|hand
null|Hand|Anatomy|false|false|C0741992|handnull|Difficult (qualifier value)|Finding|false|false||Difficulty withnull|Has difficulty doing (qualifier value)|Finding|false|false||Difficultynull|Rapid|Modifier|false|false||rapidnull|Alternating|Finding|false|false||alternatingnull|Movement|Finding|false|false||movementsnull|Structure of right hand|Anatomy|false|false|C0741992|R handnull|Hand problem|Finding|false|false|C4285005;C0018563;C0230370|handnull|Upper extremity>Hand|Anatomy|false|false|C0741992|hand
null|Hand|Anatomy|false|false|C0741992|handnull|At discharge|Time|false|false||AT DISCHARGEnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Pupil|Anatomy|false|false||Pupilsnull|Extraocular|Finding|false|false||EOMsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Cardiac attachment|Finding|false|false|C0018787|Cardiacnull|Heart|Anatomy|false|false|C1314974|Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Pansystolic murmur|Finding|false|false||holosystolic murmurnull|Heart murmur|Finding|false|false||murmurnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Erythema|Disorder|true|false||erythemanull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Awake (finding)|Finding|false|false||Awakenull|Awakening (time frame)|Time|false|false||Awakenull|cooperative|Entity|false|false||cooperativenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Mental Orientation|Finding|false|false||Orientationnull|Orientation, Spatial|Modifier|false|false||Orientation
null|Genomic Orientation|Modifier|false|false||Orientation
null|Orientation|Modifier|false|false||Orientationnull|Oriented to person|Finding|false|false||Oriented to personnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Programming Languages|Finding|false|false||Languagenull|null|Attribute|false|false||Languagenull|Languages|Entity|false|false||Languagenull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Comprehension|Finding|false|false||comprehensionnull|Neoplasm of uncertain or unknown behavior of cranial nerves|Disorder|false|false|C0027740;C0010268;C0037303|Cranial Nerves
null|Benign neoplasm of cranial nerves|Disorder|false|false|C0027740;C0010268;C0037303|Cranial Nervesnull|Cranial Nerves|Anatomy|false|false|C0004992;C0496937|Cranial Nervesnull|Bone structure of cranium|Anatomy|false|false|C0004992;C0496937|Cranialnull|Cranial|Modifier|false|false||Cranialnull|Nerve|Anatomy|false|false|C0004992;C0496937|Nervesnull|Tests (qualifier value)|Finding|false|false||tested
null|Testing|Finding|false|false||testednull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Pronator drift|Finding|true|false||pronator driftnull|Gait|Finding|false|false||Gaitnull|Steady|Modifier|false|false||steadynull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Helping Behavior|Finding|true|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Observation of Sensation|Finding|false|false||Sensation
null|Sensory perception|Finding|false|false||Sensationnull|sensory exam|Procedure|false|false||Sensationnull|Sensation quality|Modifier|false|false||Sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Lower extremity>Toes|Anatomy|false|false||Toes
null|Toes|Anatomy|false|false||Toesnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Glycosylated hemoglobin A|Drug|false|false||HbA1c
null|Glycosylated hemoglobin A|Drug|false|false||HbA1cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1cnull|KCNH1 gene|Finding|false|false||eAGnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CAT scan of head|Procedure|false|false|C0018670;C0152336|CT Headnull|null|Attribute|false|false|C0018670;C0152336|CT Headnull|Problems with head|Disorder|false|false|C0018670;C0152336|Headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|Headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0881943;C0202691;C0362076|Head
null|Head|Anatomy|false|false|C0876917;C0881943;C0202691;C0362076|Headnull|Head Device|Device|false|false||Headnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Focal|Modifier|false|false||foci ofnull|Foci|Finding|false|false||focinull|Focal|Modifier|false|false||focinull|Pathologic calcification, calcified structure|Finding|false|false||calcifications
null|Physiologic calcification|Finding|false|false||calcificationsnull|Calcified (qualifier value)|Modifier|false|false||calcificationsnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Benign Meningioma|Disorder|false|false||meningioma
null|Meningioma|Disorder|false|false||meningiomanull|Hematoma|Finding|false|false||hematomanull|Subacute to chronic|Time|false|false||subacute to chronicnull|Subacute|Time|false|false||subacutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Loss (adaptation)|Finding|false|false||Lossnull|Loss (quantitative)|LabModifier|false|false||Lossnull|Gray color|Modifier|false|false||graynull|Gray unit of radiation dose|LabModifier|false|false||graynull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Cell Differentiation process|Finding|false|false||differentiation
null|Differentiation|Finding|false|false||differentiationnull|Cellular Differentiation Qualifier|Attribute|false|false||differentiationnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|AKT1S1 wt Allele|Finding|false|false|C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0796494|lobenull|lobe|Anatomy|false|false|C0021308;C3539671;C1428707;C0333548;C1547295;C1547229|lobenull|Acute infarct|Finding|false|false|C0796494|acute infarctnull|Admission Level of Care Code - Acute|Finding|false|false|C0796494|acute
null|Acute - Triage Code|Finding|false|false|C0796494|acutenull|acute|Time|false|false||acutenull|Infarction|Finding|false|false|C0796494|infarctnull|MRI of head|Procedure|false|false|C0018670;C0152336|MRI Headnull|CYREN gene|Finding|false|false|C0018670;C0152336|MRInull|Magnetic resonance imaging service|Procedure|false|false|C0018670;C0152336|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C0018670;C0152336|MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false|C0018670;C0152336|Headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|Headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0024485;C0587658;C1824234;C0876917;C0412674;C0362076|Head
null|Head|Anatomy|false|false|C0024485;C0587658;C1824234;C0876917;C0412674;C0362076|Headnull|Head Device|Device|false|false||Headnull|Acute to subacute|Time|false|false||Acute to subacutenull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Subacute|Time|false|false||subacutenull|Bilateral|Modifier|false|false||bilateralnull|Infarction|Finding|false|false||infarctionsnull|Largest|LabModifier|false|false||largestnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|patient appearance regarding mental status exam|Procedure|false|false||Appearancenull|null|Attribute|false|false||Appearancenull|Personal appearance|Subject|false|false||Appearancenull|Appearance|Modifier|false|false||Appearancenull|Kind of quantity - Appearance|LabModifier|false|false||Appearancenull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Somewhat|Finding|false|false||somewhatnull|Heterogeneity|Modifier|false|false||heterogeneousnull|Attention - G-code|Finding|false|false||attention
null|Attention|Finding|false|false||attentionnull|follow-up|Procedure|false|false||followupnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Present|Finding|false|false||presence ofnull|Providing presence (regime/therapy)|Procedure|false|false||presencenull|Presence (property)|Modifier|false|false||presencenull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Meningioma|Disorder|false|false|C0016733;C0549224;C0162783|meningiomasnull|Table Cell Horizontal Align - left|Finding|false|false|C0016733;C0549224;C0162783|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Frontal region|Anatomy|false|false|C0025286;C1514562;C1552822|frontal region
null|frontal lobe|Anatomy|false|false|C0025286;C1514562;C1552822|frontal region
null|Prefrontal Cortex|Anatomy|false|false|C0025286;C1514562;C1552822|frontal regionnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Protein Domain|Drug|false|false|C0016733;C0549224;C0162783|regionnull|Geographic Locations|Entity|false|false||regionnull|regional|Modifier|false|false||regionnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Mass Effect|Finding|true|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Marked|Modifier|false|false||Marked
null|Massive|Modifier|false|false||Markednull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Left Ventricular Hypertrophy|Disorder|false|false|C0018827|left ventricular hypertrophynull|null|Attribute|false|false|C0018827|left ventricular hypertrophynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Ventricular hypertrophy|Disorder|false|false|C0018827|ventricular hypertrophynull|Heart Ventricle|Anatomy|false|false|C3484363;C0340279;C0020564;C0149721|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Hypertrophy|Finding|false|false|C0018827|hypertrophynull|Dental caries|Disorder|false|false|C0333343|cavity
null|Cavitation|Disorder|false|false|C0333343|cavitynull|Body cavities|Anatomy|false|false|C1510420;C0011334|cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Global|Modifier|false|false||global
null|Generalized|Modifier|false|false||globalnull|Systole|Finding|false|false||systolicnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Mild Severity of Illness Code|Finding|false|false|C4533215;C0003501|Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Aortic valve structure|Anatomy|false|false|C1547225|aortic valve
null|Chest>Aortic valve|Anatomy|false|false|C1547225|aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Aortic Valve Insufficiency|Disorder|false|false|C0003483|aortic regurgitationnull|Aorta|Anatomy|false|false|C0460152;C0232605;C2004489;C0003504|aorticnull|Regurgitation|Finding|false|false|C0003483|regurgitation
null|Regurgitates after swallowing|Finding|false|false|C0003483|regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false|C0003483|regurgitationnull|Right Ventricular Free Wall|Anatomy|false|false|C1552823;C0332296|Right ventricular free wallnull|Table Cell Horizontal Align - right|Finding|false|false|C4288280|Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Free of (attribute)|Finding|false|false|C4288280|freenull|Empty (qualifier)|Modifier|false|false||freenull|Walls of a building|Device|false|false||wallnull|Hypertrophy|Finding|false|false||hypertrophynull|Pulmonary artery structure|Anatomy|false|false|C4522268;C0039155;C2707265;C0221155;C0020538|Pulmonary arterynull|Pulmonary (intended site)|Finding|false|false|C0034052;C0226004;C0003842;C0024109|Pulmonarynull|Lung|Anatomy|false|false|C0221155;C2707265;C0020538;C4522268|Pulmonarynull|null|Attribute|false|false|C0024109;C0226004;C0003842;C0034052|Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Arterial system|Anatomy|false|false|C2707265;C0221155;C0039155;C4522268;C0020538|artery
null|Arteries|Anatomy|false|false|C2707265;C0221155;C0039155;C4522268;C0020538|arterynull|Systolic Hypertension|Disorder|false|false|C0024109;C0226004;C0003842;C0034052|systolic hypertensionnull|Systole|Finding|false|false|C0226004;C0003842;C0034052|systolicnull|Hypertensive disease|Disorder|false|false|C0226004;C0003842;C0024109;C0034052|hypertensionnull|Dilated|Finding|false|false||Dilatednull|Ascending aorta structure|Anatomy|false|false|C0869784;C1547175;C1962987|ascending aortanull|Sequencing - Ascending|Finding|false|false|C4037978;C0003483;C0003956|ascending
null|Ascend (action)|Finding|false|false|C4037978;C0003483;C0003956|ascendingnull|Ascending|Modifier|false|false||ascendingnull|Procedure on aorta|Procedure|false|false|C0003956;C4037978;C0003483|aortanull|Chest+Abdomen>Aorta|Anatomy|false|false|C1547175;C1962987;C0869784|aorta
null|Aorta|Anatomy|false|false|C1547175;C1962987;C0869784|aortanull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||CLINICALnull|Clinical|Modifier|false|false||CLINICALnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Aortic Valve Stenosis|Finding|false|false|C0003483|aortic stenosisnull|Aorta|Anatomy|false|false|C0003507|aorticnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Amorphous Calcium Carbonate|Drug|false|false|C2954192;C0152325|ACC
null|Acetyl-CoA Carboxylase 1|Drug|false|false|C2954192;C0152325|ACC
null|Acetyl-CoA Carboxylase 1|Drug|false|false|C2954192;C0152325|ACCnull|Agenesis of corpus callosum|Disorder|false|false|C2954192;C0152325|ACC
null|Aplasia Cutis Congenita|Disorder|false|false|C2954192;C0152325|ACC
null|Adrenocortical carcinoma|Disorder|false|false|C2954192;C0152325|ACCnull|ACACA wt Allele|Finding|false|false|C2954192;C0152325|ACC
null|ACACA gene|Finding|false|false|C2954192;C0152325|ACCnull|Gray matter of anterior cingulate gyrus|Anatomy|false|false|C0002880;C0272325;C3541413;C1412104;C4724142;C3541857;C0206686;C0175754;C0282160|ACC
null|Structure of forceps minor|Anatomy|false|false|C0002880;C0272325;C3541413;C1412104;C4724142;C3541857;C0206686;C0175754;C0282160|ACCnull|acetohydroxamic acid|Drug|false|false||AHA
null|acetohydroxamic acid|Drug|false|false||AHAnull|Factor 8 deficiency, acquired|Disorder|false|false|C2954192;C0152325|AHA
null|Autoimmune hemolytic anemia|Disorder|false|false|C2954192;C0152325|AHAnull|American Hospital Association|Entity|false|false||AHAnull|Heart valve disease|Disorder|false|false|C4037974;C0018787|Valvular Heart Diseasenull|Heart Diseases|Disorder|false|false|C4037974;C0018787|Heart Diseasenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|Heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|Heartnull|Chest>Heart|Anatomy|false|false|C0018824;C0153957;C0153500;C1522577;C0220845;C0162791;C0282423;C0018799;C0012634;C0795691|Heart
null|Heart|Anatomy|false|false|C0018824;C0153957;C0153500;C1522577;C0220845;C0162791;C0282423;C0018799;C0012634;C0795691|Heartnull|Disease|Disorder|false|false|C4037974;C0018787|Diseasenull|Guidelines|Finding|false|false|C4037974;C0018787|Guidelines
null|Guideline (Publication Type)|Finding|false|false|C4037974;C0018787|Guidelines
null|guiding characteristics|Finding|false|false|C4037974;C0018787|Guidelinesnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false|C4037974;C0018787|follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Echocardiography|Procedure|false|false||echocardiogramnull|year|Time|false|false||yearsnull|Endocarditis prophylaxis|Procedure|false|false||endocarditis prophylaxisnull|Endocarditis|Disorder|false|false||endocarditisnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Recommendation|Finding|false|false||recommendationsnull|ECHO protocol|Procedure|false|false||echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false||echonull|Echo <Calopterygidae>|Entity|false|false||echonull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||Clinicalnull|Clinical|Modifier|false|false||Clinicalnull|Decision|Finding|false|false||decisionsnull|Patient need for (contextual qualifier)|Finding|false|false||need fornull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|Data|Finding|false|false||datanull|Data call receiving device|Device|false|false||datanull|Data <Amphipyrinae>|Entity|false|false||datanull|Magnetic resonance angiography of vascular structure of head|Procedure|false|false|C0018670;C0152336;C0027530;C3159206|MRA Headnull|tocilizumab|Drug|false|false|C0018670;C0152336|MRA
null|tocilizumab|Drug|false|false|C0018670;C0152336|MRA
null|tocilizumab|Drug|false|false|C0018670;C0152336|MRAnull|Magnetic Resonance Angiography|Procedure|false|false|C0018670;C0152336;C0027530;C3159206|MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|Problems with head|Disorder|false|false|C0018670;C0152336;C0027530;C3159206|Headnull|Procedure on head|Procedure|false|false|C0018670;C0152336;C0027530;C3159206|Headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0812434;C0684335;C0243032;C1609165;C1636167;C0362076|Head
null|Head|Anatomy|false|false|C0876917;C0812434;C0684335;C0243032;C1609165;C1636167;C0362076|Headnull|Head Device|Device|false|false||Headnull|Passive joint movement of neck (finding)|Finding|false|false|C0018670;C0152336;C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0018670;C0152336;C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0876917;C1636167;C0362076;C0812434;C0684335;C0243032|Neck
null|Neck|Anatomy|false|false|C0876917;C1636167;C0362076;C0812434;C0684335;C0243032|Necknull|Mild Severity of Illness Code|Finding|false|false|C0004811;C0226004;C0003842|Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|atherosclerotic|Finding|false|false|C0004811;C0226004;C0003842|atheroscleroticnull|Disease|Disorder|false|false|C0226004;C0003842;C0004811|diseasenull|Structure of basilar artery|Anatomy|false|false|C0333482;C1547225;C0012634|basilar arterynull|Basilar|Modifier|false|false||basilarnull|Arterial system|Anatomy|false|false|C1547225;C0012634;C0333482|artery
null|Arteries|Anatomy|false|false|C1547225;C0012634;C0333482|arterynull|Evidence of (contextual qualifier)|Finding|false|false|C0005847|evidence ofnull|Evidence|Finding|false|false|C0005847|evidencenull|Admission Level of Care Code - Acute|Finding|false|false|C0005847|acute
null|Acute - Triage Code|Finding|false|false|C0005847|acutenull|acute|Time|false|false||acutenull|Abnormality of the vasculature|Finding|false|false|C0005847|vascular abnormalitiesnull|Blood Vessel|Anatomy|false|false|C0241657;C1547295;C1547229;C0332120;C0000768;C3887511;C0000769|vascularnull|Vascular|Modifier|false|false||vascularnull|Congenital Abnormality|Disorder|false|false|C0005847|abnormalitiesnull|teratologic|Finding|false|false|C0005847|abnormalitiesnull|Intracranial Route of Administration|Finding|false|false|C0524466;C0226004;C0003842|intracranialnull|Intracranial|Anatomy|false|false|C0397581;C1522213|intracranialnull|Procedure on artery|Procedure|false|false|C0226004;C0003842;C0524466|arteriesnull|Arteries|Anatomy|false|false|C0397581;C1522213|arteries
null|Arterial system|Anatomy|false|false|C0397581;C1522213|arteriesnull|Neurosurgical service|Entity|false|false||neurosurgical servicenull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Encounter Referral Source - emergency room|Finding|false|false||emergency roomnull|Accident and Emergency department|Device|false|false||emergency roomnull|Accident and Emergency department|Entity|false|false||emergency roomnull|Level of Care - Emergency|Finding|false|false||emergency
null|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Series|LabModifier|false|false||seriesnull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|More|LabModifier|false|false||morenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Parietal|Modifier|false|false||parietalnull|AKT1S1 wt Allele|Finding|false|false|C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0796494|lobenull|lobe|Anatomy|false|false|C1552822;C3539671;C1428707|lobenull|Table Cell Horizontal Align - left|Finding|false|false|C0796494|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Recent|Time|false|false||recentnull|Accidental Falls|Disorder|false|false||fallsnull|Falls|Finding|false|false||fallsnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Scale, LOINC Axis 5|Finding|false|false|C0222045|scale
null|Base Number|Finding|false|false|C0222045|scale
null|Scale - rank|Finding|false|false|C0222045|scalenull|Integumentary scale|Anatomy|false|false|C1947916;C0349674;C2981742;C1522412|scalenull|Weight measurement scales|Device|false|false||scalenull|Scaling|Event|false|false|C0222045|scalenull|Concern|Finding|false|false||concernnull|Hypoglycemia|Disorder|false|false||hypoglycemianull|Blood glucose below reference range (finding)|Finding|false|false||hypoglycemianull|General unsteadiness|Finding|false|false||unsteadinessnull|CYREN gene|Finding|false|false|C0018670;C0152336|MRInull|Magnetic resonance imaging service|Procedure|false|false|C0018670;C0152336|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C0018670;C0152336|MRInull|Maori Language|Entity|false|false||MRInull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917;C0024485;C0587658;C1824234|head
null|Head|Anatomy|false|false|C0362076;C0876917;C0024485;C0587658;C1824234|headnull|Head Device|Device|false|false||headnull|Benign Meningioma|Disorder|false|false||meningioma
null|Meningioma|Disorder|false|false||meningiomanull|malignant neoplasm of frontal lobe|Disorder|false|false|C0016733;C0796494|frontal lobenull|frontal lobe|Anatomy|false|false|C0153635;C3539671;C1428707;C0021308|frontal lobenull|Coronal (qualifier value)|Modifier|false|false||frontalnull|AKT1S1 wt Allele|Finding|false|false|C0016733;C0796494|lobe
null|AKT1S1 gene|Finding|false|false|C0016733;C0796494|lobenull|lobe|Anatomy|false|false|C3539671;C1428707;C0153635|lobenull|Infarction|Finding|false|false|C0016733|infarctnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Encounter Referral Source - emergency room|Finding|false|false||emergency roomnull|Accident and Emergency department|Device|false|false||emergency roomnull|Accident and Emergency department|Entity|false|false||emergency roomnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Day hospital|Device|false|false||hospital daynull|Day hospital|Entity|false|false||hospital daynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Nearly|Modifier|false|false||nearlynull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Neurology speciality|Title|false|false||neurologynull|Consultation|Procedure|false|false||consultnull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Dilantin|Drug|false|false||dilantin
null|Dilantin|Drug|false|false||dilantinnull|null|Event|false|false||checkingnull|Electroencephalography|Procedure|false|false||EEGnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Surface|Modifier|false|false||surfacenull|ECHO protocol|Procedure|false|false|C4266577;C0006104|echo
null|Extension for Community Healthcare Outcomes|Procedure|false|false|C4266577;C0006104|echonull|Echo <Calopterygidae>|Entity|false|false||echonull|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRA
null|tocilizumab|Drug|false|false||MRAnull|Magnetic Resonance Angiography|Procedure|false|false|C0027530;C3159206;C4266577;C0006104|MRAnull|MRI-Based Angiogram|Lab|false|false||MRAnull|Brain Diseases|Disorder|false|false|C4266577;C0006104;C0027530;C3159206|brainnull|Head>Brain|Anatomy|false|false|C0006111;C0812434;C0684335;C5575284;C0058928;C0243032|brain
null|Brain|Anatomy|false|false|C0006111;C0812434;C0684335;C5575284;C0058928;C0243032|brainnull|Passive joint movement of neck (finding)|Finding|false|false|C4266577;C0006104;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C4266577;C0006104;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0243032;C0006111;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0243032;C0006111;C0812434;C0684335|necknull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Embolism|Finding|false|false||embolicnull|Nature|Finding|false|false||nature
null|Natures|Finding|false|false||naturenull|Cerebrovascular accident|Disorder|false|false||strokesnull|Neurology speciality|Title|false|false||Neurologynull|3 Months|Time|false|false||3 monthsnull|month|Time|false|false||monthsnull|Repeat Object|Finding|false|false|C0018670;C0152336|repeat
null|Repeat|Finding|false|false|C0018670;C0152336|repeatnull|Repeat Pattern|Time|false|false||repeatnull|MRI of head|Procedure|false|false|C0018670;C0152336|head MRInull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0024485;C0587658;C0876917;C1705914;C0205341;C0412674;C1824234|head
null|Head|Anatomy|false|false|C0362076;C0024485;C0587658;C0876917;C1705914;C0205341;C0412674;C1824234|headnull|Head Device|Device|false|false||headnull|CYREN gene|Finding|false|false|C0018670;C0152336|MRInull|Magnetic resonance imaging service|Procedure|false|false|C0018670;C0152336|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C0018670;C0152336|MRInull|Maori Language|Entity|false|false||MRInull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|glipizide|Drug|false|false||glipizide
null|glipizide|Drug|false|false||glipizidenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Episode of|Time|false|false||episodesnull|Hypoglycemia|Disorder|false|false||hypoglycemianull|Blood glucose below reference range (finding)|Finding|false|false||hypoglycemianull|Neurologic (qualifier value)|Modifier|false|false||neurologicnull|In-House|Finding|false|false||in-housenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Right hemiparesis|Finding|false|false||right sided weaknessnull|Right sided|Modifier|false|false||right sided
null|Right|Modifier|false|false||right sidednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|General unsteadiness|Finding|false|false||unsteadinessnull|Continuous|Finding|false|false||continuednull|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||support
null|Support brand of multivitamin|Drug|false|false||supportnull|Supportive assistance|Finding|false|false||supportnull|Supportive care|Procedure|false|false||supportnull|Support - dental|Attribute|false|false||supportnull|null|Device|false|false||supportnull|short-term|Time|false|false||short termnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Term (lexical)|Finding|false|false||term
null|Term Birth|Finding|false|false||termnull|Term (temporal)|Time|false|false||termnull|Rehabilitation therapy|Procedure|false|false||rehabnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|transfers|Finding|false|false||transfersnull|Ambulate|Finding|false|false||ambulatenull|Walkers|Device|false|false||walkernull|Neurology speciality|Title|false|false||neurologynull|Neurosurgical Procedures|Procedure|false|false||neurosurgerynull|Science of neurosurgery|Title|false|false||neurosurgerynull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Ischemic stroke|Disorder|false|false||ischemic strokesnull|Ischemic|Finding|false|false||ischemicnull|Cerebrovascular accident|Disorder|false|false||strokesnull|Benign Meningioma|Disorder|false|false||meningioma
null|Meningioma|Disorder|false|false||meningiomanull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Prandin|Drug|false|false||prandin
null|Prandin|Drug|false|false||prandinnull|glipizide|Drug|false|false||glipizide
null|glipizide|Drug|false|false||glipizidenull|isosorbide|Drug|false|false||isosorbide
null|isosorbide|Drug|false|false||isosorbidenull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|allopurinol|Drug|false|false||allopurinol
null|allopurinol|Drug|false|false||allopurinolnull|torsemide|Drug|false|false||torsemide
null|torsemide|Drug|false|false||torsemidenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Lipitor|Drug|false|false||lipitor
null|Lipitor|Drug|false|false||lipitornull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|isosorbide dinitrate|Drug|false|false||Isosorbide Dinitrate
null|isosorbide dinitrate|Drug|false|false||Isosorbide Dinitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||Dailynull|torsemide|Drug|false|false||Torsemide
null|torsemide|Drug|false|false||Torsemidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|glipizide|Drug|false|false||Glipizide
null|glipizide|Drug|false|false||Glipizidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Benign Meningioma|Disorder|false|false||meningioma
null|Meningioma|Disorder|false|false||meningiomanull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Parietal|Modifier|false|false||parietalnull|Infarction|Finding|false|false||infarctnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Confusion|Disorder|false|false||Confusednull|Precaution Code - Confused|Finding|false|false||Confused
null|Clouded consciousness|Finding|false|false||Confusednull|Sometimes|Time|false|false||sometimesnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Small|LabModifier|false|false||smallnull|Cerebrovascular accident|Disorder|false|false|C4266577;C0006104|strokenull|Stroke (heart beat)|Finding|false|false|C4266577;C0006104|strokenull|LEFT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE LEFT SIDE OF THE BODY)|Modifier|false|false||left side
null|Left|Modifier|false|false||left sidenull|Table Cell Horizontal Align - left|Finding|false|false|C4266577;C0006104|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Side|Modifier|false|false||sidenull|Brain Diseases|Disorder|false|false|C4266577;C0006104|brainnull|Head>Brain|Anatomy|false|false|C0006111;C0038454;C5977286;C1552822|brain
null|Brain|Anatomy|false|false|C0006111;C0038454;C5977286;C1552822|brainnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|General Instructions|Finding|false|false||General Instructionsnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Acknowledgement Detail Type - Information|Finding|false|false||Information
null|Error severity - Information|Finding|false|false||Information
null|Information|Finding|false|false||Information
null|control act - information|Finding|false|false||Informationnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Exercise|Finding|false|false||Exercisenull|Exercise Pain Management|Procedure|false|false||Exercisenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Lifting|Event|true|false||liftingnull|Straining (finding)|Finding|true|false||strainingnull|Excessive (qualifier value)|Modifier|false|false||excessivenull|Decompression Sickness|Disorder|false|false||bendingnull|Bending - Changing basic body position|Finding|false|false||bending
null|Does bend|Finding|false|false||bendingnull|Bent|Modifier|false|false||bendingnull|Intake|Finding|false|false|C1304649|intakenull|Measurement of fluid intake|Procedure|false|false|C1304649|intake
null|Intake (treatment)|Procedure|false|false|C1304649|intakenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fibernull|Tissue fiber|Anatomy|false|false|C0225326;C1321801;C4521161;C3251814;C1512806|fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Constipation|Finding|false|false||constipationnull|Drugs, Non-Prescription|Drug|false|false||over the counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Anti-Inflammatory Agents|Drug|false|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|false|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Etc.|Finding|false|false||etcnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0872393;C0038354;C0496905;C0153943;C0154060;C0577027|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0872393;C0038354;C0496905;C0153943;C0154060;C0577027|stomach
null|Stomach|Anatomy|false|false|C0872393;C0038354;C0496905;C0153943;C0154060;C0577027|stomachnull|Prilosec|Drug|false|false||Prilosec
null|Prilosec|Drug|false|false||Prilosecnull|Protonix|Drug|false|false||Protonix
null|Protonix|Drug|false|false||Protonixnull|Pepcid|Drug|false|false||Pepcid
null|Pepcid|Drug|false|false||Pepcidnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Stomach Diseases|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Benign neoplasm of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomach
null|Carcinoma in situ of stomach|Disorder|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach problem|Finding|false|false|C3714551;C0038351;C4266636|stomachnull|Procedure on stomach|Procedure|false|false|C3714551;C0038351;C4266636|stomachnull|Stomach structure|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomach
null|Abdomen>Stomach|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomach
null|Stomach|Anatomy|false|false|C0872393;C0577027;C0038354;C0496905;C0153943;C0154060|stomachnull|Have Vulvar Irritation question|Finding|false|false||irritation
null|Irritability - emotion|Finding|false|false||irritation
null|Irritation (finding)|Finding|false|false||irritationnull|Irritation|Phenomenon|false|false||irritationnull|Make - Instruction Imperative|Finding|false|false||Make
null|Manufacturer Name|Finding|false|false||Makenull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glassnull|Chromosome 2q32-Q33 Deletion Syndrome|Disorder|false|false||glassnull|Glass Packaging Device|Device|false|false||glass
null|Glass (substance)|Device|false|false||glassnull|cow milk allergenic extract|Drug|false|false||milk
null|Milk antigen|Drug|false|false||milk
null|Milk Beverage|Drug|false|false||milk
null|Plant-Based Milk|Drug|false|false||milk
null|cow milk allergenic extract|Drug|false|false||milk
null|Milk Specimen|Drug|false|false||milk
null|Cow's milk|Drug|false|false||milk
null|null|Drug|false|false||milknull|Milk (body substance)|Finding|false|false||milk
null|Milk Specimen Code|Finding|false|false||milknull|Clearance procedure|Procedure|false|false||Clearancenull|Clearance of substance|Attribute|false|false||Clearancenull|Clearance [PK]|Phenomenon|false|false||Clearancenull|Clearance|Modifier|false|false||Clearancenull|Work|Event|false|false||worknull|Postoperative Period|Time|false|false||post-operativenull|Office Visits|Procedure|false|false||office visitnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Visit|Finding|false|false||visitnull|Make - Instruction Imperative|Finding|false|false||Make
null|Manufacturer Name|Finding|false|false||Makenull|SURE Test|Finding|false|false||surenull|Certain (qualifier value)|Modifier|false|false||surenull|Continuous|Finding|false|false||continuenull|Incentive spirometry|Procedure|false|false||incentive spirometernull|Incentive Spirometers (device)|Device|false|false||incentive spirometernull|Incentives|Modifier|false|false||incentivenull|Spirometer Device|Device|false|false||spirometernull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Call - dosing instruction fragment|Finding|false|false||CALL
null|Call (Instruction)|Finding|false|false||CALL
null|Decision|Finding|false|false||CALL
null|CHL1 gene|Finding|false|false||CALLnull|null|Attribute|false|false||SURGEONnull|Surgeon|Subject|false|false||SURGEONnull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Experience (Practice)|Finding|false|false||EXPERIENCE
null|Experience|Finding|false|false||EXPERIENCEnull|Following|Time|false|false||FOLLOWING
null|Status post|Time|false|false||FOLLOWINGnull|new onset|Finding|false|false||New onsetnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Tremor|Finding|false|false||tremorsnull|Seizures|Finding|false|false||seizuresnull|Confusion|Disorder|true|false||confusionnull|Clouded consciousness|Finding|true|false||confusionnull|Mental status changes|Finding|false|false||change in mental statusnull|null|Attribute|false|false||change in mental statusnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Changed status|LabModifier|false|false||change
null|Delta (difference)|LabModifier|false|false||changenull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Paresthesia|Disorder|false|false|C0278454;C0015385|tinglingnull|Has tingling sensation|Finding|false|false||tinglingnull|Weakness|Finding|false|false|C0278454;C0015385|weakness
null|Asthenia|Finding|false|false|C0278454;C0015385|weaknessnull|All extremities|Anatomy|false|false|C0030554;C3714552;C0004093|extremities
null|Limb structure|Anatomy|false|false|C0030554;C3714552;C0004093|extremitiesnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Headache|Finding|false|false||headachenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than or Equal To|LabModifier|false|false||greater than or equal tonull|Greater Than or Equal To|LabModifier|false|false||greater than or equalnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Equal|Modifier|false|false||equal tonull|Relational Operator - Equal|Finding|false|false||equalnull|Equal|Modifier|false|false||equalnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions