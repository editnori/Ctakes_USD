 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
CARDIOTHORACIC|156,170
<EOL>|170,171
<EOL>|172,173
lisinopril|185,195
<EOL>|195,196
<EOL>|197,198
Attending|198,207
:|207,208
_|209,210
_|210,211
_|211,212
<EOL>|212,213
<EOL>|214,215
Substernal|232,242
chest|243,248
pain|249,253
and|254,257
throat|258,264
tightness|265,274
with|275,279
exertion|280,288
<EOL>|288,289
<EOL>|289,290
<EOL>|291,292
Major|292,297
Surgical|298,306
or|307,309
Invasive|310,318
Procedure|319,328
:|328,329
<EOL>|329,330
_|330,331
_|331,332
_|332,333
<EOL>|333,334
1.|334,336
Off|337,340
pump|341,345
coronary|346,354
artery|355,361
bypass|362,368
graft|369,374
x3|375,377
,|377,378
left|379,383
internal|384,392
<EOL>|393,394
mammary|394,401
artery|402,408
to|409,411
left|412,416
anterior|417,425
descending|426,436
artery|437,443
and|444,447
saphenous|448,457
<EOL>|458,459
vein|459,463
grafts|464,470
to|471,473
diagonal|474,482
,|482,483
and|484,487
obtuse|488,494
marginal|495,503
arteries|504,512
.|512,513
<EOL>|513,514
2.|514,516
Endoscopic|517,527
harvesting|528,538
of|539,541
the|542,545
long|546,550
saphenous|551,560
vein|561,565
.|565,566
<EOL>|566,567
<EOL>|567,568
<EOL>|569,570
This|598,602
is|603,605
a|606,607
_|608,609
_|609,610
_|610,611
patient|612,619
with|620,624
extensive|625,634
coronary|635,643
artery|644,650
<EOL>|651,652
disease|652,659
history|660,667
with|668,672
previous|673,681
stenting|682,690
presented|691,700
again|701,706
with|707,711
<EOL>|712,713
symptoms|713,721
and|722,725
was|726,729
investigated|730,742
and|743,746
found|747,752
to|753,755
have|756,760
a|761,762
significant|763,774
<EOL>|775,776
lesion|776,782
in|783,785
the|786,789
left|790,794
anterior|795,803
descending|804,814
artery|815,821
diagonal|822,830
and|831,834
the|835,838
<EOL>|839,840
obtuse|840,846
marginal|847,855
arteries|856,864
.|864,865
Left|867,871
ventricular|872,883
function|884,892
is|893,895
well|896,900
<EOL>|901,902
preserved|902,911
and|912,915
she|916,919
was|920,923
electively|924,934
admitted|935,943
for|944,947
off|948,951
pump|952,956
coronary|957,965
<EOL>|966,967
artery|967,973
bypass|974,980
grafting|981,989
.|989,990
<EOL>|990,991
<EOL>|991,992
<EOL>|993,994
Coronary|1016,1024
artery|1025,1031
disease|1032,1039
(|1039,1040
s|1040,1041
/|1041,1042
p|1042,1043
MI|1044,1046
_|1047,1048
_|1048,1049
_|1049,1050
,|1050,1051
BMS|1052,1055
to|1056,1058
proximal|1059,1067
LAD|1068,1071
_|1072,1073
_|1073,1074
_|1074,1075
,|1075,1076
<EOL>|1077,1078
DES|1078,1081
to|1082,1084
mid|1085,1088
LAD|1089,1092
_|1093,1094
_|1094,1095
_|1095,1096
,|1096,1097
DES|1098,1101
to|1102,1104
edge|1105,1109
ISR|1110,1113
of|1114,1116
mid|1117,1120
LAD|1121,1124
DES|1125,1128
and|1129,1132
stenosis|1133,1141
<EOL>|1142,1143
distal|1143,1149
to|1150,1152
stent|1153,1158
_|1159,1160
_|1160,1161
_|1161,1162
,|1162,1163
DES|1164,1167
to|1168,1170
OM1|1171,1174
,|1174,1175
_|1176,1177
_|1177,1178
_|1178,1179
.|1179,1180
<EOL>|1181,1182
diastolic|1182,1191
congestive|1192,1202
heart|1203,1208
failure|1209,1216
<EOL>|1216,1217
Hypertension|1217,1229
<EOL>|1229,1230
Dyslipidemia|1230,1242
<EOL>|1242,1243
Morbid|1243,1249
obesity|1250,1257
<EOL>|1257,1258
COPD|1258,1262
<EOL>|1262,1263
GERD|1263,1267
<EOL>|1267,1268
Rt|1268,1270
rotator|1271,1278
cuff|1279,1283
injury|1284,1290
/|1290,1291
bursitis|1291,1299
(|1299,1300
outpt|1300,1305
_|1306,1307
_|1307,1308
_|1308,1309
,|1309,1310
<EOL>|1311,1312
Migraines|1312,1321
,|1321,1322
<EOL>|1323,1324
Depression|1324,1334
/|1334,1335
Anxiety|1335,1342
<EOL>|1342,1343
DJD|1343,1346
<EOL>|1346,1347
Hemorrhoids|1347,1358
<EOL>|1359,1360
Rosacea|1360,1367
<EOL>|1368,1369
Left|1369,1373
foot|1374,1378
tendion|1379,1386
repair|1387,1393
<EOL>|1393,1394
<EOL>|1395,1396
:|1410,1411
<EOL>|1411,1412
_|1412,1413
_|1413,1414
_|1414,1415
<EOL>|1415,1416
:|1430,1431
<EOL>|1431,1432
She|1432,1435
was|1436,1439
a|1440,1441
ward|1442,1446
of|1447,1449
the|1450,1453
_|1454,1455
_|1455,1456
_|1456,1457
and|1458,1461
does|1462,1466
not|1467,1470
know|1471,1475
her|1476,1479
family|1480,1486
.|1486,1487
<EOL>|1489,1490
<EOL>|1490,1491
<EOL>|1492,1493
<EOL>|1507,1508
Pulse|1523,1528
:|1528,1529
86|1530,1532
Resp|1533,1537
:|1537,1538
20|1538,1540
O2|1542,1544
sat|1545,1548
:|1548,1549
98|1549,1551
%|1551,1552
<EOL>|1552,1553
B|1553,1554
/|1554,1555
P|1555,1556
Right|1558,1563
:|1563,1564
132|1565,1568
/|1568,1569
68|1569,1571
Left|1574,1578
:|1578,1579
<EOL>|1579,1580
Height|1580,1586
:|1586,1587
5|1588,1589
'|1589,1590
2|1590,1591
Weight|1595,1601
:|1601,1602
210|1602,1605
<EOL>|1606,1607
<EOL>|1607,1608
General|1608,1615
:|1615,1616
AAOx3|1617,1622
,|1622,1623
NAD|1624,1627
<EOL>|1628,1629
Skin|1629,1633
:|1633,1634
Dry|1635,1638
[|1639,1640
x|1640,1641
]|1641,1642
intact|1643,1649
[|1650,1651
x|1651,1652
]|1652,1653
<EOL>|1653,1654
HEENT|1654,1659
:|1659,1660
PERRLA|1661,1667
[|1668,1669
x|1669,1670
]|1670,1671
EOMI|1672,1676
[|1677,1678
x|1678,1679
]|1679,1680
<EOL>|1680,1681
Neck|1681,1685
:|1685,1686
Supple|1688,1694
[|1695,1696
x|1696,1697
]|1697,1698
Full|1699,1703
ROM|1704,1707
[|1708,1709
x|1709,1710
]|1710,1711
<EOL>|1711,1712
Chest|1712,1717
:|1717,1718
Lungs|1719,1724
clear|1725,1730
bilaterally|1731,1742
[|1743,1744
x|1744,1745
]|1745,1746
<EOL>|1746,1747
Heart|1747,1752
:|1752,1753
RRR|1754,1757
[|1758,1759
x|1759,1760
]|1760,1761
Irregular|1763,1772
[|1773,1774
]|1774,1775
Murmur|1777,1783
[|1784,1785
]|1785,1786
grade|1787,1792
_|1793,1794
_|1794,1795
_|1795,1796
_|1796,1797
_|1797,1798
_|1798,1799
<EOL>|1799,1800
Abdomen|1800,1807
:|1807,1808
Soft|1809,1813
[|1814,1815
x|1815,1816
]|1816,1817
non-distended|1817,1830
[|1831,1832
x|1832,1833
]|1833,1834
non-tender|1834,1844
[|1845,1846
x|1846,1847
]|1847,1848
bowel|1848,1853
sounds|1854,1860
<EOL>|1861,1862
+|1862,1863
[|1863,1864
x|1864,1865
]|1865,1866
<EOL>|1866,1867
Extremities|1867,1878
:|1878,1879
Warm|1880,1884
[|1885,1886
x|1886,1887
]|1887,1888
,|1888,1889
well|1890,1894
-|1894,1895
perfused|1895,1903
[|1904,1905
x|1905,1906
]|1906,1907
Edema|1909,1914
[|1915,1916
]|1916,1917
_|1918,1919
_|1919,1920
_|1920,1921
_|1921,1922
_|1922,1923
<EOL>|1923,1924
Varicosities|1924,1936
:|1936,1937
None|1938,1942
[|1943,1944
x|1944,1945
]|1945,1946
<EOL>|1946,1947
Neuro|1947,1952
:|1952,1953
Grossly|1954,1961
intact|1962,1968
[|1969,1970
x|1970,1971
]|1971,1972
<EOL>|1972,1973
<EOL>|1973,1974
Pulses|1974,1980
:|1980,1981
<EOL>|1981,1982
Femoral|1982,1989
Right|1995,2000
:|2000,2001
+|2002,2003
2|2003,2004
Left|2006,2010
:|2010,2011
+|2011,2012
2|2012,2013
<EOL>|2013,2014
DP|2014,2016
Right|2027,2032
:|2032,2033
+|2033,2034
2|2034,2035
Left|2038,2042
:|2042,2043
+|2043,2044
2|2044,2045
<EOL>|2045,2046
_|2046,2047
_|2047,2048
_|2048,2049
Right|2060,2065
:|2065,2066
+|2066,2067
2|2067,2068
Left|2071,2075
:|2075,2076
+|2076,2077
2|2077,2078
<EOL>|2078,2079
Radial|2079,2085
Right|2092,2097
:|2097,2098
cath|2098,2102
site|2103,2107
Left|2109,2113
:|2113,2114
+|2114,2115
2|2115,2116
<EOL>|2116,2117
<EOL>|2117,2118
Carotid|2118,2125
Bruit|2126,2131
:|2131,2132
None|2133,2137
<EOL>|2143,2144
<EOL>|2144,2145
<EOL>|2146,2147
Pertinent|2147,2156
Results|2157,2164
:|2164,2165
<EOL>|2165,2166
Echocargiogram|2166,2180
_|2181,2182
_|2182,2183
_|2183,2184
<EOL>|2184,2185
LEFT|2185,2189
ATRIUM|2190,2196
:|2196,2197
Normal|2198,2204
LA|2205,2207
size|2208,2212
.|2212,2213
<EOL>|2214,2215
RIGHT|2215,2220
ATRIUM|2221,2227
/|2227,2228
INTERATRIAL|2228,2239
SEPTUM|2240,2246
:|2246,2247
Normal|2248,2254
RA|2255,2257
size|2258,2262
.|2262,2263
A|2264,2265
catheter|2266,2274
or|2275,2277
<EOL>|2278,2279
pacing|2279,2285
wire|2286,2290
is|2291,2293
seen|2294,2298
in|2299,2301
the|2302,2305
RA|2306,2308
and|2309,2312
extending|2313,2322
into|2323,2327
the|2328,2331
RV|2332,2334
.|2334,2335
<EOL>|2336,2337
Left|2337,2341
-|2341,2342
to|2342,2344
-|2344,2345
right|2345,2350
shunt|2351,2356
across|2357,2363
the|2364,2367
interatrial|2368,2379
septum|2380,2386
at|2387,2389
rest|2390,2394
.|2394,2395
<EOL>|2396,2397
LEFT|2397,2401
VENTRICLE|2402,2411
:|2411,2412
Wall|2413,2417
thickness|2418,2427
and|2428,2431
cavity|2432,2438
_|2439,2440
_|2440,2441
_|2441,2442
were|2443,2447
<EOL>|2448,2449
obtained|2449,2457
from|2458,2462
2D|2463,2465
images|2466,2472
.|2472,2473
Normal|2474,2480
regional|2481,2489
LV|2490,2492
systolic|2493,2501
function|2502,2510
.|2510,2511
<EOL>|2512,2513
Overall|2513,2520
normal|2521,2527
LVEF|2528,2532
(|2533,2534
>|2534,2535
55|2535,2537
%|2537,2538
)|2538,2539
.|2539,2540
<EOL>|2541,2542
RIGHT|2542,2547
VENTRICLE|2548,2557
:|2557,2558
Normal|2559,2565
RV|2566,2568
chamber|2569,2576
size|2577,2581
and|2582,2585
free|2586,2590
wall|2591,2595
motion|2596,2602
.|2602,2603
<EOL>|2604,2605
AORTA|2605,2610
:|2610,2611
Normal|2612,2618
diameter|2619,2627
of|2628,2630
aorta|2631,2636
at|2637,2639
the|2640,2643
sinus|2644,2649
,|2649,2650
ascending|2651,2660
and|2661,2664
arch|2665,2669
<EOL>|2670,2671
levels|2671,2677
.|2677,2678
Simple|2679,2685
atheroma|2686,2694
in|2695,2697
ascending|2698,2707
aorta|2708,2713
.|2713,2714
Normal|2715,2721
descending|2722,2732
<EOL>|2733,2734
aorta|2734,2739
diameter|2740,2748
.|2748,2749
Simple|2750,2756
atheroma|2757,2765
in|2766,2768
descending|2769,2779
aorta|2780,2785
.|2785,2786
<EOL>|2787,2788
AORTIC|2788,2794
VALVE|2795,2800
:|2800,2801
Normal|2802,2808
aortic|2809,2815
valve|2816,2821
leaflets|2822,2830
(|2831,2832
3|2832,2833
)|2833,2834
.|2834,2835
No|2836,2838
AS|2839,2841
.|2841,2842
No|2843,2845
AR|2846,2848
.|2848,2849
<EOL>|2850,2851
MITRAL|2851,2857
VALVE|2858,2863
:|2863,2864
Normal|2865,2871
mitral|2872,2878
valve|2879,2884
leaflets|2885,2893
with|2894,2898
trivial|2899,2906
MR|2907,2909
.|2909,2910
<EOL>|2911,2912
_|2912,2913
_|2913,2914
_|2914,2915
VALVE|2916,2921
:|2921,2922
Normal|2923,2929
tricuspid|2930,2939
valve|2940,2945
leaflets|2946,2954
with|2955,2959
trivial|2960,2967
<EOL>|2968,2969
TR|2969,2971
.|2971,2972
<EOL>|2973,2974
PULMONIC|2974,2982
VALVE|2983,2988
/|2988,2989
PULMONARY|2989,2998
ARTERY|2999,3005
:|3005,3006
Normal|3007,3013
pulmonic|3014,3022
valve|3023,3028
leaflet|3029,3036
.|3036,3037
<EOL>|3038,3039
No|3039,3041
PS|3042,3044
.|3044,3045
Physiologic|3046,3057
PR|3058,3060
.|3060,3061
<EOL>|3062,3063
PERICARDIUM|3063,3074
:|3074,3075
No|3076,3078
pericardial|3079,3090
effusion|3091,3099
.|3099,3100
<EOL>|3101,3102
Conclusions|3102,3113
<EOL>|3115,3116
Pre|3116,3119
operative|3120,3129
:|3129,3130
<EOL>|3130,3131
The|3131,3134
left|3135,3139
atrium|3140,3146
is|3147,3149
normal|3150,3156
in|3157,3159
size|3160,3164
.|3164,3165
There|3166,3171
is|3172,3174
a|3175,3176
small|3177,3182
PFO|3183,3186
with|3187,3191
a|3192,3193
<EOL>|3194,3195
left|3195,3199
-|3199,3200
to|3200,3202
-|3202,3203
right|3203,3208
shunt|3209,3214
across|3215,3221
the|3222,3225
interatrial|3226,3237
septum|3238,3244
.|3244,3245
Regional|3246,3254
left|3255,3259
<EOL>|3260,3261
ventricular|3261,3272
wall|3273,3277
motion|3278,3284
is|3285,3287
normal|3288,3294
.|3294,3295
Overall|3296,3303
left|3304,3308
ventricular|3309,3320
<EOL>|3321,3322
systolic|3322,3330
function|3331,3339
is|3340,3342
normal|3343,3349
(|3350,3351
LVEF|3351,3355
>|3355,3356
55|3356,3358
%|3358,3359
)|3359,3360
.|3360,3361
Right|3362,3367
ventricular|3368,3379
<EOL>|3380,3381
chamber|3381,3388
size|3389,3393
and|3394,3397
free|3398,3402
wall|3403,3407
motion|3408,3414
are|3415,3418
normal|3419,3425
.|3425,3426
The|3427,3430
diameters|3431,3440
of|3441,3443
<EOL>|3444,3445
aorta|3445,3450
at|3451,3453
the|3454,3457
sinus|3458,3463
,|3463,3464
ascending|3465,3474
and|3475,3478
arch|3479,3483
levels|3484,3490
are|3491,3494
normal|3495,3501
.|3501,3502
There|3503,3508
<EOL>|3509,3510
are|3510,3513
simple|3514,3520
atheroma|3521,3529
in|3530,3532
the|3533,3536
ascending|3537,3546
aorta|3547,3552
.|3552,3553
There|3554,3559
are|3560,3563
simple|3564,3570
<EOL>|3571,3572
atheroma|3572,3580
in|3581,3583
the|3584,3587
descending|3588,3598
thoracic|3599,3607
aorta|3608,3613
.|3613,3614
The|3615,3618
aortic|3619,3625
valve|3626,3631
<EOL>|3632,3633
leaflets|3633,3641
(|3642,3643
3|3643,3644
)|3644,3645
appear|3646,3652
structurally|3653,3665
normal|3666,3672
with|3673,3677
good|3678,3682
leaflet|3683,3690
<EOL>|3691,3692
excursion|3692,3701
and|3702,3705
no|3706,3708
aortic|3709,3715
stenosis|3716,3724
or|3725,3727
aortic|3728,3734
regurgitation|3735,3748
.|3748,3749
The|3750,3753
<EOL>|3754,3755
mitral|3755,3761
valve|3762,3767
appears|3768,3775
structurally|3776,3788
normal|3789,3795
with|3796,3800
trivial|3801,3808
mitral|3809,3815
<EOL>|3816,3817
regurgitation|3817,3830
.|3830,3831
There|3832,3837
is|3838,3840
no|3841,3843
pericardial|3844,3855
effusion|3856,3864
.|3864,3865
<EOL>|3866,3867
<EOL>|3867,3868
Chest|3868,3873
X-Ray|3874,3879
_|3880,3881
_|3881,3882
_|3882,3883
<EOL>|3884,3885
There|3885,3890
is|3891,3893
mild|3894,3898
-|3898,3899
to|3899,3901
-|3901,3902
moderate|3902,3910
cardiomegaly|3911,3923
.|3923,3924
Bilateral|3926,3935
pleural|3936,3943
<EOL>|3944,3945
effusions|3945,3954
are|3955,3958
<EOL>|3959,3960
small|3960,3965
.|3965,3966
Aside|3968,3973
from|3974,3978
atelectasis|3979,3990
in|3991,3993
the|3994,3997
left|3998,4002
lower|4003,4008
lobe|4009,4013
,|4013,4014
the|4015,4018
lungs|4019,4024
<EOL>|4025,4026
are|4026,4029
grossly|4030,4037
clear|4038,4043
.|4043,4044
Almost|4046,4052
complete|4053,4061
resolution|4062,4072
of|4073,4075
atelectasis|4076,4087
in|4088,4090
<EOL>|4091,4092
the|4092,4095
left|4096,4100
upper|4101,4106
lobe|4107,4111
.|4111,4112
Sternal|4114,4121
wires|4122,4127
are|4128,4131
aligned|4132,4139
.|4139,4140
Widened|4142,4149
<EOL>|4150,4151
mediastinum|4151,4162
has|4163,4166
improved|4167,4175
.|4175,4176
A|4178,4179
small|4180,4185
air|4186,4189
-|4189,4190
fluid|4190,4195
level|4196,4201
in|4202,4204
the|4205,4208
<EOL>|4209,4210
retrosternal|4210,4222
region|4223,4229
suggests|4230,4238
the|4239,4242
presence|4243,4251
of|4252,4254
a|4255,4256
tiny|4257,4261
pneumothorax|4262,4274
<EOL>|4275,4276
and|4276,4279
small|4280,4285
effusion|4286,4294
.|4294,4295
These|4297,4302
are|4303,4306
most|4307,4311
likely|4312,4318
located|4319,4326
in|4327,4329
the|4330,4333
left|4334,4338
<EOL>|4339,4340
side|4340,4344
.|4344,4345
<EOL>|4346,4347
<EOL>|4347,4348
_|4348,4349
_|4349,4350
_|4350,4351
06|4352,4354
:|4354,4355
05AM|4355,4359
BLOOD|4360,4365
WBC|4366,4369
-|4369,4370
11|4370,4372
.|4372,4373
7|4373,4374
*|4374,4375
RBC|4376,4379
-|4379,4380
3|4380,4381
.|4381,4382
06|4382,4384
*|4384,4385
Hgb|4386,4389
-|4389,4390
10|4390,4392
.|4392,4393
4|4393,4394
*|4394,4395
Hct|4396,4399
-|4399,4400
30|4400,4402
.|4402,4403
5|4403,4404
*|4404,4405
<EOL>|4406,4407
MCV|4407,4410
-|4410,4411
100|4411,4414
*|4414,4415
MCH|4416,4419
-|4419,4420
33|4420,4422
.|4422,4423
9|4423,4424
*|4424,4425
MCHC|4426,4430
-|4430,4431
34.0|4431,4435
RDW|4436,4439
-|4439,4440
13.5|4440,4444
Plt|4445,4448
_|4449,4450
_|4450,4451
_|4451,4452
<EOL>|4452,4453
_|4453,4454
_|4454,4455
_|4455,4456
06|4457,4459
:|4459,4460
15AM|4460,4464
BLOOD|4465,4470
WBC|4471,4474
-|4474,4475
11|4475,4477
.|4477,4478
1|4478,4479
*|4479,4480
RBC|4481,4484
-|4484,4485
3|4485,4486
.|4486,4487
23|4487,4489
*|4489,4490
Hgb|4491,4494
-|4494,4495
11|4495,4497
.|4497,4498
1|4498,4499
*|4499,4500
Hct|4501,4504
-|4504,4505
32|4505,4507
.|4507,4508
1|4508,4509
*|4509,4510
<EOL>|4511,4512
MCV|4512,4515
-|4515,4516
99|4516,4518
*|4518,4519
MCH|4520,4523
-|4523,4524
34|4524,4526
.|4526,4527
4|4527,4528
*|4528,4529
MCHC|4530,4534
-|4534,4535
34.6|4535,4539
RDW|4540,4543
-|4543,4544
13.3|4544,4548
Plt|4549,4552
_|4553,4554
_|4554,4555
_|4555,4556
<EOL>|4556,4557
_|4557,4558
_|4558,4559
_|4559,4560
08|4561,4563
:|4563,4564
20AM|4564,4568
BLOOD|4569,4574
WBC|4575,4578
-|4578,4579
14|4579,4581
.|4581,4582
0|4582,4583
*|4583,4584
RBC|4585,4588
-|4588,4589
3|4589,4590
.|4590,4591
26|4591,4593
*|4593,4594
Hgb|4595,4598
-|4598,4599
10|4599,4601
.|4601,4602
8|4602,4603
*|4603,4604
Hct|4605,4608
-|4608,4609
32|4609,4611
.|4611,4612
3|4612,4613
*|4613,4614
<EOL>|4615,4616
MCV|4616,4619
-|4619,4620
99|4620,4622
*|4622,4623
MCH|4624,4627
-|4627,4628
33|4628,4630
.|4630,4631
2|4631,4632
*|4632,4633
MCHC|4634,4638
-|4638,4639
33.4|4639,4643
RDW|4644,4647
-|4647,4648
13.3|4648,4652
Plt|4653,4656
_|4657,4658
_|4658,4659
_|4659,4660
<EOL>|4660,4661
_|4661,4662
_|4662,4663
_|4663,4664
06|4665,4667
:|4667,4668
05AM|4668,4672
BLOOD|4673,4678
Na|4679,4681
-|4681,4682
137|4682,4685
K|4686,4687
-|4687,4688
4.1|4688,4691
Cl|4692,4694
-|4694,4695
97|4695,4697
<EOL>|4697,4698
_|4698,4699
_|4699,4700
_|4700,4701
06|4702,4704
:|4704,4705
15AM|4705,4709
BLOOD|4710,4715
Glucose|4716,4723
-|4723,4724
161|4724,4727
*|4727,4728
UreaN|4729,4734
-|4734,4735
19|4735,4737
Creat|4738,4743
-|4743,4744
1.1|4744,4747
Na|4748,4750
-|4750,4751
136|4751,4754
<EOL>|4755,4756
K|4756,4757
-|4757,4758
4.0|4758,4761
Cl|4762,4764
-|4764,4765
97|4765,4767
HCO3|4768,4772
-|4772,4773
29|4773,4775
AnGap|4776,4781
-|4781,4782
14|4782,4784
<EOL>|4784,4785
_|4785,4786
_|4786,4787
_|4787,4788
08|4789,4791
:|4791,4792
00AM|4792,4796
BLOOD|4797,4802
Glucose|4803,4810
-|4810,4811
230|4811,4814
*|4814,4815
UreaN|4816,4821
-|4821,4822
14|4822,4824
Creat|4825,4830
-|4830,4831
0.9|4831,4834
Na|4835,4837
-|4837,4838
136|4838,4841
<EOL>|4842,4843
K|4843,4844
-|4844,4845
4.1|4845,4848
Cl|4849,4851
-|4851,4852
98|4852,4854
HCO3|4855,4859
-|4859,4860
26|4860,4862
AnGap|4863,4868
-|4868,4869
16|4869,4871
<EOL>|4871,4872
_|4872,4873
_|4873,4874
_|4874,4875
08|4876,4878
:|4878,4879
20AM|4879,4883
BLOOD|4884,4889
Glucose|4890,4897
-|4897,4898
238|4898,4901
*|4901,4902
UreaN|4903,4908
-|4908,4909
16|4909,4911
Creat|4912,4917
-|4917,4918
1.0|4918,4921
Na|4922,4924
-|4924,4925
134|4925,4928
<EOL>|4929,4930
K|4930,4931
-|4931,4932
4.6|4932,4935
Cl|4936,4938
-|4938,4939
100|4939,4942
HCO3|4943,4947
-|4947,4948
22|4948,4950
AnGap|4951,4956
-|4956,4957
17|4957,4959
<EOL>|4959,4960
_|4960,4961
_|4961,4962
_|4962,4963
:|4963,4964
00AM|4964,4968
BLOOD|4969,4974
Glucose|4975,4982
-|4982,4983
98|4983,4985
UreaN|4986,4991
-|4991,4992
13|4992,4994
Creat|4995,5000
-|5000,5001
0.9|5001,5004
Na|5005,5007
-|5007,5008
136|5008,5011
<EOL>|5012,5013
K|5013,5014
-|5014,5015
4.7|5015,5018
Cl|5019,5021
-|5021,5022
106|5022,5025
HCO|5026,5029
_|5029,5030
_|5030,5031
_|5031,5032
AnGap|5033,5038
-|5038,5039
12|5039,5041
<EOL>|5041,5042
<EOL>|5043,5044
The|5067,5070
patient|5071,5078
was|5079,5082
brought|5083,5090
to|5091,5093
the|5094,5097
Operating|5098,5107
Room|5108,5112
on|5113,5115
_|5116,5117
_|5117,5118
_|5118,5119
where|5120,5125
<EOL>|5126,5127
the|5127,5130
patient|5131,5138
underwent|5139,5148
Off|5149,5152
pump|5153,5157
coronary|5158,5166
artery|5167,5173
bypass|5174,5180
graft|5181,5186
x3|5187,5189
,|5189,5190
<EOL>|5191,5192
left|5192,5196
internal|5197,5205
mammary|5206,5213
artery|5214,5220
to|5221,5223
left|5224,5228
anterior|5229,5237
descending|5238,5248
artery|5249,5255
<EOL>|5256,5257
and|5257,5260
saphenous|5261,5270
vein|5271,5275
grafts|5276,5282
to|5283,5285
diagonal|5286,5294
,|5294,5295
and|5296,5299
obtuse|5300,5306
marginal|5307,5315
<EOL>|5315,5316
arteries|5316,5324
.|5324,5325
Endoscopic|5326,5336
harvesting|5337,5347
of|5348,5350
the|5351,5354
long|5355,5359
saphenous|5360,5369
vein|5370,5374
.|5374,5375
<EOL>|5375,5376
Overall|5376,5383
the|5384,5387
patient|5388,5395
tolerated|5396,5405
the|5406,5409
procedure|5410,5419
well|5420,5424
and|5425,5428
<EOL>|5429,5430
post-operatively|5430,5446
was|5447,5450
transferred|5451,5462
to|5463,5465
the|5466,5469
CVICU|5470,5475
in|5476,5478
stable|5479,5485
<EOL>|5486,5487
condition|5487,5496
for|5497,5500
recovery|5501,5509
and|5510,5513
invasive|5514,5522
monitoring|5523,5533
.|5533,5534
She|5535,5538
required|5539,5547
<EOL>|5548,5549
Nitroglycerin|5549,5562
for|5563,5566
hypertension|5567,5579
her|5580,5583
first|5584,5589
night|5590,5595
post|5596,5600
op|5601,5603
but|5604,5607
was|5608,5611
<EOL>|5612,5613
transitioned|5613,5625
to|5626,5628
oral|5629,5633
betablocker|5634,5645
and|5646,5649
diuretics|5650,5659
.|5659,5660
POD|5661,5664
1|5665,5666
found|5667,5672
the|5673,5676
<EOL>|5677,5678
patient|5678,5685
extubated|5686,5695
,|5695,5696
alert|5697,5702
and|5703,5706
oriented|5707,5715
and|5716,5719
breathing|5720,5729
comfortably|5730,5741
.|5741,5742
<EOL>|5743,5744
The|5745,5748
patient|5749,5756
was|5757,5760
neurologically|5761,5775
intact|5776,5782
and|5783,5786
hemodynamically|5787,5802
<EOL>|5803,5804
stable|5804,5810
.|5810,5811
The|5812,5815
patient|5816,5823
was|5824,5827
transferred|5828,5839
to|5840,5842
the|5843,5846
telemetry|5847,5856
floor|5857,5862
for|5863,5866
<EOL>|5867,5868
further|5868,5875
recovery|5876,5884
.|5884,5885
Chest|5886,5891
tubes|5892,5897
and|5898,5901
pacing|5902,5908
wires|5909,5914
were|5915,5919
discontinued|5920,5932
<EOL>|5933,5934
without|5934,5941
complication|5942,5954
.|5954,5955
She|5956,5959
was|5960,5963
started|5964,5971
on|5972,5974
plavix|5975,5981
due|5982,5985
to|5986,5988
being|5989,5994
<EOL>|5995,5996
done|5996,6000
off|6001,6004
pump|6005,6009
and|6010,6013
will|6014,6018
it|6019,6021
need|6022,6026
to|6027,6029
be|6030,6032
continued|6033,6042
for|6043,6046
six|6047,6050
months|6051,6057
.|6057,6058
<EOL>|6059,6060
Blood|6060,6065
sugars|6066,6072
were|6073,6077
closely|6078,6085
monitored|6086,6095
and|6096,6099
she|6100,6103
was|6104,6107
restarted|6108,6117
on|6118,6120
her|6121,6124
<EOL>|6125,6126
home|6126,6130
regime|6131,6137
which|6138,6143
have|6144,6148
slowly|6149,6155
improved|6156,6164
.|6164,6165
The|6166,6169
patient|6170,6177
was|6178,6181
<EOL>|6182,6183
evaluated|6183,6192
by|6193,6195
the|6196,6199
physical|6200,6208
therapy|6209,6216
service|6217,6224
for|6225,6228
assistance|6229,6239
with|6240,6244
<EOL>|6245,6246
strength|6246,6254
and|6255,6258
mobility|6259,6267
.|6267,6268
By|6270,6272
the|6273,6276
time|6277,6281
of|6282,6284
discharge|6285,6294
on|6295,6297
POD|6298,6301
5|6302,6303
the|6304,6307
<EOL>|6308,6309
patient|6309,6316
was|6317,6320
ambulating|6321,6331
freely|6332,6338
,|6338,6339
the|6340,6343
wound|6344,6349
was|6350,6353
healing|6354,6361
and|6362,6365
pain|6366,6370
<EOL>|6371,6372
was|6372,6375
controlled|6376,6386
with|6387,6391
oral|6392,6396
analgesics|6397,6407
.|6407,6408
The|6410,6413
patient|6414,6421
was|6422,6425
discharged|6426,6436
<EOL>|6437,6438
home|6438,6442
with|6443,6447
visiting|6448,6456
nurse|6457,6462
services|6463,6471
in|6472,6474
good|6475,6479
condition|6480,6489
with|6490,6494
<EOL>|6495,6496
appropriate|6496,6507
follow|6508,6514
up|6515,6517
instructions|6518,6530
.|6530,6531
<EOL>|6531,6532
<EOL>|6532,6533
<EOL>|6534,6535
Medications|6535,6546
on|6547,6549
Admission|6550,6559
:|6559,6560
<EOL>|6560,6561
Preadmission|6561,6573
medications|6574,6585
listed|6586,6592
are|6593,6596
correct|6597,6604
and|6605,6608
complete|6609,6617
.|6617,6618
<EOL>|6620,6621
Information|6621,6632
was|6633,6636
obtained|6637,6645
from|6646,6650
webOMR|6651,6657
.|6657,6658
<EOL>|6658,6659
1.|6659,6661
Atorvastatin|6662,6674
40|6675,6677
mg|6678,6680
PO|6681,6683
DAILY|6684,6689
<EOL>|6690,6691
2.|6691,6693
Albuterol|6694,6703
Inhaler|6704,6711
2|6712,6713
PUFF|6714,6718
IH|6719,6721
Q4H|6722,6725
:|6725,6726
PRN|6726,6729
wheezing|6730,6738
<EOL>|6739,6740
3.|6740,6742
Benzonatate|6743,6754
100|6755,6758
mg|6759,6761
PO|6762,6764
TID|6765,6768
:|6768,6769
PRN|6769,6772
tos|6773,6776
<EOL>|6777,6778
4.|6778,6780
Clopidogrel|6781,6792
75|6793,6795
mg|6796,6798
PO|6799,6801
DAILY|6802,6807
<EOL>|6808,6809
5.|6809,6811
Fluticasone|6812,6823
Propionate|6824,6834
110mcg|6835,6841
2|6842,6843
PUFF|6844,6848
IH|6849,6851
BID|6852,6855
<EOL>|6856,6857
6.|6857,6859
Glargine|6860,6868
80|6869,6871
Units|6872,6877
Bedtime|6878,6885
<EOL>|6885,6886
Insulin|6886,6893
SC|6894,6896
Sliding|6897,6904
Scale|6905,6910
using|6911,6916
HUM|6917,6920
Insulin|6921,6928
<EOL>|6928,6929
7.|6929,6931
Isosorbide|6932,6942
Mononitrate|6943,6954
(|6955,6956
Extended|6956,6964
Release|6965,6972
)|6972,6973
60|6974,6976
mg|6977,6979
PO|6980,6982
DAILY|6983,6988
<EOL>|6989,6990
8.|6990,6992
Metoprolol|6993,7003
Succinate|7004,7013
XL|7014,7016
100|7017,7020
mg|7021,7023
PO|7024,7026
DAILY|7027,7032
<EOL>|7033,7034
9.|7034,7036
Metronidazole|7037,7050
Gel|7051,7054
0.75|7055,7059
%|7059,7060
-|7060,7061
Vaginal|7061,7068
1|7069,7070
Appl|7071,7075
VG|7076,7078
HS|7079,7081
<EOL>|7082,7083
10.|7083,7086
Naproxen|7087,7095
500|7096,7099
mg|7100,7102
PO|7103,7105
Q8H|7106,7109
:|7109,7110
PRN|7110,7113
pain|7114,7118
<EOL>|7119,7120
11|7120,7122
.|7122,7123
Nitroglycerin|7124,7137
SL|7138,7140
0.4|7141,7144
mg|7145,7147
SL|7148,7150
PRN|7151,7154
cp|7155,7157
<EOL>|7158,7159
12.|7159,7162
Oxycodone|7163,7172
-|7172,7173
Acetaminophen|7173,7186
(|7187,7188
5mg|7188,7191
-|7191,7192
325mg|7192,7197
)|7197,7198
1|7199,7200
TAB|7201,7204
PO|7205,7207
Q6H|7208,7211
:|7211,7212
PRN|7212,7215
pain|7216,7220
<EOL>|7221,7222
13|7222,7224
.|7224,7225
Pantoprazole|7226,7238
40|7239,7241
mg|7242,7244
PO|7245,7247
Q12H|7248,7252
<EOL>|7253,7254
14.|7254,7257
Ropinirole|7258,7268
0.25|7269,7273
mg|7274,7276
PO|7277,7279
QPM|7280,7283
<EOL>|7284,7285
15.|7285,7288
Valsartan|7289,7298
80|7299,7301
mg|7302,7304
PO|7305,7307
DAILY|7308,7313
<EOL>|7314,7315
16|7315,7317
.|7317,7318
Aspirin|7319,7326
325|7327,7330
mg|7331,7333
PO|7334,7336
DAILY|7337,7342
<EOL>|7343,7344
17.|7344,7347
Vitamin|7348,7355
D|7356,7357
400|7358,7361
UNIT|7362,7366
PO|7367,7369
DAILY|7370,7375
<EOL>|7376,7377
<EOL>|7377,7378
<EOL>|7379,7380
Discharge|7380,7389
Medications|7390,7401
:|7401,7402
<EOL>|7402,7403
1.|7403,7405
Aspirin|7406,7413
EC|7414,7416
81|7417,7419
mg|7420,7422
PO|7423,7425
DAILY|7426,7431
<EOL>|7432,7433
2.|7433,7435
Atorvastatin|7436,7448
40|7449,7451
mg|7452,7454
PO|7455,7457
DAILY|7458,7463
<EOL>|7464,7465
RX|7465,7467
*|7468,7469
atorvastatin|7469,7481
40|7482,7484
mg|7485,7487
1|7488,7489
tablet|7490,7496
(|7496,7497
s|7497,7498
)|7498,7499
by|7500,7502
mouth|7503,7508
daily|7509,7514
Disp|7515,7519
#|7520,7521
*|7521,7522
30|7522,7524
<EOL>|7525,7526
Tablet|7526,7532
Refills|7533,7540
:|7540,7541
*|7541,7542
0|7542,7543
<EOL>|7543,7544
3.|7544,7546
Clopidogrel|7547,7558
75|7559,7561
mg|7562,7564
PO|7565,7567
DAILY|7568,7573
<EOL>|7574,7575
RX|7575,7577
*|7578,7579
clopidogrel|7579,7590
75|7591,7593
mg|7594,7596
1|7597,7598
tablet|7599,7605
(|7605,7606
s|7606,7607
)|7607,7608
by|7609,7611
mouth|7612,7617
daily|7618,7623
Disp|7624,7628
#|7629,7630
*|7630,7631
90|7631,7633
<EOL>|7634,7635
Tablet|7635,7641
Refills|7642,7649
:|7649,7650
*|7650,7651
1|7651,7652
<EOL>|7652,7653
4.|7653,7655
Fluticasone|7656,7667
Propionate|7668,7678
110mcg|7679,7685
2|7686,7687
PUFF|7688,7692
IH|7693,7695
BID|7696,7699
<EOL>|7700,7701
RX|7701,7703
*|7704,7705
fluticasone|7705,7716
[|7717,7718
Flovent|7718,7725
HFA|7726,7729
]|7729,7730
220|7731,7734
mcg|7735,7738
2|7739,7740
puffs|7741,7746
twice|7747,7752
a|7753,7754
day|7755,7758
Disp|7759,7763
<EOL>|7764,7765
#|7765,7766
*|7766,7767
1|7767,7768
Inhaler|7769,7776
Refills|7777,7784
:|7784,7785
*|7785,7786
0|7786,7787
<EOL>|7787,7788
5.|7788,7790
Glargine|7791,7799
50|7800,7802
Units|7803,7808
Bedtime|7809,7816
<EOL>|7816,7817
Insulin|7817,7824
SC|7825,7827
Sliding|7828,7835
Scale|7836,7841
using|7842,7847
HUM|7848,7851
Insulin|7852,7859
<EOL>|7859,7860
6.|7860,7862
Oxycodone|7863,7872
-|7872,7873
Acetaminophen|7873,7886
(|7887,7888
5mg|7888,7891
-|7891,7892
325mg|7892,7897
)|7897,7898
1|7899,7900
TAB|7901,7904
PO|7905,7907
Q6H|7908,7911
:|7911,7912
PRN|7912,7915
pain|7916,7920
<EOL>|7921,7922
RX|7922,7924
*|7925,7926
oxycodone|7926,7935
-|7935,7936
acetaminophen|7936,7949
5|7950,7951
mg|7952,7954
-|7954,7955
325|7955,7958
mg|7959,7961
1|7962,7963
tablet|7964,7970
(|7970,7971
s|7971,7972
)|7972,7973
by|7974,7976
mouth|7977,7982
Q|7983,7984
4|7985,7986
<EOL>|7987,7988
hrs|7988,7991
Disp|7992,7996
#|7997,7998
*|7998,7999
30|7999,8001
Tablet|8002,8008
Refills|8009,8016
:|8016,8017
*|8017,8018
0|8018,8019
<EOL>|8019,8020
7.|8020,8022
Pantoprazole|8023,8035
40|8036,8038
mg|8039,8041
PO|8042,8044
Q24H|8045,8049
<EOL>|8050,8051
RX|8051,8053
*|8054,8055
pantoprazole|8055,8067
40|8068,8070
mg|8071,8073
1|8074,8075
tablet|8076,8082
(|8082,8083
s|8083,8084
)|8084,8085
by|8086,8088
mouth|8089,8094
daily|8095,8100
Disp|8101,8105
#|8106,8107
*|8107,8108
30|8108,8110
<EOL>|8111,8112
Tablet|8112,8118
Refills|8119,8126
:|8126,8127
*|8127,8128
0|8128,8129
<EOL>|8129,8130
8.|8130,8132
Ropinirole|8133,8143
0.25|8144,8148
mg|8149,8151
PO|8152,8154
QPM|8155,8158
<EOL>|8159,8160
9.|8160,8162
Furosemide|8163,8173
40|8174,8176
mg|8177,8179
PO|8180,8182
DAILY|8183,8188
Duration|8189,8197
:|8197,8198
7|8199,8200
Days|8201,8205
<EOL>|8206,8207
RX|8207,8209
*|8210,8211
furosemide|8211,8221
[|8222,8223
Lasix|8223,8228
]|8228,8229
40|8230,8232
mg|8233,8235
1|8236,8237
tablet|8238,8244
(|8244,8245
s|8245,8246
)|8246,8247
by|8248,8250
mouth|8251,8256
daily|8257,8262
Disp|8263,8267
#|8268,8269
*|8269,8270
7|8270,8271
<EOL>|8272,8273
Tablet|8273,8279
Refills|8280,8287
:|8287,8288
*|8288,8289
0|8289,8290
<EOL>|8290,8291
10.|8291,8294
Ibuprofen|8295,8304
600|8305,8308
mg|8309,8311
PO|8312,8314
Q6H|8315,8318
:|8318,8319
PRN|8319,8322
pain|8323,8327
<EOL>|8328,8329
take|8329,8333
with|8334,8338
food|8339,8343
<EOL>|8344,8345
RX|8345,8347
*|8348,8349
ibuprofen|8349,8358
600|8359,8362
mg|8363,8365
1|8366,8367
tablet|8368,8374
(|8374,8375
s|8375,8376
)|8376,8377
by|8378,8380
mouth|8381,8386
three|8387,8392
times|8393,8398
a|8399,8400
day|8401,8404
Disp|8405,8409
<EOL>|8410,8411
#|8411,8412
*|8412,8413
90|8413,8415
Tablet|8416,8422
Refills|8423,8430
:|8430,8431
*|8431,8432
0|8432,8433
<EOL>|8433,8434
11.|8434,8437
Metoprolol|8438,8448
Tartrate|8449,8457
25|8458,8460
mg|8461,8463
PO|8464,8466
TID|8467,8470
<EOL>|8471,8472
Hold|8472,8476
for|8477,8480
HR|8481,8483
<|8484,8485
55|8486,8488
or|8489,8491
SBP|8492,8495
<|8496,8497
90|8498,8500
and|8501,8504
call|8505,8509
medical|8510,8517
provider|8518,8526
.|8526,8527
<EOL>|8528,8529
RX|8529,8531
*|8532,8533
metoprolol|8533,8543
tartrate|8544,8552
25|8553,8555
mg|8556,8558
1|8559,8560
tablet|8561,8567
(|8567,8568
s|8568,8569
)|8569,8570
by|8571,8573
mouth|8574,8579
three|8580,8585
times|8586,8591
a|8592,8593
<EOL>|8594,8595
day|8595,8598
Disp|8599,8603
#|8604,8605
*|8605,8606
90|8606,8608
Tablet|8609,8615
Refills|8616,8623
:|8623,8624
*|8624,8625
1|8625,8626
<EOL>|8626,8627
12.|8627,8630
Potassium|8631,8640
Chloride|8641,8649
20|8650,8652
mEq|8653,8656
PO|8657,8659
DAILY|8660,8665
<EOL>|8666,8667
RX|8667,8669
*|8670,8671
potassium|8671,8680
chloride|8681,8689
20|8690,8692
mEq|8693,8696
1|8697,8698
tablet|8699,8705
by|8706,8708
mouth|8709,8714
daily|8715,8720
Disp|8721,8725
#|8726,8727
*|8727,8728
7|8728,8729
<EOL>|8730,8731
Tablet|8731,8737
Refills|8738,8745
:|8745,8746
*|8746,8747
0|8747,8748
<EOL>|8748,8749
13.|8749,8752
Albuterol|8753,8762
Inhaler|8763,8770
2|8771,8772
PUFF|8773,8777
IH|8778,8780
Q4H|8781,8784
:|8784,8785
PRN|8785,8788
wheezing|8789,8797
<EOL>|8798,8799
RX|8799,8801
*|8802,8803
albuterol|8803,8812
2|8814,8815
puffs|8816,8821
PRN|8822,8825
Q|8826,8827
4|8828,8829
hrs|8830,8833
Disp|8834,8838
#|8839,8840
*|8840,8841
1|8841,8842
Inhaler|8843,8850
Refills|8851,8858
:|8858,8859
*|8859,8860
0|8860,8861
<EOL>|8861,8862
14.|8862,8865
Vitamin|8866,8873
D|8874,8875
400|8876,8879
UNIT|8880,8884
PO|8885,8887
DAILY|8888,8893
<EOL>|8894,8895
<EOL>|8895,8896
<EOL>|8897,8898
Discharge|8898,8907
Disposition|8908,8919
:|8919,8920
<EOL>|8920,8921
Home|8921,8925
With|8926,8930
Service|8931,8938
<EOL>|8938,8939
<EOL>|8940,8941
Facility|8941,8949
:|8949,8950
<EOL>|8950,8951
_|8951,8952
_|8952,8953
_|8953,8954
<EOL>|8954,8955
<EOL>|8956,8957
_|8957,8958
_|8958,8959
_|8959,8960
Diagnosis|8961,8970
:|8970,8971
<EOL>|8971,8972
Coronary|8972,8980
artery|8981,8987
disease|8988,8995
(|8995,8996
s|8996,8997
/|8997,8998
p|8998,8999
MI|9000,9002
_|9003,9004
_|9004,9005
_|9005,9006
,|9006,9007
BMS|9008,9011
to|9012,9014
proximal|9015,9023
LAD|9024,9027
_|9028,9029
_|9029,9030
_|9030,9031
,|9031,9032
<EOL>|9033,9034
DES|9034,9037
to|9038,9040
mid|9041,9044
LAD|9045,9048
_|9049,9050
_|9050,9051
_|9051,9052
,|9052,9053
DES|9054,9057
to|9058,9060
edge|9061,9065
ISR|9066,9069
of|9070,9072
mid|9073,9076
LAD|9077,9080
DES|9081,9084
and|9085,9088
stenosis|9089,9097
<EOL>|9098,9099
distal|9099,9105
to|9106,9108
stent|9109,9114
_|9115,9116
_|9116,9117
_|9117,9118
,|9118,9119
DES|9120,9123
to|9124,9126
OM1|9127,9130
,|9130,9131
_|9132,9133
_|9133,9134
_|9134,9135
.|9135,9136
<EOL>|9137,9138
diastolic|9138,9147
congestive|9148,9158
heart|9159,9164
failure|9165,9172
<EOL>|9172,9173
Hypertension|9173,9185
<EOL>|9185,9186
Dyslipidemia|9186,9198
<EOL>|9198,9199
Morbid|9199,9205
obesity|9206,9213
<EOL>|9213,9214
COPD|9214,9218
<EOL>|9218,9219
GERD|9219,9223
<EOL>|9223,9224
Rt|9224,9226
rotator|9227,9234
cuff|9235,9239
injury|9240,9246
/|9246,9247
bursitis|9247,9255
(|9255,9256
outpt|9256,9261
_|9262,9263
_|9263,9264
_|9264,9265
,|9265,9266
<EOL>|9267,9268
Migraines|9268,9277
,|9277,9278
<EOL>|9279,9280
Depression|9280,9290
/|9290,9291
Anxiety|9291,9298
<EOL>|9298,9299
DJD|9299,9302
<EOL>|9302,9303
Hemorrhoids|9303,9314
<EOL>|9315,9316
Rosacea|9316,9323
<EOL>|9324,9325
Left|9325,9329
foot|9330,9334
tendion|9335,9342
repair|9343,9349
<EOL>|9349,9350
<EOL>|9350,9351
<EOL>|9352,9353
Alert|9374,9379
and|9380,9383
oriented|9384,9392
x3|9393,9395
nonfocal|9396,9404
<EOL>|9404,9405
Ambulating|9405,9415
,|9415,9416
gait|9417,9421
steady|9422,9428
<EOL>|9428,9429
Sternal|9429,9436
pain|9437,9441
managed|9442,9449
with|9450,9454
oral|9455,9459
analgesics|9460,9470
<EOL>|9470,9471
Sternal|9471,9478
Incision|9479,9487
-|9488,9489
healing|9490,9497
well|9498,9502
,|9502,9503
no|9504,9506
erythema|9507,9515
or|9516,9518
drainage|9519,9527
<EOL>|9527,9528
<EOL>|9529,9530
<EOL>|9530,9531
<EOL>|9532,9533
Please|9557,9563
shower|9564,9570
daily|9571,9576
including|9577,9586
washing|9587,9594
incisions|9595,9604
gently|9605,9611
with|9612,9616
mild|9617,9621
<EOL>|9622,9623
soap|9623,9627
,|9627,9628
no|9629,9631
baths|9632,9637
or|9638,9640
swimming|9641,9649
,|9649,9650
and|9651,9654
look|9655,9659
at|9660,9662
your|9663,9667
incisions|9668,9677
<EOL>|9677,9678
Please|9678,9684
NO|9685,9687
lotions|9688,9695
,|9695,9696
cream|9697,9702
,|9702,9703
powder|9704,9710
,|9710,9711
or|9712,9714
ointments|9715,9724
to|9725,9727
incisions|9728,9737
<EOL>|9737,9738
Each|9738,9742
morning|9743,9750
you|9751,9754
should|9755,9761
weigh|9762,9767
yourself|9768,9776
and|9777,9780
then|9781,9785
in|9786,9788
the|9789,9792
evening|9793,9800
<EOL>|9801,9802
take|9802,9806
your|9807,9811
temperature|9812,9823
,|9823,9824
these|9825,9830
should|9831,9837
be|9838,9840
written|9841,9848
down|9849,9853
on|9854,9856
the|9857,9860
chart|9861,9866
<EOL>|9866,9867
No|9867,9869
driving|9870,9877
for|9878,9881
approximately|9882,9895
one|9896,9899
month|9900,9905
and|9906,9909
while|9910,9915
taking|9916,9922
<EOL>|9923,9924
narcotics|9924,9933
,|9933,9934
will|9935,9939
be|9940,9942
discussed|9943,9952
at|9953,9955
follow|9956,9962
up|9963,9965
appointment|9966,9977
with|9978,9982
<EOL>|9983,9984
surgeon|9984,9991
when|9992,9996
you|9997,10000
will|10001,10005
be|10006,10008
able|10009,10013
to|10014,10016
drive|10017,10022
<EOL>|10022,10023
No|10023,10025
lifting|10026,10033
more|10034,10038
than|10039,10043
10|10044,10046
pounds|10047,10053
for|10054,10057
10|10058,10060
weeks|10061,10066
<EOL>|10066,10067
<EOL>|10067,10068
*|10068,10069
*|10069,10070
Please|10070,10076
call|10077,10081
cardiac|10082,10089
surgery|10090,10097
office|10098,10104
with|10105,10109
any|10110,10113
questions|10114,10123
or|10124,10126
<EOL>|10127,10128
concerns|10128,10136
_|10137,10138
_|10138,10139
_|10139,10140
.|10140,10141
Answering|10142,10151
service|10152,10159
will|10160,10164
contact|10165,10172
on|10173,10175
call|10176,10180
<EOL>|10181,10182
person|10182,10188
during|10189,10195
off|10196,10199
hours|10200,10205
*|10205,10206
*|10206,10207
<EOL>|10207,10208
Females|10208,10215
:|10215,10216
Please|10217,10223
wear|10224,10228
bra|10229,10232
to|10233,10235
reduce|10236,10242
pulling|10243,10250
on|10251,10253
incision|10254,10262
,|10262,10263
avoid|10264,10269
<EOL>|10270,10271
rubbing|10271,10278
on|10279,10281
lower|10282,10287
edge|10288,10292
<EOL>|10292,10293
<EOL>|10293,10294
<EOL>|10295,10296
Followup|10296,10304
Instructions|10305,10317
:|10317,10318
<EOL>|10318,10319
_|10319,10320
_|10320,10321
_|10321,10322
<EOL>|10322,10323

