 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|27,28
_|28,29
_|29,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
ORTHOPAEDICS|153,165
<EOL>|165,166
<EOL>|167,168
Allergies|168,177
:|177,178
<EOL>|179,180
meropenem|180,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Chief|210,215
Complaint|216,225
:|225,226
<EOL>|226,227
left|227,231
hip|232,235
pain|236,240
<EOL>|240,241
<EOL>|242,243
Major|243,248
Surgical|249,257
or|258,260
Invasive|261,269
Procedure|270,279
:|279,280
<EOL>|280,281
Closed|281,287
reduction|288,297
and|298,301
percutaneous|302,314
pinning|315,322
,|322,323
left|324,328
<EOL>|328,329
femoral|329,336
neck|337,341
fracture|342,350
<EOL>|350,351
<EOL>|351,352
<EOL>|353,354
History|354,361
of|362,364
Present|365,372
Illness|373,380
:|380,381
<EOL>|381,382
This|382,386
is|387,389
a|390,391
_|392,393
_|393,394
_|394,395
yo|396,398
woman|399,404
in|405,407
her|408,411
USOH|412,416
until|417,422
the|423,426
day|427,430
of|431,433
presentation|434,446
<EOL>|447,448
when|448,452
she|453,456
sustained|457,466
a|467,468
mechanical|469,479
fall|480,484
onto|485,489
her|490,493
left|494,498
lower|499,504
<EOL>|505,506
extremity|506,515
with|516,520
immediate|521,530
pain|531,535
,|535,536
inability|537,546
to|547,549
ambulate|550,558
.|558,559
The|561,564
<EOL>|565,566
patient|566,573
denies|574,580
LOC|581,584
,|584,585
premonitory|586,597
symptoms|598,606
and|607,610
ROS|611,614
is|615,617
otherwise|618,627
at|628,630
<EOL>|631,632
baseline|632,640
.|640,641
<EOL>|642,643
<EOL>|643,644
<EOL>|645,646
Past|646,650
Medical|651,658
History|659,666
:|666,667
<EOL>|667,668
Anemia|668,674
<EOL>|676,677
Borderline|677,687
cholesterol|688,699
<EOL>|701,702
Recurrent|702,711
C.|712,714
Diff|715,719
<EOL>|721,722
Flatulence|722,732
<EOL>|734,735
Heart|735,740
Murmur|741,747
<EOL>|749,750
Hypertension|750,762
<EOL>|764,765
Hypothyroidism|765,779
<EOL>|781,782
Mitral|782,788
Regurgitation|789,802
<EOL>|804,805
Osteoporosis|805,817
<EOL>|819,820
Pneumonia|820,829
<EOL>|831,832
Sinusitis|832,841
<EOL>|843,844
Sjo|844,847
_|847,848
_|848,849
_|849,850
<EOL>|852,853
<EOL>|854,855
Social|855,861
History|862,869
:|869,870
<EOL>|870,871
_|871,872
_|872,873
_|873,874
<EOL>|874,875
Family|875,881
History|882,889
:|889,890
<EOL>|890,891
Long|891,895
history|896,903
of|904,906
hypertension|907,919
in|920,922
her|923,926
family|927,933
.|933,934
Father|936,942
's|942,944
family|945,951
has|952,955
<EOL>|956,957
a|957,958
history|959,966
of|967,969
multiple|970,978
cancers|979,986
.|986,987
She|989,992
has|993,996
a|997,998
grandfather|999,1010
with|1011,1015
a|1016,1017
<EOL>|1018,1019
history|1019,1026
of|1027,1029
stomach|1030,1037
cancer|1038,1044
and|1045,1048
an|1049,1051
uncle|1052,1057
with|1058,1062
a|1063,1064
history|1065,1072
of|1073,1075
throat|1076,1082
<EOL>|1083,1084
cancer|1084,1090
.|1090,1091
No|1093,1095
history|1096,1103
of|1104,1106
colon|1107,1112
cancers|1113,1120
.|1120,1121
Father|1122,1128
had|1129,1132
stroke|1133,1139
.|1139,1140
No|1141,1143
<EOL>|1144,1145
family|1145,1151
h|1152,1153
/|1153,1154
o|1154,1155
MI|1156,1158
.|1158,1159
Mother|1160,1166
had|1167,1170
a|1171,1172
heart|1173,1178
valve|1179,1184
replaced|1185,1193
.|1193,1194
<EOL>|1194,1195
<EOL>|1195,1196
<EOL>|1197,1198
Physical|1198,1206
Exam|1207,1211
:|1211,1212
<EOL>|1212,1213
On|1213,1215
admission|1216,1225
:|1225,1226
<EOL>|1227,1228
Pelvis|1228,1234
stable|1235,1241
to|1242,1244
AP|1245,1247
and|1248,1251
lateral|1252,1259
compression|1260,1271
.|1271,1272
<EOL>|1274,1275
BLE|1275,1278
skin|1279,1283
clean|1284,1289
and|1290,1293
intact|1294,1300
<EOL>|1301,1302
LLE|1302,1305
<EOL>|1305,1306
Shortened|1306,1315
and|1316,1319
externally|1320,1330
rotated|1331,1338
,|1338,1339
painful|1340,1347
with|1348,1352
internal|1353,1361
or|1362,1364
<EOL>|1365,1366
external|1366,1374
rotation|1375,1383
of|1384,1386
the|1387,1390
hip|1391,1394
.|1394,1395
<EOL>|1397,1398
Thighs|1398,1404
and|1405,1408
leg|1409,1412
compartments|1413,1425
soft|1426,1430
<EOL>|1431,1432
Saphenous|1432,1441
,|1441,1442
Sural|1443,1448
,|1448,1449
Deep|1450,1454
peroneal|1455,1463
,|1463,1464
Superficial|1465,1476
peroneal|1477,1485
SILT|1486,1490
<EOL>|1491,1492
_|1492,1493
_|1493,1494
_|1494,1495
FHS|1496,1499
_|1500,1501
_|1501,1502
_|1502,1503
TA|1504,1506
Peroneals|1507,1516
Fire|1517,1521
<EOL>|1522,1523
1|1523,1524
+|1524,1525
_|1526,1527
_|1527,1528
_|1528,1529
and|1530,1533
DP|1534,1536
pulses|1537,1543
<EOL>|1544,1545
Knee|1545,1549
stable|1550,1556
to|1557,1559
varus|1560,1565
and|1566,1569
valgus|1570,1576
stress|1577,1583
.|1583,1584
<EOL>|1587,1588
Negative|1588,1596
anterior|1597,1605
,|1605,1606
posterior|1607,1616
drawer|1617,1623
signs|1624,1629
.|1629,1630
<EOL>|1632,1633
<EOL>|1633,1634
On|1634,1636
discharge|1637,1646
:|1646,1647
<EOL>|1648,1649
NAD|1649,1652
,|1652,1653
A|1654,1655
+|1655,1656
Ox3|1656,1659
<EOL>|1659,1660
INcision|1660,1668
:|1668,1669
dressing|1670,1678
changed|1679,1686
_|1687,1688
_|1688,1689
_|1689,1690
-|1691,1692
c|1693,1694
/|1694,1695
d|1695,1696
/|1696,1697
i|1697,1698
<EOL>|1698,1699
Neurovascularly|1699,1714
intact|1715,1721
,|1721,1722
strenght|1723,1731
intact|1732,1738
,|1738,1739
SILT|1740,1744
s|1745,1746
/|1746,1747
s|1747,1748
/|1748,1749
dp|1749,1751
/|1751,1752
sp|1752,1754
/|1754,1755
t|1755,1756
<EOL>|1757,1758
distributions|1758,1771
<EOL>|1771,1772
WWP|1772,1775
,|1775,1776
2|1777,1778
+|1778,1779
DP|1780,1782
pulse|1783,1788
<EOL>|1788,1789
<EOL>|1789,1790
<EOL>|1791,1792
Pertinent|1792,1801
Results|1802,1809
:|1809,1810
<EOL>|1810,1811
Hip|1811,1814
XR|1815,1817
_|1818,1819
_|1819,1820
_|1820,1821
:|1821,1822
IMPRESSION|1823,1833
:|1833,1834
Impacted|1836,1844
left|1845,1849
subcapital|1850,1860
femoral|1861,1868
neck|1869,1873
<EOL>|1874,1875
fracture|1875,1883
.|1883,1884
<EOL>|1884,1885
<EOL>|1886,1887
Brief|1887,1892
Hospital|1893,1901
Course|1902,1908
:|1908,1909
<EOL>|1909,1910
On|1910,1912
_|1913,1914
_|1914,1915
_|1915,1916
the|1917,1920
pt|1921,1923
was|1924,1927
admitted|1928,1936
to|1937,1939
the|1940,1943
ortho|1944,1949
trauma|1950,1956
service|1957,1964
and|1965,1968
<EOL>|1969,1970
found|1970,1975
to|1976,1978
have|1979,1983
a|1984,1985
valgus|1986,1992
impacted|1993,2001
left|2002,2006
femoral|2007,2014
neck|2015,2019
hip|2020,2023
fracture|2024,2032
,|2032,2033
<EOL>|2034,2035
for|2035,2038
which|2039,2044
she|2045,2048
underwent|2049,2058
closed|2059,2065
reduction|2066,2075
and|2076,2079
percutaneous|2080,2092
<EOL>|2093,2094
pinning|2094,2101
,|2101,2102
left|2103,2107
<EOL>|2107,2108
femoral|2108,2115
neck|2116,2120
fracture|2121,2129
by|2130,2132
Dr.|2133,2136
_|2137,2138
_|2138,2139
_|2139,2140
<EOL>|2140,2141
<EOL>|2141,2142
On|2142,2144
_|2145,2146
_|2146,2147
_|2147,2148
the|2149,2152
patient|2153,2160
was|2161,2164
noted|2165,2170
to|2171,2173
be|2174,2176
recovering|2177,2187
well|2188,2192
from|2193,2197
<EOL>|2198,2199
surgery|2199,2206
.|2206,2207
She|2208,2211
became|2212,2218
hypotensive|2219,2230
with|2231,2235
physical|2236,2244
therapy|2245,2252
,|2252,2253
which|2254,2259
<EOL>|2260,2261
normalized|2261,2271
after|2272,2277
stopping|2278,2286
exercise|2287,2295
.|2295,2296
<EOL>|2297,2298
<EOL>|2298,2299
On|2299,2301
_|2302,2303
_|2303,2304
_|2304,2305
the|2306,2309
patient|2310,2317
continued|2318,2327
to|2328,2330
do|2331,2333
well|2334,2338
.|2338,2339
She|2340,2343
was|2344,2347
seen|2348,2352
by|2353,2355
<EOL>|2356,2357
physical|2357,2365
therapy|2366,2373
and|2374,2377
cleared|2378,2385
for|2386,2389
discharge|2390,2399
to|2400,2402
a|2403,2404
rehab|2405,2410
facility|2411,2419
.|2419,2420
<EOL>|2421,2422
SOcial|2422,2428
work|2429,2433
saw|2434,2437
pt|2438,2440
for|2441,2444
her|2445,2448
difficulty|2449,2459
coping|2460,2466
with|2467,2471
decreased|2472,2481
<EOL>|2482,2483
mobility|2483,2491
.|2491,2492
Her|2493,2496
labs|2497,2501
showed|2502,2508
sodium|2509,2515
level|2516,2521
of|2522,2524
130|2525,2528
,|2528,2529
unchanged|2530,2539
from|2540,2544
<EOL>|2545,2546
_|2546,2547
_|2547,2548
_|2548,2549
and|2550,2553
similar|2554,2561
to|2562,2564
132|2565,2568
on|2569,2571
admission|2572,2581
.|2581,2582
She|2583,2586
was|2587,2590
given|2591,2596
instructions|2597,2609
<EOL>|2610,2611
to|2611,2613
f|2614,2615
/|2615,2616
u|2616,2617
with|2618,2622
Dr.|2623,2626
_|2627,2628
_|2628,2629
_|2629,2630
in|2631,2633
clinic|2634,2640
in|2641,2643
2|2644,2645
weeks|2646,2651
,|2651,2652
and|2653,2656
will|2657,2661
be|2662,2664
on|2665,2667
<EOL>|2668,2669
lovenox|2669,2676
subq|2677,2681
40|2682,2684
mg|2685,2687
daily|2688,2693
in|2694,2696
the|2697,2700
interim|2701,2708
.|2708,2709
<EOL>|2710,2711
<EOL>|2711,2712
<EOL>|2713,2714
Medications|2714,2725
on|2726,2728
Admission|2729,2738
:|2738,2739
<EOL>|2739,2740
The|2740,2743
Preadmission|2744,2756
Medication|2757,2767
list|2768,2772
is|2773,2775
accurate|2776,2784
and|2785,2788
complete|2789,2797
.|2797,2798
<EOL>|2798,2799
1.|2799,2801
Levothyroxine|2802,2815
Sodium|2816,2822
75|2823,2825
mcg|2826,2829
PO|2830,2832
DAILY|2833,2838
<EOL>|2839,2840
2.|2840,2842
Lisinopril|2843,2853
5|2854,2855
mg|2856,2858
PO|2859,2861
DAILY|2862,2867
<EOL>|2868,2869
3.|2869,2871
MethylPHENIDATE|2872,2887
(|2888,2889
Ritalin|2889,2896
)|2896,2897
2.5|2898,2901
mg|2902,2904
PO|2905,2907
BID|2908,2911
<EOL>|2912,2913
4.|2913,2915
mirtazapine|2916,2927
30|2928,2930
mg|2931,2933
Oral|2934,2938
QHS|2939,2942
<EOL>|2943,2944
<EOL>|2944,2945
<EOL>|2946,2947
Discharge|2947,2956
Medications|2957,2968
:|2968,2969
<EOL>|2969,2970
1.|2970,2972
Levothyroxine|2973,2986
Sodium|2987,2993
75|2994,2996
mcg|2997,3000
PO|3001,3003
DAILY|3004,3009
<EOL>|3010,3011
2.|3011,3013
Lisinopril|3014,3024
5|3025,3026
mg|3027,3029
PO|3030,3032
DAILY|3033,3038
<EOL>|3039,3040
3.|3040,3042
MethylPHENIDATE|3043,3058
(|3059,3060
Ritalin|3060,3067
)|3067,3068
2.5|3069,3072
mg|3073,3075
PO|3076,3078
BID|3079,3082
<EOL>|3083,3084
4.|3084,3086
mirtazapine|3087,3098
30|3099,3101
mg|3102,3104
Oral|3105,3109
QHS|3110,3113
<EOL>|3114,3115
5.|3115,3117
Acetaminophen|3118,3131
1000|3132,3136
mg|3137,3139
PO|3140,3142
TID|3143,3146
<EOL>|3147,3148
6.|3148,3150
Aluminum|3151,3159
-|3159,3160
Magnesium|3160,3169
Hydrox|3170,3176
.|3176,3177
-|3177,3178
Simethicone|3178,3189
_|3190,3191
_|3191,3192
_|3192,3193
ml|3194,3196
PO|3197,3199
QID|3200,3203
:|3203,3204
PRN|3204,3207
<EOL>|3208,3209
Dyspepsia|3209,3218
<EOL>|3219,3220
7.|3220,3222
Artificial|3223,3233
Tears|3234,3239
_|3240,3241
_|3241,3242
_|3242,3243
DROP|3244,3248
BOTH|3249,3253
EYES|3254,3258
PRN|3259,3262
dry|3263,3266
eyes|3267,3271
<EOL>|3272,3273
8.|3273,3275
Biotene|3276,3283
Dry|3284,3287
Mouth|3288,3293
Rinse|3294,3299
(|3300,3301
saliva|3301,3307
substitution|3308,3320
combo|3321,3326
no|3327,3329
.8|3329,3331
)|3331,3332
1|3333,3334
<EOL>|3335,3336
application|3336,3347
Mucous|3348,3354
Membrane|3355,3363
q2hr|3364,3368
<EOL>|3369,3370
9.|3370,3372
Bisacodyl|3373,3382
10|3383,3385
mg|3386,3388
PO|3389,3391
/|3391,3392
PR|3392,3394
DAILY|3395,3400
:|3400,3401
PRN|3401,3404
Constipation|3405,3417
<EOL>|3418,3419
10|3419,3421
.|3421,3422
Calcium|3423,3430
Carbonate|3431,3440
1250|3441,3445
mg|3446,3448
PO|3449,3451
TID|3452,3455
<EOL>|3456,3457
11.|3457,3460
Docusate|3461,3469
Sodium|3470,3476
100|3477,3480
mg|3481,3483
PO|3484,3486
BID|3487,3490
<EOL>|3491,3492
12.|3492,3495
Enoxaparin|3496,3506
Sodium|3507,3513
40|3514,3516
mg|3517,3519
SC|3520,3522
DAILY|3523,3528
DVT|3529,3532
prophylaxis|3533,3544
Duration|3545,3553
:|3553,3554
<EOL>|3555,3556
14|3556,3558
Days|3559,3563
Start|3564,3569
:|3569,3570
_|3571,3572
_|3572,3573
_|3573,3574
,|3574,3575
First|3576,3581
Dose|3582,3586
:|3586,3587
Next|3588,3592
Routine|3593,3600
Administration|3601,3615
<EOL>|3616,3617
Time|3617,3621
<EOL>|3622,3623
RX|3623,3625
*|3626,3627
enoxaparin|3627,3637
40|3638,3640
mg|3641,3643
/|3643,3644
0.4|3644,3647
mL|3648,3650
40|3651,3653
mg|3654,3656
subq|3657,3661
daily|3662,3667
Disp|3668,3672
#|3673,3674
*|3674,3675
14|3675,3677
Syringe|3678,3685
<EOL>|3686,3687
Refills|3687,3694
:|3694,3695
*|3695,3696
0|3696,3697
<EOL>|3697,3698
13.|3698,3701
Milk|3702,3706
of|3707,3709
Magnesia|3710,3718
30|3719,3721
ml|3722,3724
PO|3725,3727
BID|3728,3731
:|3731,3732
PRN|3732,3735
Dyspepsia|3736,3745
<EOL>|3746,3747
14.|3747,3750
Multivitamins|3751,3764
1|3765,3766
CAP|3767,3770
PO|3771,3773
DAILY|3774,3779
<EOL>|3780,3781
15.|3781,3784
OxycoDONE|3785,3794
(|3795,3796
Immediate|3796,3805
Release|3806,3813
)|3813,3814
2.5|3816,3819
mg|3820,3822
PO|3823,3825
Q6H|3826,3829
:|3829,3830
PRN|3830,3833
pain|3834,3838
<EOL>|3839,3840
RX|3840,3842
*|3843,3844
oxycodone|3844,3853
5|3854,3855
mg|3856,3858
_|3859,3860
_|3860,3861
_|3861,3862
tablet|3863,3869
(|3869,3870
s|3870,3871
)|3871,3872
by|3873,3875
mouth|3876,3881
every|3882,3887
four|3888,3892
hours|3893,3898
Disp|3899,3903
<EOL>|3904,3905
#|3905,3906
*|3906,3907
60|3907,3909
Tablet|3910,3916
Refills|3917,3924
:|3924,3925
*|3925,3926
0|3926,3927
<EOL>|3927,3928
16|3928,3930
.|3930,3931
Pantoprazole|3932,3944
40|3945,3947
mg|3948,3950
PO|3951,3953
Q24H|3954,3958
<EOL>|3959,3960
17.|3960,3963
Senna|3964,3969
2|3970,3971
TAB|3972,3975
PO|3976,3978
HS|3979,3981
<EOL>|3982,3983
18.|3983,3986
Vitamin|3987,3994
D|3995,3996
800|3997,4000
UNIT|4001,4005
PO|4006,4008
DAILY|4009,4014
<EOL>|4015,4016
<EOL>|4016,4017
<EOL>|4018,4019
Discharge|4019,4028
Disposition|4029,4040
:|4040,4041
<EOL>|4041,4042
Extended|4042,4050
Care|4051,4055
<EOL>|4055,4056
<EOL>|4057,4058
Facility|4058,4066
:|4066,4067
<EOL>|4067,4068
_|4068,4069
_|4069,4070
_|4070,4071
<EOL>|4071,4072
<EOL>|4073,4074
Discharge|4074,4083
Diagnosis|4084,4093
:|4093,4094
<EOL>|4094,4095
left|4095,4099
femoral|4100,4107
neck|4108,4112
fracture|4113,4121
<EOL>|4121,4122
<EOL>|4122,4123
<EOL>|4124,4125
Discharge|4125,4134
Condition|4135,4144
:|4144,4145
<EOL>|4145,4146
Mental|4146,4152
Status|4153,4159
:|4159,4160
Clear|4161,4166
and|4167,4170
coherent|4171,4179
.|4179,4180
<EOL>|4180,4181
Level|4181,4186
of|4187,4189
Consciousness|4190,4203
:|4203,4204
Alert|4205,4210
and|4211,4214
interactive|4215,4226
.|4226,4227
<EOL>|4227,4228
Activity|4228,4236
Status|4237,4243
:|4243,4244
Out|4245,4248
of|4249,4251
Bed|4252,4255
with|4256,4260
assistance|4261,4271
to|4272,4274
chair|4275,4280
or|4281,4283
<EOL>|4284,4285
wheelchair|4285,4295
.|4295,4296
<EOL>|4296,4297
<EOL>|4297,4298
<EOL>|4299,4300
Discharge|4300,4309
Instructions|4310,4322
:|4322,4323
<EOL>|4323,4324
MEDICATIONS|4324,4335
:|4335,4336
<EOL>|4336,4337
<EOL>|4337,4338
-|4338,4339
Please|4340,4346
take|4347,4351
all|4352,4355
medications|4356,4367
as|4368,4370
prescribed|4371,4381
by|4382,4384
your|4385,4389
physicians|4390,4400
<EOL>|4401,4402
at|4402,4404
discharge|4405,4414
.|4414,4415
<EOL>|4415,4416
<EOL>|4416,4417
-|4417,4418
Continue|4419,4427
all|4428,4431
home|4432,4436
medications|4437,4448
unless|4449,4455
specifically|4456,4468
instructed|4469,4479
<EOL>|4480,4481
to|4481,4483
stop|4484,4488
by|4489,4491
your|4492,4496
surgeon|4497,4504
.|4504,4505
<EOL>|4505,4506
<EOL>|4506,4507
-|4507,4508
Do|4509,4511
not|4512,4515
drink|4516,4521
alcohol|4522,4529
,|4529,4530
drive|4531,4536
a|4537,4538
motor|4539,4544
vehicle|4545,4552
,|4552,4553
or|4554,4556
operate|4557,4564
<EOL>|4565,4566
machinery|4566,4575
while|4576,4581
taking|4582,4588
narcotic|4589,4597
pain|4598,4602
relievers|4603,4612
.|4612,4613
<EOL>|4613,4614
<EOL>|4614,4615
-|4615,4616
Narcotic|4617,4625
pain|4626,4630
relievers|4631,4640
can|4641,4644
cause|4645,4650
constipation|4651,4663
,|4663,4664
so|4665,4667
you|4668,4671
should|4672,4678
<EOL>|4679,4680
drink|4680,4685
eight|4686,4691
8oz|4692,4695
glasses|4696,4703
of|4704,4706
water|4707,4712
daily|4713,4718
and|4719,4722
take|4723,4727
a|4728,4729
stool|4730,4735
softener|4736,4744
<EOL>|4745,4746
(|4746,4747
colace|4747,4753
)|4753,4754
to|4755,4757
prevent|4758,4765
this|4766,4770
side|4771,4775
effect|4776,4782
.|4782,4783
<EOL>|4783,4784
<EOL>|4784,4785
<EOL>|4786,4787
<EOL>|4787,4788
ANTICOAGULATION|4788,4803
:|4803,4804
<EOL>|4804,4805
<EOL>|4805,4806
-|4806,4807
Please|4808,4814
take|4815,4819
lovenox|4820,4827
40mg|4828,4832
daily|4833,4838
for|4839,4842
2|4843,4844
weeks|4845,4850
<EOL>|4850,4851
<EOL>|4851,4852
<EOL>|4853,4854
<EOL>|4854,4855
WOUND|4855,4860
CARE|4861,4865
:|4865,4866
<EOL>|4866,4867
<EOL>|4867,4868
-|4868,4869
You|4870,4873
can|4874,4877
get|4878,4881
the|4882,4885
wound|4886,4891
wet|4892,4895
/|4895,4896
take|4896,4900
a|4901,4902
shower|4903,4909
starting|4910,4918
3|4919,4920
days|4921,4925
after|4926,4931
<EOL>|4932,4933
your|4933,4937
surgery|4938,4945
.|4945,4946
You|4948,4951
may|4952,4955
wash|4956,4960
gently|4961,4967
with|4968,4972
soap|4973,4977
and|4978,4981
water|4982,4987
,|4987,4988
and|4989,4992
pat|4993,4996
<EOL>|4997,4998
the|4998,5001
incision|5002,5010
dry|5011,5014
after|5015,5020
showering|5021,5030
.|5030,5031
<EOL>|5033,5034
<EOL>|5034,5035
-|5035,5036
No|5037,5039
baths|5040,5045
or|5046,5048
swimming|5049,5057
for|5058,5061
at|5062,5064
least|5065,5070
4|5071,5072
weeks|5073,5078
.|5078,5079
<EOL>|5079,5080
<EOL>|5080,5081
-|5081,5082
Any|5083,5086
stitches|5087,5095
or|5096,5098
staples|5099,5106
that|5107,5111
need|5112,5116
to|5117,5119
be|5120,5122
removed|5123,5130
will|5131,5135
be|5136,5138
taken|5139,5144
<EOL>|5145,5146
out|5146,5149
at|5150,5152
your|5153,5157
2|5158,5159
-|5159,5160
week|5160,5164
follow|5165,5171
up|5172,5174
appointment|5175,5186
.|5186,5187
<EOL>|5187,5188
<EOL>|5188,5189
-|5189,5190
No|5191,5193
dressing|5194,5202
is|5203,5205
needed|5206,5212
if|5213,5215
wound|5216,5221
continues|5222,5231
to|5232,5234
be|5235,5237
non-draining|5238,5250
.|5250,5251
<EOL>|5251,5252
<EOL>|5252,5253
<EOL>|5254,5255
<EOL>|5255,5256
ACTIVITY|5256,5264
AND|5265,5268
WEIGHT|5269,5275
BEARING|5276,5283
:|5283,5284
<EOL>|5284,5285
<EOL>|5285,5286
touch|5286,5291
-|5291,5292
down|5292,5296
weight|5297,5303
-|5303,5304
bearing|5304,5311
LLE|5312,5315
<EOL>|5315,5316
Physical|5316,5324
Therapy|5325,5332
:|5332,5333
<EOL>|5333,5334
Touch|5334,5339
-|5339,5340
down|5340,5344
weight|5345,5351
bearing|5352,5359
LLE|5360,5363
<EOL>|5363,5364
Treatments|5364,5374
Frequency|5375,5384
:|5384,5385
<EOL>|5385,5386
WOUND|5386,5391
CARE|5392,5396
:|5396,5397
<EOL>|5397,5398
<EOL>|5398,5399
-|5399,5400
You|5401,5404
can|5405,5408
get|5409,5412
the|5413,5416
wound|5417,5422
wet|5423,5426
/|5426,5427
take|5427,5431
a|5432,5433
shower|5434,5440
starting|5441,5449
3|5450,5451
days|5452,5456
after|5457,5462
<EOL>|5463,5464
your|5464,5468
surgery|5469,5476
.|5476,5477
You|5479,5482
may|5483,5486
wash|5487,5491
gently|5492,5498
with|5499,5503
soap|5504,5508
and|5509,5512
water|5513,5518
,|5518,5519
and|5520,5523
pat|5524,5527
<EOL>|5528,5529
the|5529,5532
incision|5533,5541
dry|5542,5545
after|5546,5551
showering|5552,5561
.|5561,5562
<EOL>|5564,5565
<EOL>|5565,5566
-|5566,5567
No|5568,5570
baths|5571,5576
or|5577,5579
swimming|5580,5588
for|5589,5592
at|5593,5595
least|5596,5601
4|5602,5603
weeks|5604,5609
.|5609,5610
<EOL>|5610,5611
<EOL>|5611,5612
-|5612,5613
Any|5614,5617
stitches|5618,5626
or|5627,5629
staples|5630,5637
that|5638,5642
need|5643,5647
to|5648,5650
be|5651,5653
removed|5654,5661
will|5662,5666
be|5667,5669
taken|5670,5675
<EOL>|5676,5677
out|5677,5680
at|5681,5683
your|5684,5688
2|5689,5690
-|5690,5691
week|5691,5695
follow|5696,5702
up|5703,5705
appointment|5706,5717
.|5717,5718
<EOL>|5718,5719
<EOL>|5719,5720
-|5720,5721
No|5722,5724
dressing|5725,5733
is|5734,5736
needed|5737,5743
if|5744,5746
wound|5747,5752
continues|5753,5762
to|5763,5765
be|5766,5768
non-draining|5769,5781
.|5781,5782
<EOL>|5782,5783
<EOL>|5783,5784
<EOL>|5785,5786
Followup|5786,5794
Instructions|5795,5807
:|5807,5808
<EOL>|5808,5809
_|5809,5810
_|5810,5811
_|5811,5812
<EOL>|5812,5813

