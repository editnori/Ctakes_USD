CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Locally Advanced Gastric Carcinoma|Disorder|false|false|C0038351|Locally advanced gastric carcinomanull|Locally|Modifier|false|false||Locallynull|Stomach Carcinoma|Disorder|false|false|C0038351|gastric carcinomanull|Stomach|Anatomy|false|false|C5206813;C0699791|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Carcinoma|Disorder|false|false||carcinomanull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cystoscopy|Procedure|false|false||Cystoscopynull|Foley catheter|Device|false|false||foley catheternull|Catheter placement|Procedure|false|false||catheter placementnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Therapeutic Laparoscopy|Procedure|false|false||Laparoscopy
null|Laparoscopy|Procedure|false|false||Laparoscopynull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Endoscopy of stomach|Procedure|false|false||Gastroscopynull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|Locally|Modifier|false|false||locallynull|Stomach|Anatomy|false|false||gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Cure (remedy)|Finding|false|false||curativenull|Curative - procedure intent|Procedure|false|false||curativenull|Act Mood - intent|Finding|false|false||intent
null|null|Finding|false|false||intentnull|intent|Modifier|false|false||intentnull|removal technique|Procedure|false|false||surgical resection
null|Excision|Procedure|false|false||surgical resectionnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|completion - ResponseLevel|Modifier|false|false||completion
null|Complete|Modifier|false|false||completionnull|Induce (action)|Finding|false|false||inductionnull|Induction procedure|Procedure|false|false||inductionnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Neoadjuvant Chemotherapy|Procedure|false|false||neoadjuvant chemotherapynull|Neoadjuvant Therapy|Procedure|false|false||neoadjuvantnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Overall Publication Type|Finding|false|false||Overallnull|Overall|Modifier|false|false||Overallnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|aspects of adverse effects|Finding|false|false||side effects
null|Adverse effects|Finding|false|false||side effectsnull|Side|Modifier|false|false||sidenull|Effect|Modifier|false|false||effectsnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Right upper extremity|Anatomy|false|false|C0085649;C0522035;C1552823;C0013604|right upper extremitynull|Table Cell Horizontal Align - right|Finding|false|false|C1140618;C0230329|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Edema of the upper extremity|Finding|false|false|C0015385;C1140618;C0230329|upper extremity edemanull|Upper Extremity|Anatomy|false|false|C0522035;C0085649;C1552823;C0013604|upper extremitynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Peripheral edema|Finding|false|false|C0230329;C1140618;C0015385|extremity edemanull|Limb structure|Anatomy|false|false|C0522035;C0013604;C0085649|extremitynull|Edema|Finding|false|false|C0015385;C1140618;C0230329|edemanull|null|Attribute|false|false||edemanull|Thrombosis|Finding|false|false||thrombosisnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|ug/g|LabModifier|false|false||mg/kgnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Compliance behavior|Finding|false|false||compliantnull|Compliant (qualifier value)|Modifier|false|false||compliantnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Chills|Finding|false|false||chillsnull|Weight Loss|Finding|false|false||weight loss
null|Losing Weight (question)|Finding|false|false||weight lossnull|Measured weight loss (observable entity)|LabModifier|false|false||weight lossnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Melena|Finding|false|false||melenanull|Hematochezia|Disorder|false|false||hematochezianull|Blood in stool|Finding|false|false||hematochezianull|Hematuria|Disorder|false|false||hematurianull|Recent|Time|false|false||recentnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|With staging|Finding|false|false||stagingnull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Disease|Disorder|true|false||diseasenull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Invasive|Modifier|false|false||invasivenull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Open|Modifier|false|false||opennull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Partial gastrectomy with anastomosis to duodenum|Procedure|false|false||distal gastrectomy
null|Billroth I Procedure|Procedure|false|false||distal gastrectomynull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Gastrectomy|Procedure|false|false||gastrectomynull|Lymph node excision|Procedure|false|false||lymphadenectomynull|Risk|Finding|false|false||risksnull|Benefit|LabModifier|false|false||benefitsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|detail - Response Level|Finding|false|false||detailnull|Details|Modifier|false|false||detailnull|Separate|Modifier|false|false||separatenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|Prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|Prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|Prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|Prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|Prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|Prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0006826;C0376358;C0600139;C0496923;C0154088;C0033575;C0154009|Prostate
null|Prostate|Anatomy|false|false|C0006826;C0376358;C0600139;C0496923;C0154088;C0033575;C0154009|Prostatenull|Thyroid carcinoma|Disorder|false|false|C0040132|cancer, Thyroidnull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Thyroid Nodule|Disorder|false|false|C0040132|Thyroid nodulenull|null|Finding|false|false|C0040132|Thyroid nodulenull|THYROID DIAGNOSTIC RADIOPHARMACEUTICALS|Drug|false|false|C0040132|Thyroid
null|THYROID|Drug|false|false|C0040132|Thyroid
null|THYROID|Drug|false|false|C0040132|Thyroid
null|thyroid (USP)|Drug|false|false|C0040132|Thyroid
null|thyroid (USP)|Drug|false|false|C0040132|Thyroid
null|thyroid (USP)|Drug|false|false|C0040132|Thyroidnull|Thyroid Diseases|Disorder|false|false|C0040132|Thyroidnull|examination of thyroid|Procedure|false|false|C0040132|Thyroidnull|Thyroid Gland|Anatomy|false|false|C0549473;C0040137;C2116082;C3540038;C0040134;C5781115;C2228489;C0040128|Thyroidnull|Hypothyroidism|Disorder|false|false||Hypothyroidnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Diverticulosis|Disorder|false|false||Diverticulosisnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|butyl phosphorotrithioate|Drug|false|false||def
null|butyl phosphorotrithioate|Drug|false|false||defnull|UTP25 gene|Finding|false|false||defnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|History of surgery|Finding|false|false||Past Surgical Historynull|history of prior surgery|Finding|false|false||Surgical Historynull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527;C1548801|Prostate cancer
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527;C1548801|Prostate cancernull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|Prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|Prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|Prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|Prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009;C0376358;C0600139;C0006826|Prostate
null|Prostate|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009;C0376358;C0600139;C0006826|Prostatenull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527;C1548801|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|External route|Finding|false|false|C1548801|externalnull|Body Site Modifier - External|Anatomy|false|false|C0521134;C0376358;C0600139;C0338248;C0006826|externalnull|Code System Type - External|Modifier|false|false||external
null|External|Modifier|false|false||externalnull|Beam -- chemical|Drug|false|false||beam
null|Beam -- chemical|Drug|false|false||beamnull|carmustine/cytarabine/etoposide/melphalan regimen|Procedure|false|false|C1548801|beamnull|Beam - rays of radiation or stream of particles|Phenomenon|false|false||beamnull|Repair of Achilles tendon|Procedure|false|false|C0001074;C0001074;C1305378;C0817321;C0039508|Achilles tendon repairnull|Structure of achilles tendon|Anatomy|false|false|C0043240;C4319951;C0407029;C0565350;C0374711;C1705181|Achilles tendon
null|null|Anatomy|false|false|C0043240;C4319951;C0407029;C0565350;C0374711;C1705181|Achilles tendonnull|Structure of achilles tendon|Anatomy|false|false|C0374711;C1705181;C0407029;C0565350;C0043240;C4319951|Achillesnull|Plastic repair of tendon|Procedure|false|false|C0817321;C0001074;C0001074;C1305378;C0039508|tendon repairnull|Tendon structure|Anatomy|false|false|C0043240;C4319951;C0374711;C1705181;C0407029;C0565350|tendonnull|Repair|Finding|false|false|C0001074;C1305378;C0039508;C0817321;C0001074|repair
null|Wound Healing|Finding|false|false|C0001074;C1305378;C0039508;C0817321;C0001074|repairnull|Repair - Remedial Action|Procedure|false|false|C0001074;C0039508;C0817321;C0001074;C1305378|repair
null|Surgical repair|Procedure|false|false|C0001074;C0039508;C0817321;C0001074;C1305378|repairnull|Right tibia|Anatomy|false|false|C0565350;C0407029;C0043240;C4319951;C1552823;C0374711;C1705181|right tibianull|Table Cell Horizontal Align - right|Finding|false|false|C0817321|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|tibia and fibula|Anatomy|false|false||tibia and fibulanull|Bone structure of tibia|Anatomy|false|false||tibianull|Tibia <Rostellariidae>|Entity|false|false||tibianull|Fibula|Anatomy|false|false||fibulanull|Tonsillectomy|Procedure|false|false||Tonsillectomynull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Lymphoma|Disorder|false|false||Lymphomanull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|null|Modifier|false|false||with typenull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Data|Finding|false|false||Datanull|Data call receiving device|Device|false|false||Datanull|Data <Amphipyrinae>|Entity|false|false||Datanull|Last|Modifier|false|false||lastnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|scleranull|examination of sclera|Procedure|false|false|C0036410|scleranull|Sclera|Anatomy|false|false|C0205180;C0036412;C2228481|scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|Respiratory distress|Finding|true|false||respiratory distressnull|Respiratory attachment|Finding|true|false||respiratory
null|respiratory|Finding|true|false||respiratory
null|null|Finding|true|false||respiratory
null|Respiratory specimen|Finding|true|false||respiratorynull|Respiratory rate|Attribute|true|false||respiratorynull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Psychiatric problem|Disorder|false|false||PSYCH
null|Mental disorders|Disorder|false|false||PSYCHnull|Insight|Finding|false|false||insightnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Mood (psychological function)|Finding|false|false||mood
null|mood (physical finding)|Finding|false|false||mood
null|Mood (attribute)|Finding|false|false||moodnull|null|Attribute|false|false||moodnull|Traumatic Wound|Disorder|false|false|C2338258|WOUND
null|Wounds and Injuries|Disorder|false|false|C2338258|WOUND
null|Traumatic injury|Disorder|false|false|C2338258|WOUNDnull|Route of Administration - Wound|Finding|false|false|C2338258|WOUND
null|null|Finding|false|false|C2338258|WOUND
null|Specimen Type - Wound|Finding|false|false|C2338258|WOUNDnull|Surgical wound|Disorder|false|false|C2338258|Incisionnull|Surgical incisions|Procedure|false|false|C2338258|Incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C1549529;C1547965;C1550680;C0184898;C3263723;C0043251;C0043250|Incisionnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Male Gender|Finding|false|false||Malenull|Male, Self-Reported|Subject|false|false||Male
null|Males|Subject|false|false||Malenull|Male Phenotype|Modifier|false|false||Malenull|Invasive|Modifier|false|false||invasivenull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Open|Modifier|false|false||opennull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Gastrectomy|Procedure|false|false||gastrectomynull|Lymph node excision|Procedure|false|false|C0038351|lymphadenectomynull|Locally|Modifier|false|false||locallynull|Stomach|Anatomy|false|false|C0024203|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Carcinoma|Disorder|false|false||carcinomanull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Quadrant|Modifier|false|false||quadrantnull|Port - alcoholic beverage|Drug|false|false||portnull|Implanted Port Access Device|Device|false|false||port
null|Port (physical object)|Device|false|false||port
null|Data Port|Device|false|false||port
null|Harbor|Device|false|false||portnull|Insufflation route|Finding|false|false||insufflationnull|Insufflation|Procedure|false|false|C0230177|insufflationnull|Structure of right upper quadrant of abdomen|Anatomy|false|false|C1552823;C0021634|right upper quadrantnull|RUQ - Right upper quadrant|Modifier|false|false||right upper quadrantnull|Table Cell Horizontal Align - right|Finding|false|false|C0230177|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Quadrant|Modifier|false|false||quadrantnull|Port - alcoholic beverage|Drug|false|false|C0028977|portnull|Implanted Port Access Device|Device|false|false||port
null|Port (physical object)|Device|false|false||port
null|Data Port|Device|false|false||port
null|Harbor|Device|false|false||portnull|Omentum|Anatomy|false|false|C0452253|omentumnull|Structure of transverse mesocolon|Anatomy|false|false|C5575035;C0750873;C0009373;C0154061;C0496907|transverse mesocolonnull|Anatomical transverse plane|Modifier|false|false||transverse
null|Transverse plane|Modifier|false|false||transversenull|Mesocolon|Anatomy|false|false|C5575035;C0750873;C0009373;C0154061;C0496907|mesocolonnull|Well (answer to question)|Finding|false|false|C0025483;C0230254|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0025483;C0230254|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0025483;C0230254|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0025483;C0230254|colonnull|COLON PROBLEM|Finding|false|false|C0025483;C0230254;C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Obvious|Modifier|false|false||obviousnull|peritoneal|Anatomy|false|false|C0333562|peritoneal
null|Peritoneum|Anatomy|false|false|C0333562|peritonealnull|Deposition (morphologic abnormality)|Finding|false|false|C0442034;C0031153|depositsnull|peritoneal|Anatomy|false|false||peritoneal
null|Peritoneum|Anatomy|false|false||peritonealnull|Four quadrants|Modifier|false|false||four quadrantsnull|carcinomatosis of unspecified behavior|Disorder|false|false||carcinomatosis
null|Carcinomatosis|Disorder|false|false||carcinomatosisnull|Bad|Modifier|false|false||poorlynull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Neoplasm of uncertain or unknown behavior of peritoneum|Disorder|false|false|C0031153;C4482223;C0230198|peritoneum
null|Benign neoplasm of peritoneum|Disorder|false|false|C0031153;C4482223;C0230198|peritoneumnull|Serous layer of peritoneum|Anatomy|false|false|C0496874;C0496954|peritoneum
null|Peritoneum|Anatomy|false|false|C0496874;C0496954|peritoneum
null|Abdomen>Peritoneum|Anatomy|false|false|C0496874;C0496954|peritoneumnull|Indication of (contextual qualifier)|Finding|false|false||reasonnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Ward (environment)|Device|false|false||wardsnull|Ward (environment)|Entity|false|false||wardsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Hospitalization|Procedure|false|false||hospitalizationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Initially|Time|false|false||initiallynull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCAnull|Posterior cortical atrophy syndrome|Disorder|false|false|C0149576|PCA
null|Familial lichen amyloidosis|Disorder|false|false|C0149576|PCAnull|PCA Message Structure|Finding|false|false|C0149576|PCA
null|CHOANAL ATRESIA, POSTERIOR|Finding|false|false|C0149576|PCA
null|FLVCR1 gene|Finding|false|false|C0149576|PCAnull|Patient controlled intravenous analgesia|Procedure|false|false|C0149576|PCA
null|Passive Cutaneous Anaphylaxis|Procedure|false|false|C0149576|PCA
null|Patient-Controlled Analgesia|Procedure|false|false|C0149576|PCAnull|Structure of posterior cerebral artery|Anatomy|false|false|C0034330;C0030131;C0268398;C4275079;C0220723;C1836722;C1549860;C0078944;C5968782;C0030625|PCAnull|Principal Component Analysis|LabModifier|false|false||PCAnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Describes Very Well|Finding|false|false||very well
null|Can Do Very Well|Finding|false|false||very well
null|Very Well|Finding|false|false||very wellnull|Very good (qualifier value)|Modifier|false|false||very wellnull|Very|Modifier|false|false||verynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Cardiovascular system|Anatomy|false|false||cardiovascular
null|Cardiovascular|Anatomy|false|false||cardiovascularnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Pulmonary (intended site)|Finding|false|false|C0024109|PULMONARYnull|Lung|Anatomy|false|false|C4522268;C2707265|PULMONARYnull|null|Attribute|false|false|C0024109|PULMONARYnull|Pulmonary (qualifier value)|Modifier|false|false||PULMONARYnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Language Ability Proficiency - Good|Finding|false|false|C0024109|Good
null|Language Proficiency - Good|Finding|false|false|C0024109|Goodnull|Specimen Quality - Good|Modifier|false|false||Good
null|Good|Modifier|false|false||Goodnull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C1610541;C1551023;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Toilet procedure|Procedure|false|false||toiletnull|Commodes|Device|false|false||toiletnull|Early Ambulation|Procedure|false|false||early ambulationnull|Early|Time|false|false||earlynull|Ambulation|Finding|false|false||ambulation
null|Walking (function)|Finding|false|false||ambulationnull|Incentive spirometry|Procedure|false|false||incentive spirometrynull|Incentives|Modifier|false|false||incentivenull|Spirometry|Procedure|false|false||spirometrynull|Hospitalization|Procedure|false|false||hospitalizationnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Nurses|Subject|false|false||nursenull|Unable|Finding|false|false||unablenull|Pass (indicator)|Finding|false|false||passnull|Attempt|Event|false|false||attemptnull|Type of Agreement - Standard|Finding|false|false||standard
null|Standard (document)|Finding|false|false||standardnull|Standard base excess calculation technique|Procedure|false|false||standardnull|Standard (qualifier)|Modifier|false|false||standardnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Usual|Modifier|false|false||usualnull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Techniques|Finding|false|false||techniquenull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|HL7 Version 2.5 - Application|Finding|false|false||application
null|Application Document|Finding|false|false||application
null|Computer Application|Finding|false|false||application
null|Regulatory Application|Finding|false|false||application
null|Apply|Finding|false|false||applicationnull|Application procedure|Procedure|false|false||applicationnull|Application - unit of product usage|LabModifier|false|false||applicationnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|catheter device|Device|false|false||cathetersnull|Unable|Finding|false|false||unablenull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009|prostatenull|Urology|Title|false|false||Urologynull|Flexible|Modifier|false|false||flexiblenull|Cystoscopes|Device|false|false||cystoscopenull|Neoplasm of uncertain or unknown behavior of urethra|Disorder|false|false|C0041967|urethra
null|Urethral Diseases|Disorder|false|false|C0041967|urethra
null|Benign neoplasm of urethra|Disorder|false|false|C0041967|urethra
null|Malignant neoplasm of urethra|Disorder|false|false|C0041967|urethranull|Urethra specimen code|Finding|false|false|C0041967|urethra
null|Urethra specimen|Finding|false|false|C0041967|urethranull|Procedure on urethra|Procedure|false|false|C0041967|urethranull|Urethra|Anatomy|false|false|C0153620;C0041969;C0496929;C0154019;C0810170;C1550675;C1547951|urethranull|Flexible|Modifier|false|false||flexiblenull|Guidewire Device|Device|false|false||guidewirenull|Cystoscopes|Device|false|false||cystoscopenull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0872388;C0496930;C0154017;C0154091|bladdernull|Scope|Finding|false|false||scopenull|Council (ethnic group)|Subject|false|false||councilnull|WIPF2 gene|Finding|false|false||wirenull|Wire Device|Device|false|false||wire
null|Bone Wires|Device|false|false||wirenull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0005682;C0033572;C4266527|prostate
null|Prostatic Diseases|Disorder|false|false|C0005682;C0033572;C4266527|prostate
null|Carcinoma in situ of prostate|Disorder|false|false|C0005682;C0033572;C4266527|prostate
null|Benign neoplasm of prostate|Disorder|false|false|C0005682;C0033572;C4266527|prostatenull|Structure of prostate (body structure)|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009|prostate
null|Prostate|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009|prostatenull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496923;C0154088;C0033575;C0154009;C0872388;C0496930;C0154017;C0154091|bladdernull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Urology|Title|false|false||urologynull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|Urination|Finding|false|false||voiding
null|Voids|Finding|false|false||voidingnull|Clinical Trials|Procedure|false|false||trialnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|true|false||antibiotics
null|Antibiotics|Drug|true|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|true|false||antibiotics
null|Antibiotics, Gynecological|Drug|true|false||antibiotics
null|antibiotics, intestinal|Drug|true|false||antibiotics
null|Antibiotic throat preparations|Drug|true|false||antibiotics
null|Antibiotics, Antitubercular|Drug|true|false||antibiotics
null|Antibiotics for systemic use|Drug|true|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|true|false||antibioticsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Heme|Drug|false|false||HEME
null|Heme|Drug|false|false||HEMEnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C5239664|BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|DVT prophylaxis|Procedure|false|false|C5239664|DVT prophylaxisnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2926618;C0199176;C0853245;C4546282|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Prophylactic treatment|Procedure|false|false|C5239664|prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Early Ambulation|Procedure|false|false||early ambulationnull|Early|Time|false|false||earlynull|Ambulation|Finding|false|false||ambulation
null|Walking (function)|Finding|false|false||ambulationnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Medical Devices|Device|false|false||devices
null|device aspects|Device|false|false||devices
null|Devices|Device|false|false||devicesnull|TCF21 wt Allele|Finding|false|false||POD1
null|CORO7 gene|Finding|false|false||POD1
null|TCF21 gene|Finding|false|false||POD1null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Foley catheter|Device|false|false||Foley catheternull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Appropriate|Modifier|false|false||appropriatenull|Visit User Code - Teaching|Finding|false|false||teachingnull|Teaching aspects|Procedure|false|false||teaching
null|Education (procedure)|Procedure|false|false||teachingnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Teaching|Finding|false|false||teachingnull|Teaching aspects|Procedure|false|false||teaching
null|Education (procedure)|Procedure|false|false||teachingnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Comprehension|Finding|false|false||understandingnull|Agreement (document)|Finding|false|false||agreement
null|Agreement|Finding|false|false||agreementnull|null|Attribute|false|false||agreementnull|Discharge plan|Finding|false|false||discharge plannull|Discharge Planning|Procedure|false|false||discharge plannull|null|Attribute|false|false||discharge plannull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|prescription document|Finding|false|false||Prescriptionnull|Prescription (procedure)|Procedure|false|false||Prescriptionnull|Prescription (attribute)|Attribute|false|false||Prescriptionnull|Bio-Throid|Drug|false|false||BIO-THROID
null|Bio-Throid|Drug|false|false||BIO-THROID
null|Bio-Throid|Drug|false|false||BIO-THROIDnull|Bio-Throid|Drug|false|false||Bio-Throid
null|Bio-Throid|Drug|false|false||Bio-Throid
null|Bio-Throid|Drug|false|false||Bio-Throidnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|enoxaparin|Drug|false|false||ENOXAPARIN
null|enoxaparin|Drug|false|false||ENOXAPARINnull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Syringes|Device|false|false||syringenull|Syringe (unit of presentation)|LabModifier|false|false||syringe
null|Syringe Dosing Unit|LabModifier|false|false||syringenull|Daily|Time|false|false||dailynull|omeprazole|Drug|false|false||OMEPRAZOLE
null|omeprazole|Drug|false|false||OMEPRAZOLEnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|ubiquinol|Drug|false|false||UBIQUINOL
null|ubiquinol|Drug|false|false||UBIQUINOLnull|ubiquinol|Drug|false|false||ubiquinol
null|ubiquinol|Drug|false|false||ubiquinolnull|Oral cavity|Anatomy|false|false|C1561538;C1561539|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Drugs, Non-Prescription|Drug|false|false||OTCnull|OTC gene|Finding|false|false||OTCnull|ferrous sulfate|Drug|false|false||FERROUS SULFATE
null|ferrous sulfate|Drug|false|false||FERROUS SULFATEnull|Ferrous|Drug|false|false||FERROUSnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATE
null|Sulfates, Inorganic|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|sulfate ion|Drug|false|false||SULFATE
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||SULFATEnull|ferrous sulfate|Drug|false|false||ferrous sulfate
null|ferrous sulfate|Drug|false|false||ferrous sulfatenull|Ferrous|Drug|false|false||ferrousnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Lactobacillus combination no.4|Entity|false|false||LACTOBACILLUS COMBINATION NO.4null|Lactobacillus|Entity|false|false||LACTOBACILLUSnull|combination - answer to question|Finding|false|false||COMBINATIONnull|combination of objects|Entity|false|false||COMBINATIONnull|Combined|Modifier|false|false||COMBINATIONnull|Probiotics|Entity|false|false||PROBIOTICnull|Dosage|LabModifier|false|false||Dosagenull|Uncertainty|Finding|false|false||uncertainnull|Transaction counts and value totals - provider|Finding|false|false||Provider
null|Provider|Finding|false|false||Providernull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Low dose|LabModifier|false|false||low dosenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Constipation|Finding|false|false||constipationnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Malignant neoplasm of stomach stage IV|Disorder|false|false|C0038351|Metastatic gastric cancernull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Malignant neoplasm of stomach|Disorder|false|false|C0038351|gastric cancer
null|Stomach Carcinoma|Disorder|false|false|C0038351|gastric cancernull|Stomach|Anatomy|false|false|C0278498;C0024623;C0699791;C0006826|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Malignant Neoplasms|Disorder|false|false|C0038351|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Urethral Stenosis|Disorder|false|false|C0041967|Urethral stricturenull|Urethral stricture|Finding|false|false|C0041967|Urethral stricturenull|Urethral Dosage Form|Drug|false|false|C0041967|Urethralnull|Intraurethral Route of Administration|Finding|false|false|C0041967|Urethralnull|Urethra|Anatomy|false|false|C1522518;C1261287;C0041974;C2349082;C4551691|Urethralnull|Urethral (intended site)|Modifier|false|false||Urethralnull|Stenosis|Finding|false|false|C0041967|stricturenull|Stenosis Morphology|Modifier|false|false||stricturenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Malignant neoplasm of stomach|Disorder|false|false|C0038351|gastric cancer
null|Stomach Carcinoma|Disorder|false|false|C0038351|gastric cancernull|Stomach|Anatomy|false|false|C0024623;C0699791;C0006826|gastricnull|Gastric (qualifier value)|Modifier|false|false||gastricnull|Malignant Neoplasms|Disorder|false|false|C0038351|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Robot Device|Device|false|false||Robot
null|null|Device|false|false||Robotnull|Laparoscopy|Procedure|false|false||laparoscopicnull|Laparoscopic approach|Modifier|false|false||laparoscopicnull|Subtotal gastrectomy|Procedure|false|false||partial gastrectomynull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Gastrectomy|Procedure|false|false||gastrectomynull|Endoscopy of stomach|Procedure|false|false||gastroscopynull|complication aspects|Finding|true|false||complications
null|Complication|Finding|true|false||complicationsnull|null|Attribute|true|false||complicationsnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Feces|Finding|false|false||stoolingnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false|C0230028;C0226896|pain
null|Pain|Finding|false|false|C0230028;C0226896|painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false|C0230028;C0226896|medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1549543;C0030193;C4284232;C1527415|mouth
null|Oral region|Anatomy|false|false|C1549543;C0030193;C4284232;C1527415|mouthnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Recommendation|Finding|false|false||recommendationsnull|Uneventful|Finding|false|false||uneventfulnull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Activity (animal life circumstance)|Finding|false|false||ACTIVITY
null|Physical activity|Finding|false|false||ACTIVITYnull|Activities|Event|false|false||ACTIVITYnull|null|Modifier|false|false||ACTIVITYnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Prior functioning.stairs|Finding|false|false||stairsnull|Several|LabModifier|false|false||severalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Distance|LabModifier|false|false||distancesnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Visit|Finding|false|false||visitnull|Light Exercise|Finding|false|false||light exercisenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Feeling comfortable|Finding|false|false||comfortablenull|Slow|Modifier|false|false||Slowlynull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Heavy (weight) (qualifier value)|Modifier|false|false||Heavy
null|Heavy (amount)|Modifier|false|false||Heavynull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Sensory perception|Finding|false|false||sensenull|Slow|Modifier|false|false||slowlynull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|true|false||liftingnull|10 pounds|Finding|true|false||10 poundsnull|Pounds|LabModifier|false|false||poundsnull|More|LabModifier|false|false||morenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Sexual Activity|Finding|false|false||sexual activity
null|Sex Behavior|Finding|false|false||sexual activitynull|Sex Behavior|Finding|false|false||sexualnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Feelings|Finding|false|false||FEELnull|Feel Weak (question)|Finding|false|false||feel weak
null|Weakness|Finding|false|false||feel weaknull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Neutrophil Activation Probe Imaging Agent|Drug|false|false||napnull|CTNNBL1 gene|Finding|false|false||nap
null|Napping|Finding|false|false||napnull|Neapolitan Language|Entity|false|false||napnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|LITAF gene|Finding|false|false||Simplenull|Simple|Modifier|false|false||Simplenull|exhaust|Drug|false|false||exhaustnull|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throatnull|Pharyngitis|Disorder|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore Throat|Finding|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore to touch|Finding|false|false||sore
null|Sore skin|Finding|false|false||sorenull|Sore sensation quality|Modifier|false|false||sorenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Anterior portion of neck|Anatomy|false|false|C0031350;C1950455;C3244654;C0723402;C0242429;C1550663;C1547926|throat
null|Throat|Anatomy|false|false|C0031350;C1950455;C3244654;C0723402;C0242429;C1550663;C1547926|throat
null|Pharyngeal structure|Anatomy|false|false|C0031350;C1950455;C3244654;C0723402;C0242429;C1550663;C1547926|throatnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Throat|Anatomy|false|false|C1550663;C1547926;C1950455;C0543467;C0038895;C1457907;C1547138|throat
null|Anterior portion of neck|Anatomy|false|false|C1550663;C1547926;C1950455;C0543467;C0038895;C1457907;C1547138|throat
null|Pharyngeal structure|Anatomy|false|false|C1550663;C1547926;C1950455;C0543467;C0038895;C1457907;C1547138|throatnull|Level of Care - Surgery|Finding|false|false|C0230069;C3665375;C0031354|surgery
null|Surgical procedure finding|Finding|false|false|C0230069;C3665375;C0031354|surgery
null|Surgical aspects|Finding|false|false|C0230069;C3665375;C0031354|surgerynull|Operative Surgical Procedures|Procedure|false|false|C0230069;C3665375;C0031354|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Intestines|Anatomy|false|false||BOWELSnull|Constipation|Finding|false|false||Constipationnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Adverse effects|Finding|false|false||side effectnull|Side|Modifier|false|false||sidenull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Gentle Laxative|Drug|false|false||gentle laxative
null|Gentle Laxative|Drug|false|false||gentle laxativenull|Gentle|Drug|false|false||gentle
null|Gentle|Drug|false|false||gentlenull|Laxatives|Drug|false|false||laxativenull|cow milk allergenic extract|Drug|false|false||milk
null|Milk antigen|Drug|false|false||milk
null|Milk Beverage|Drug|false|false||milk
null|Plant-Based Milk|Drug|false|false||milk
null|cow milk allergenic extract|Drug|false|false||milk
null|Milk Specimen|Drug|false|false||milk
null|Cow's milk|Drug|false|false||milk
null|null|Drug|false|false||milknull|Milk (body substance)|Finding|false|false||milk
null|Milk Specimen Code|Finding|false|false||milknull|magnesium oxide|Drug|false|false||magnesia
null|magnesium oxide|Drug|false|false||magnesianull|Townes syndrome|Disorder|false|false||tbsnull|Toxicity Burden Score|Finding|false|false||tbs
null|SALL1 gene|Finding|false|false||tbs
null|SALL1 wt Allele|Finding|false|false||tbsnull|theta-burst stimulation|Procedure|false|false||tbsnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|prescription document|Finding|true|false||prescriptionnull|Prescription (procedure)|Procedure|true|false||prescriptionnull|Prescription (attribute)|Attribute|true|false||prescriptionnull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|Defecation|Finding|true|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|true|false||movementnull|Have Pain|Finding|false|false||have painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Intestines|Anatomy|false|false||bowelsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|ActInformationPrivacyReason - operations|Finding|false|false||operations
null|HL7PublishingSubSection - operations|Finding|false|false||operations
null|Surgical aspects|Finding|false|false||operationsnull|Operation Activity|Event|false|false||operationsnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Anti-Diarrhea|Drug|false|false||anti-diarrhea
null|Anti-Diarrhea|Drug|false|false||anti-diarrheanull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Feel Ill Question|Finding|false|false||feel ill
null|Malaise|Finding|false|false||feel ill
null|Feeling bad emotionally|Finding|false|false||feel illnull|Malaise|Finding|false|false||illnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Pain management (procedure)|Procedure|false|false||PAIN MANAGEMENTnull|Pain Management (specialty)|Title|false|false||PAIN MANAGEMENTnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Disease Management|Procedure|false|false||MANAGEMENTnull|Management Occupations|Subject|false|false||MANAGEMENTnull|Management procedure|Event|false|false||MANAGEMENT
null|Administration occupational activities|Event|false|false||MANAGEMENTnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|24 Hours|Time|false|false||24 hoursnull|Hour|Time|false|false||hoursnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Increase|Finding|false|false||increasenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Dosage|LabModifier|false|false||dosesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|Constipation|Finding|false|false||constipationnull|Slow|Modifier|false|false||Slowlynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Sharp pain|Finding|false|false||sharp painnull|Sharp sensation quality|Finding|false|false||sharp
null|SPEN wt Allele|Finding|false|false||sharp
null|SPEN gene|Finding|false|false||sharpnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Several|LabModifier|false|false||severalnull|Hour|Time|false|false||hoursnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C2926613;C1549543;C0030193;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C2926613;C1549543;C0030193;C0008031|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Tightness sensation quality|Modifier|false|false||tightnessnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Wheezing|Finding|false|false||wheezingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Nature|Finding|false|false||nature
null|Natures|Finding|false|false||naturenull|Quality|Modifier|false|false||qualitynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Nausea and vomiting|Finding|false|false||nausea and vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Dehydration|Disorder|false|false||dehydratednull|Xerostomia|Disorder|false|false|C0230028;C0226896|dry mouthnull|Oral cavity|Anatomy|false|false|C0795691;C0043352;C0425583;C0153957;C0153500|mouth
null|Oral region|Anatomy|false|false|C0795691;C0043352;C0425583;C0153957;C0153500|mouthnull|Tachycardia|Finding|false|false|C4037974;C0018787|rapid heart beatnull|Rapid|Modifier|false|false||rapidnull|Heart beat|Finding|false|false|C4037974;C0018787;C0230028;C0226896|heart beatnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787;C0230028;C0226896|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787;C0230028;C0226896|heartnull|HEART PROBLEM|Finding|false|false|C0230028;C0226896;C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0425583;C0795691;C0039231|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0425583;C0795691;C0039231|heartnull|feeling dizzy|Finding|false|false||feeling dizzynull|Dizziness|Finding|false|false||dizzynull|Faint - appearance|Finding|false|false||faint
null|Syncope|Finding|false|false||faintnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Additional|Finding|false|false||Additionalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|In Urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urine
null|Portion of urine|Finding|false|false||urinenull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONSnull|Medications|Finding|false|false||MEDICATIONSnull|null|Attribute|false|false||MEDICATIONS
null|null|Attribute|false|false||MEDICATIONSnull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Take|Procedure|false|false||takenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Wound care management|Procedure|false|false||WOUND CARE
null|wound care|Procedure|false|false||WOUND CAREnull|Wound Care kit|Device|false|false||WOUND CAREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|In care (finding)|Finding|false|false||CARE
null|Continuity Assessment Record and Evaluation|Finding|false|false||CAREnull|care activity|Event|false|false||CAREnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Wound Dressings (device)|Device|false|false||dressings
null|Medical dressing|Device|false|false||dressingsnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Bandage Dosage Form|Drug|false|false||bandagenull|Bandage|Device|false|false||bandagenull|strip medical device|Device|false|false||stripsnull|Swimming|Finding|false|false||swimnull|Fenamole|Drug|false|false||pat
null|Fenamole|Drug|false|false||patnull|Paroxysmal atrial tachycardia|Disorder|false|false||patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||pat
null|protein acetyltransferase activity|Finding|false|false||patnull|Thermoacoustic Computed Tomography|Procedure|false|false||patnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Steri-Strip|Device|false|false||steri stripsnull|Silene|Entity|false|false||sterinull|strip medical device|Device|false|false||stripsnull|week|Time|false|false||weeksnull|Still|Disorder|false|false||stillnull|Two weeks|Time|false|false||two weeksnull|week|Time|false|false||weeksnull|Along edge (qualifier value)|Modifier|false|false||edgesnull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|Soak Administration|Finding|false|false||soaknull|Soak (procedure)|Procedure|false|false||soaknull|Swimming|Finding|false|false||swimnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Surgical Team|Modifier|false|false||surgical teamnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Team|Subject|false|false||teamnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Smell Perception|Finding|false|false||smellingnull|Bloody|Finding|false|false||bloodynull|Hemorrhagic|Modifier|false|false||bloodynull|Pus specimen|Drug|false|false||pusnull|Pus Specimen Code|Finding|false|false||pus
null|Pus|Finding|false|false||pusnull|Pashtu language|Entity|false|false||pusnull|Etc.|Finding|false|false||etcnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Site of incision|Modifier|false|false||incision sitenull|Surgical wound|Disorder|false|false|C1515974;C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258;C1515974|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0332803;C1546778;C0184898|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Opening|Modifier|false|false||opening
null|Open|Modifier|false|false||openingnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C1549543;C0030193;C0332803|incisionnull|Increased pain|Finding|false|false||increased painnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Administration Method - Pain|Finding|false|false|C2338258|pain
null|Pain|Finding|false|false|C2338258|painnull|null|Attribute|false|false||painnull|Contusions|Disorder|false|false||bruisingnull|reported bruising (history)|Finding|false|false||bruisingnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false|C1123023;C4520765|infectionnull|Infection|Finding|false|false||infectionnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C0009450;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C0009450;C1546781;C0444099|skinnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Increased pain|Finding|false|false||increased painnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Rapid|Modifier|false|false||quicknull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||return tonull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Usual|Modifier|false|false||usualnull|Life|Finding|false|false||lifenull|Laser-Induced Fluorescence Endoscopy|Procedure|false|false||lifenull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Foley catheter|Device|false|false||Foley catheternull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0872388|bladdernull|Urology|Title|false|false||urologynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|Appointments|Event|false|false||appointmentnull|Urology|Title|false|false||Urologynull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|MDF AttributeType - Number|Finding|false|false||numbernull|Count of entities|LabModifier|false|false||number
null|Numbers|LabModifier|false|false||numbernull|Appointments|Event|false|false||appointmentnull|Attempt|Event|false|false||attemptnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Exhausted|Finding|false|false||Emptynull|Empty (qualifier)|Modifier|false|false||Emptynull|Bag Data Type|Finding|false|false||bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|Nursing Staff|Subject|false|false||nursing staffnull|Breast Feeding|Finding|false|false||nursingnull|RNAx nursing therapy actions|Procedure|false|false||nursingnull|Discipline of Nursing|Title|false|false||nursingnull|Encounter Special Courtesy - staff|Finding|false|false||staffnull|Staff|Subject|false|false||staffnull|On Staff|Modifier|false|false||staffnull|Leg bag|Device|false|false||leg bagnull|Leg|Anatomy|false|false|C1552710|leg
null|Lower Extremity|Anatomy|false|false|C1552710|legnull|Bag Data Type|Finding|false|false|C1140621;C0023216|bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Tripping|Phenomenon|false|false||tripsnull|Smaller|Modifier|false|false||smallernull|Small|LabModifier|false|false||smallernull|Bag Data Type|Finding|false|false||bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|null|Device|false|false||strapsnull|Leg|Anatomy|false|false|C1553498;C1549632;C1548341|leg
null|Lower Extremity|Anatomy|false|false|C1553498;C1549632;C1548341|legnull|Visit User Code - Home|Finding|false|false|C1140621;C0023216|home
null|Address type - Home|Finding|false|false|C1140621;C0023216|homenull|home health encounter|Procedure|false|false|C1140621;C0023216|homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Smaller|Modifier|false|false||smallernull|Small|LabModifier|false|false||smallernull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Bag Data Type|Finding|false|false||bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|More|LabModifier|false|false||morenull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Persons|Subject|false|false||peoplenull|Greater|LabModifier|false|false||larger
null|Large|LabModifier|false|false||largernull|BAD protein, human|Drug|false|false||bad
null|BAD protein, human|Drug|false|false||badnull|Brachial Amyotrophic Diplegia|Disorder|false|false||badnull|BAD gene|Finding|false|false||badnull|Banda language|Entity|false|false||badnull|Bad|Modifier|false|false||badnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions