 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|244,255|false|false|false|||Varenicline
Event|Event|Allergies|258,267|false|false|false|||Attending
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Disorder|Disease or Syndrome|Chief Complaint|293,299|false|false|false|C0002871|Anemia|Anemia
Event|Event|Chief Complaint|293,299|false|false|false|||Anemia
Event|Event|Chief Complaint|301,307|false|false|false|||Melena
Finding|Pathologic Function|Chief Complaint|301,307|false|false|false|C0025222|Melena|Melena
Event|Event|Chief Complaint|309,312|false|false|false|||SOB
Finding|Sign or Symptom|Chief Complaint|309,312|false|false|false|C0013404|Dyspnea|SOB
Finding|Classification|Chief Complaint|315,320|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|321,329|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|333,351|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|342,351|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|342,351|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|342,351|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|342,351|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|342,351|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|359,368|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|Chief Complaint|359,368|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|History of Present Illness|423,430|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|423,430|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|423,430|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|423,430|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|423,433|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|434,438|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|History of Present Illness|434,438|false|false|false|||Afib
Lab|Laboratory or Test Result|History of Present Illness|434,438|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Drug|Organic Chemical|History of Present Illness|442,449|false|false|false|C3159309|Xarelto|Xarelto
Drug|Pharmacologic Substance|History of Present Illness|442,449|false|false|false|C3159309|Xarelto|Xarelto
Disorder|Disease or Syndrome|History of Present Illness|451,455|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|451,455|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|451,455|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|451,455|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|457,460|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|457,460|false|false|false|||HTN
Anatomy|Anatomical Structure|History of Present Illness|462,465|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|History of Present Illness|462,465|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|History of Present Illness|462,465|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|History of Present Illness|462,465|false|false|false|C2347441|Pad Dosage Form|PAD
Event|Event|History of Present Illness|462,465|false|false|false|||PAD
Finding|Gene or Genome|History of Present Illness|462,465|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|462,465|false|false|false|C3814046|PAD Regimen|PAD
Event|Event|History of Present Illness|471,479|false|false|false|||presents
Finding|Finding|History of Present Illness|484,492|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|History of Present Illness|484,492|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Event|History of Present Illness|493,497|false|false|false|||labs
Lab|Laboratory or Test Result|History of Present Illness|493,497|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|History of Present Illness|503,508|false|false|false|||noted
Event|Event|History of Present Illness|515,520|false|false|false|||tarry
Finding|Finding|History of Present Illness|515,520|false|false|false|C4069282|Tarry|tarry
Finding|Body Substance|History of Present Illness|522,527|false|false|false|C0015733|Feces|stool
Event|Event|History of Present Illness|540,549|false|false|false|||presented
Disorder|Disease or Syndrome|History of Present Illness|553,556|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|553,556|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|553,556|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|553,556|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|553,556|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|553,556|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|553,556|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|553,556|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|553,556|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|553,556|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|553,556|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|580,585|false|false|false|||noted
Drug|Biomedical or Dental Material|History of Present Illness|623,631|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|623,631|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|632,635|false|false|false|||Hct
Procedure|Laboratory Procedure|History of Present Illness|632,635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|632,635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Finding|Finding|History of Present Illness|679,685|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Finding|Gene or Genome|History of Present Illness|679,685|false|false|false|C0423899;C1414153;C3539536|ARID1B wt Allele;ARID3A gene;Above average intellect|bright
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|679,689|false|false|false|C1096868|DC Red No. 8|bright red
Drug|Organic Chemical|History of Present Illness|679,689|false|false|false|C1096868|DC Red No. 8|bright red
Finding|Finding|History of Present Illness|679,689|false|false|false|C1272329|Bright red color (finding)|bright red
Finding|Finding|History of Present Illness|686,689|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|History of Present Illness|686,689|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Disorder|Disease or Syndrome|History of Present Illness|690,695|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|690,695|false|false|false|||blood
Finding|Body Substance|History of Present Illness|690,695|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|History of Present Illness|714,722|false|false|false|||believes
Disorder|Disease or Syndrome|History of Present Illness|732,743|false|false|false|C0019112|Hemorrhoids|hemorrhoids
Event|Event|History of Present Illness|732,743|false|false|false|||hemorrhoids
Disorder|Disease or Syndrome|History of Present Illness|745,748|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|745,748|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|745,748|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|745,748|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|745,748|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|745,748|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|745,748|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|745,748|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|745,748|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|745,748|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|745,748|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|749,755|false|false|false|||called
Event|Event|History of Present Illness|763,769|false|false|false|||agreed
Event|Event|History of Present Illness|773,777|false|false|false|||come
Event|Event|History of Present Illness|794,805|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|History of Present Illness|794,805|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|History of Present Illness|794,805|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|History of Present Illness|818,824|false|false|false|||showed
Disorder|Anatomical Abnormality|History of Present Illness|834,839|false|false|false|C0032584|polyps|polyp
Event|Event|History of Present Illness|834,839|false|false|false|||polyp
Disorder|Disease or Syndrome|History of Present Illness|842,862|false|false|false|C0265034|Internal hemorrhoids|internal hemorrhoids
Disorder|Disease or Syndrome|History of Present Illness|851,862|false|false|false|C0019112|Hemorrhoids|hemorrhoids
Event|Event|History of Present Illness|851,862|false|false|false|||hemorrhoids
Disorder|Disease or Syndrome|History of Present Illness|868,882|false|false|false|C1510475|Diverticulosis|diverticulosis
Event|Event|History of Present Illness|868,882|false|false|false|||diverticulosis
Event|Event|History of Present Illness|893,895|false|false|false|||BM
Event|Event|History of Present Illness|946,955|false|false|false|||complains
Event|Event|History of Present Illness|959,968|false|false|false|||increased
Finding|Finding|History of Present Illness|959,968|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|History of Present Illness|959,968|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Sign or Symptom|History of Present Illness|970,980|false|false|false|C0239313|exercise induced|exertional
Finding|Sign or Symptom|History of Present Illness|970,988|false|false|false|C0743838|Exertional fatigue|exertional fatigue
Event|Event|History of Present Illness|981,988|false|false|false|||fatigue
Finding|Sign or Symptom|History of Present Illness|981,988|false|false|false|C0015672|Fatigue|fatigue
Event|Event|History of Present Illness|1002,1009|false|false|false|||feeling
Event|Event|History of Present Illness|1015,1018|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|1015,1018|false|false|false|C0013404|Dyspnea|SOB
Drug|Biomedical or Dental Material|History of Present Illness|1029,1037|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1029,1037|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1029,1037|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|1071,1078|false|false|false|||noticed
Event|Event|History of Present Illness|1083,1090|false|false|false|||becomes
Finding|Sign or Symptom|History of Present Illness|1105,1118|false|false|false|C0848168|out (of) breath|out of breath
Finding|Body Substance|History of Present Illness|1112,1118|false|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|1120,1127|false|false|false|||walking
Finding|Daily or Recreational Activity|History of Present Illness|1120,1127|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|History of Present Illness|1120,1127|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|History of Present Illness|1120,1127|false|false|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|History of Present Illness|1131,1139|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Individual Behavior|History of Present Illness|1131,1139|false|false|false|C0561942;C2362653;C2584300|Climbing;Does climb;climbing (history)|climbing
Finding|Daily or Recreational Activity|History of Present Illness|1131,1146|false|false|false|C1290942|Climbing stairs|climbing stairs
Event|Event|History of Present Illness|1140,1146|false|false|false|||stairs
Finding|Finding|History of Present Illness|1140,1146|false|false|false|C4300351|Prior functioning.stairs|stairs
Event|Event|History of Present Illness|1154,1161|false|false|false|||becomes
Event|Event|History of Present Illness|1162,1165|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|1162,1165|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|1174,1180|false|false|false|||stairs
Finding|Finding|History of Present Illness|1174,1180|false|false|false|C4300351|Prior functioning.stairs|stairs
Drug|Biomedical or Dental Material|History of Present Illness|1196,1201|false|false|false|C1706085|Block Dosage Form|block
Event|Event|History of Present Illness|1196,1201|false|false|false|||block
Finding|Body Substance|History of Present Illness|1196,1201|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|History of Present Illness|1196,1201|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|History of Present Illness|1196,1201|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Event|Event|History of Present Illness|1203,1212|false|false|false|||requiring
Event|Event|History of Present Illness|1221,1225|false|false|false|||stop
Disorder|Disease or Syndrome|History of Present Illness|1234,1239|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|1240,1243|false|false|false|||use
Drug|Organic Chemical|History of Present Illness|1244,1253|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|History of Present Illness|1244,1253|false|false|false|C0001927|albuterol|albuterol
Event|Event|History of Present Illness|1254,1261|false|false|false|||inhaler
Finding|Functional Concept|History of Present Illness|1254,1261|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Event|Event|History of Present Illness|1267,1271|false|false|false|||used
Event|Event|History of Present Illness|1275,1278|false|false|false|||use
Event|Event|History of Present Illness|1289,1292|false|false|false|||use
Event|Event|History of Present Illness|1297,1304|false|false|false|||inhaler
Finding|Functional Concept|History of Present Illness|1297,1304|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Disorder|Disease or Syndrome|History of Present Illness|1309,1314|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|1309,1314|false|false|false|||times
Finding|Idea or Concept|History of Present Illness|1319,1322|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1319,1322|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|1332,1336|false|false|false|||uses
Disorder|Disease or Syndrome|History of Present Illness|1351,1356|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|History of Present Illness|1359,1362|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1359,1362|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Pharmacologic Substance|History of Present Illness|1367,1377|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|History of Present Illness|1367,1377|false|false|false|||nebulizers
Finding|Idea or Concept|History of Present Illness|1386,1389|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1386,1389|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|1397,1403|true|false|false|||denies
Event|Event|History of Present Illness|1408,1414|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1408,1414|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1416,1422|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1416,1422|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|1424,1430|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|1424,1430|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1424,1430|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1431,1436|true|false|false|||vomit
Finding|Body Substance|History of Present Illness|1431,1436|true|false|false|C0042963;C0042965|Vomiting;Vomitus|vomit
Finding|Sign or Symptom|History of Present Illness|1431,1436|true|false|false|C0042963;C0042965|Vomiting;Vomitus|vomit
Event|Event|History of Present Illness|1438,1446|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1438,1446|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1438,1446|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|1448,1455|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|1448,1455|true|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|History of Present Illness|1458,1462|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|History of Present Illness|1458,1462|false|false|false|||rash
Finding|Pathologic Function|History of Present Illness|1458,1462|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|1458,1462|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Functional Concept|History of Present Illness|1464,1477|false|false|false|C1283932|Unintentional|unintentional
Finding|Finding|History of Present Illness|1464,1489|false|false|false|C2363736|Unintentional weight loss|unintentional weight loss
Attribute|Clinical Attribute|History of Present Illness|1478,1484|false|false|false|C0944911||weight
Event|Event|History of Present Illness|1478,1484|false|false|false|||weight
Finding|Finding|History of Present Illness|1478,1484|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1478,1484|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1478,1484|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|1478,1489|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|1478,1489|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|1485,1489|false|false|false|||loss
Finding|Finding|History of Present Illness|1485,1489|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Idea or Concept|History of Present Illness|1508,1515|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1516,1522|false|false|false|||vitals
Lab|Laboratory or Test Result|History of Present Illness|1550,1554|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|1555,1566|false|false|false|||significant
Finding|Idea or Concept|History of Present Illness|1555,1566|false|false|false|C0750502|Significant|significant
Anatomy|Cell|History of Present Illness|1572,1575|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1572,1575|false|false|false|||WBC
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1580,1583|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|History of Present Illness|1580,1583|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|History of Present Illness|1580,1583|false|false|false|||HGB
Finding|Gene or Genome|History of Present Illness|1580,1583|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|History of Present Illness|1580,1583|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|History of Present Illness|1588,1591|false|false|false|||HCT
Procedure|Laboratory Procedure|History of Present Illness|1588,1591|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1588,1591|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Drug|Biomedical or Dental Material|History of Present Illness|1603,1611|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1603,1611|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1603,1611|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Virus|History of Present Illness|1635,1638|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|History of Present Illness|1635,1638|false|false|false|||MCV
Lab|Laboratory or Test Result|History of Present Illness|1635,1638|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|History of Present Illness|1635,1638|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1635,1638|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Event|Event|History of Present Illness|1639,1642|false|false|false|||PLT
Procedure|Laboratory Procedure|History of Present Illness|1639,1642|false|false|false|C0201617|Primed lymphocyte test|PLT
Attribute|Clinical Attribute|History of Present Illness|1657,1660|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1657,1660|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1657,1660|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1657,1660|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Disorder|Neoplastic Process|History of Present Illness|1665,1668|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|History of Present Illness|1665,1668|false|false|false|||PTT
Procedure|Laboratory Procedure|History of Present Illness|1665,1668|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Functional Concept|History of Present Illness|1674,1678|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|History of Present Illness|1674,1678|false|false|false|C0201682|Chemical procedure|Chem
Procedure|Laboratory Procedure|History of Present Illness|1674,1680|false|false|false|C2237045|Basic metabolic panel|Chem 7
Event|Event|History of Present Illness|1685,1691|false|false|false|||normal
Drug|Organic Chemical|History of Present Illness|1707,1716|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|History of Present Illness|1707,1716|false|false|false|C0001927|albuterol|albuterol
Drug|Biomedical or Dental Material|History of Present Illness|1717,1721|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|History of Present Illness|1717,1721|false|false|false|||nebs
Event|Event|History of Present Illness|1726,1733|false|false|false|||started
Finding|Finding|History of Present Illness|1734,1739|false|false|false|C3714655|On IV|on IV
Drug|Inorganic Chemical|History of Present Illness|1747,1753|false|false|false|C0036082|Saline Solution|saline
Drug|Pharmacologic Substance|History of Present Illness|1747,1753|false|false|false|C0036082|Saline Solution|saline
Event|Event|History of Present Illness|1747,1753|false|false|false|||saline
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1747,1753|false|false|false|C0450082|Saline method|saline
Event|Event|History of Present Illness|1759,1767|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1759,1767|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1759,1767|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1759,1767|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|History of Present Illness|1769,1775|false|false|false|||vitals
Event|Activity|History of Present Illness|1830,1837|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|1830,1837|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1830,1837|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|1845,1850|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|1851,1858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1851,1858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1851,1858|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1863,1869|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1863,1869|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Mental Process|History of Present Illness|1874,1889|false|false|false|C0018592|Happiness|in good spirits
Finding|Idea or Concept|History of Present Illness|1877,1881|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Food|History of Present Illness|1882,1889|false|false|false|C0301611|distilled alcoholic beverage|spirits
Event|Event|History of Present Illness|1882,1889|false|false|false|||spirits
Event|Event|History of Present Illness|1896,1901|false|false|false|||notes
Disorder|Disease or Syndrome|History of Present Illness|1920,1925|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|1920,1925|false|false|false|||blood
Finding|Body Substance|History of Present Illness|1920,1925|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|History of Present Illness|1920,1936|false|false|false|C0267596|Rectal hemorrhage|blood per rectum
Finding|Functional Concept|History of Present Illness|1926,1936|false|false|false|C1527425;C4048189|Per rectum;Rectal Route of Administration|per rectum
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1930,1936|false|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|rectum
Disorder|Disease or Syndrome|History of Present Illness|1930,1936|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Disorder|Neoplastic Process|History of Present Illness|1930,1936|false|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|rectum
Event|Event|History of Present Illness|1930,1936|false|false|false|||rectum
Procedure|Health Care Activity|History of Present Illness|1930,1936|false|false|false|C0869814|Procedure on rectum|rectum
Event|Event|History of Present Illness|1944,1953|false|false|false|||underwear
Disorder|Disease or Syndrome|Past Medical History|1982,1988|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|Past Medical History|1982,1988|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1989,1993|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1989,1993|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1989,1993|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1989,1993|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Hazardous or Poisonous Substance|Past Medical History|1994,2001|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|Past Medical History|1994,2001|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|Past Medical History|1994,2001|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|Past Medical History|1994,2001|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Attribute|Clinical Attribute|Past Medical History|1994,2005|false|false|false|C4522050||Tobacco use
Finding|Finding|Past Medical History|1994,2005|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Finding|Individual Behavior|Past Medical History|1994,2005|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Event|Event|Past Medical History|2002,2005|false|false|false|||use
Finding|Functional Concept|Past Medical History|2002,2005|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Past Medical History|2002,2005|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Disorder|Disease or Syndrome|Past Medical History|2007,2034|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|Peripheral Arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2018,2026|false|false|false|C0003842|Arteries|Arterial
Disorder|Disease or Syndrome|Past Medical History|2018,2034|false|false|false|C0852949|Arteriopathic disease|Arterial disease
Disorder|Disease or Syndrome|Past Medical History|2027,2034|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|2027,2034|false|false|false|||disease
Finding|Functional Concept|Past Medical History|2047,2053|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Past Medical History|2047,2053|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2054,2059|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2054,2068|false|false|false|C0850459|iliac stents|iliac stenting
Event|Event|Past Medical History|2060,2068|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2060,2068|false|false|false|C2348535|Stenting|stenting
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2070,2076|false|false|false|C0018792|Heart Atrium|ATRIAL
Disorder|Disease or Syndrome|Past Medical History|2070,2088|false|false|false|C0546959|Atrial tachycardia|ATRIAL TACHYCARDIA
Finding|Finding|Past Medical History|2070,2088|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|ATRIAL TACHYCARDIA
Event|Event|Past Medical History|2077,2088|false|false|false|||TACHYCARDIA
Finding|Finding|Past Medical History|2077,2088|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|TACHYCARDIA
Finding|Finding|Past Medical History|2090,2098|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|2090,2109|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|2099,2104|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|2099,2104|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|2099,2109|false|true|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|2099,2109|false|true|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|2105,2109|false|true|false|C2598155||PAIN
Event|Event|Past Medical History|2105,2109|false|false|false|||PAIN
Finding|Functional Concept|Past Medical History|2105,2109|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|2105,2109|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Past Medical History|2112,2120|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|2112,2132|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|Past Medical History|2121,2132|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|Past Medical History|2121,2132|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|Past Medical History|2134,2142|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|2134,2154|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|Past Medical History|2143,2154|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|Past Medical History|2143,2154|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2156,2164|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2156,2171|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2165,2171|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|2165,2171|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|2173,2180|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2173,2180|false|false|false|||DISEASE
Event|Event|Past Medical History|2183,2191|false|false|false|||HEADACHE
Finding|Sign or Symptom|Past Medical History|2183,2191|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2193,2196|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2193,2196|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|2193,2196|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|2193,2196|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|2193,2196|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|2193,2196|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2193,2196|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2193,2208|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|2197,2208|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|2197,2208|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|2197,2208|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2197,2208|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|Past Medical History|2210,2224|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|2210,2224|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|2210,2224|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Past Medical History|2226,2238|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|2226,2238|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|2241,2255|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Disorder|Disease or Syndrome|Past Medical History|2257,2263|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|Past Medical History|2257,2270|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|Past Medical History|2257,2270|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|Past Medical History|2264,2270|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|Past Medical History|2264,2270|false|false|false|||ZOSTER
Drug|Hazardous or Poisonous Substance|Past Medical History|2272,2279|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Past Medical History|2272,2279|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Past Medical History|2272,2279|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Past Medical History|2272,2279|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2272,2285|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2280,2285|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Past Medical History|2280,2285|false|false|false|||ABUSE
Event|Event|Past Medical History|2280,2285|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Past Medical History|2280,2285|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2287,2293|false|false|false|C0018792|Heart Atrium|ATRIAL
Disorder|Disease or Syndrome|Past Medical History|2295,2307|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|2295,2307|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2310,2317|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|Past Medical History|2310,2317|false|false|false|||ANXIETY
Finding|Sign or Symptom|Past Medical History|2310,2317|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Past Medical History|2318,2334|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Past Medical History|2318,2343|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Event|Event|Past Medical History|2335,2343|false|false|false|||BLEEDING
Finding|Pathologic Function|Past Medical History|2335,2343|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Past Medical History|2345,2359|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|2345,2359|false|false|false|||OSTEOARTHRITIS
Finding|Functional Concept|Past Medical History|2362,2377|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|Past Medical History|2362,2400|false|true|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|Past Medical History|2378,2392|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|Past Medical History|2378,2400|false|true|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|2393,2400|false|true|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2393,2400|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|2393,2421|false|false|false|C0085096|Peripheral Vascular Diseases|DISEASE, PERIPHERAL VASCULAR
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2413,2421|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|Past Medical History|2423,2430|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|2423,2430|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|2432,2440|false|false|false|C0086543|Cataract|CATARACT
Event|Event|Past Medical History|2432,2440|false|false|false|||CATARACT
Finding|Finding|Past Medical History|2432,2440|false|false|false|C1690964|cataract on exam (physical finding)|CATARACT
Finding|Finding|Past Medical History|2432,2448|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Finding|Intellectual Product|Past Medical History|2432,2448|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2432,2448|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|CATARACT SURGERY
Event|Event|Past Medical History|2441,2448|false|false|false|||SURGERY
Finding|Finding|Past Medical History|2441,2448|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Past Medical History|2441,2448|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Past Medical History|2441,2448|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2441,2448|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Finding|Past Medical History|2455,2462|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Past Medical History|2455,2462|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Past Medical History|2455,2462|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2455,2462|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Finding|Functional Concept|Past Medical History|2476,2482|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Finding|Intellectual Product|Past Medical History|2476,2482|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2476,2495|false|false|false|C1261084|Common iliac artery structure|COMMON ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2483,2488|false|false|false|C0020889|Bone structure of ilium|ILIAC
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2483,2495|false|false|false|C0020887|Structure of iliac artery|ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2489,2495|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|2489,2495|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Event|Event|Past Medical History|2496,2504|false|false|false|||STENTING
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2496,2504|false|false|false|C2348535|Stenting|STENTING
Event|Event|Past Medical History|2511,2523|false|false|false|||BUNIONECTOMY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2511,2523|false|false|false|C1542057|Silver bunionectomy|BUNIONECTOMY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2526,2529|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2526,2529|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|2526,2529|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|2526,2529|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|2526,2529|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|2526,2529|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2526,2529|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2526,2541|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|2530,2541|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|2530,2541|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|2530,2541|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2530,2541|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2550,2558|false|false|false|C3841297|Cesarean|CESAREAN
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2550,2566|false|false|false|C0007876|Cesarean section|CESAREAN SECTION
Drug|Substance|Past Medical History|2559,2566|false|false|false|C1522472|section sample|SECTION
Event|Event|Past Medical History|2559,2566|false|false|false|||SECTION
Finding|Intellectual Product|Past Medical History|2559,2566|false|false|false|C1551341;C1552858|Act Class - Section;Html Link Type - section|SECTION
Procedure|Laboratory Procedure|Past Medical History|2559,2566|false|false|false|C0700320|Sectioning technique|SECTION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2569,2577|false|false|false|C0017067|Ganglia|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2569,2577|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2569,2582|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION CYST
Disorder|Anatomical Abnormality|Past Medical History|2578,2582|false|false|false|C0010709|Cyst|CYST
Event|Event|Past Medical History|2578,2582|false|false|false|||CYST
Finding|Body Substance|Past Medical History|2578,2582|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Intellectual Product|Past Medical History|2578,2582|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Idea or Concept|Family Medical History|2621,2627|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2634,2637|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|2634,2637|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|2640,2646|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2640,2646|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|2657,2664|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2657,2664|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2657,2664|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2672,2679|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2672,2679|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2672,2679|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2688,2696|false|false|false|||Physical
Finding|Finding|Family Medical History|2688,2696|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|2688,2696|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|2688,2696|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|2702,2711|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|Family Medical History|2712,2720|false|false|false|||PHYSICAL
Finding|Finding|Family Medical History|2712,2720|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|2712,2720|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|2712,2720|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|2712,2725|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|2712,2725|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|Family Medical History|2721,2725|false|false|false|||EXAM
Finding|Functional Concept|Family Medical History|2721,2725|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|2721,2725|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|Family Medical History|2778,2785|false|false|false|||GENERAL
Finding|Classification|Family Medical History|2778,2785|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|2778,2785|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|Family Medical History|2787,2791|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|Family Medical History|2792,2801|false|false|false|||nourished
Finding|Finding|Family Medical History|2803,2807|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|2808,2817|false|false|false|||appearing
Event|Event|Family Medical History|2829,2836|false|false|false|||sitting
Disorder|Disease or Syndrome|Family Medical History|2844,2847|true|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|Family Medical History|2844,2847|true|false|false|||bed
Finding|Intellectual Product|Family Medical History|2844,2847|true|false|false|C2346952|Bachelor of Education|bed
Attribute|Clinical Attribute|Family Medical History|2848,2853|true|false|false|C5890168||Alert
Drug|Organic Chemical|Family Medical History|2848,2853|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Family Medical History|2848,2853|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Family Medical History|2848,2853|true|false|false|||Alert
Finding|Finding|Family Medical History|2848,2853|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Family Medical History|2848,2853|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Family Medical History|2848,2853|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Family Medical History|2855,2863|true|false|false|||oriented
Finding|Intellectual Product|Family Medical History|2868,2873|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Family Medical History|2874,2882|true|false|false|||distress
Finding|Finding|Family Medical History|2874,2882|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|2874,2882|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|2885,2890|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2892,2898|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|2892,2898|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|2892,2898|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|2892,2898|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|2899,2908|false|false|false|||anicteric
Finding|Finding|Family Medical History|2899,2908|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2910,2913|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|2910,2913|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|2915,2925|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|2926,2931|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|2926,2931|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|2934,2938|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Family Medical History|2934,2938|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Family Medical History|2934,2938|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|Family Medical History|2940,2946|true|false|false|||supple
Finding|Functional Concept|Family Medical History|2940,2946|true|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|2948,2951|true|false|false|||JVP
Finding|Finding|Family Medical History|2948,2951|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|2956,2964|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2969,2972|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|2969,2972|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|2969,2972|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|2969,2972|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2975,2980|true|false|false|C0024109|Lung|LUNGS
Event|Event|Family Medical History|2982,2987|false|false|false|||Clear
Finding|Idea or Concept|Family Medical History|2982,2987|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Family Medical History|2991,3003|false|false|false|||auscultation
Procedure|Diagnostic Procedure|Family Medical History|2991,3003|false|false|false|C0004339|Auscultation|auscultation
Drug|Inorganic Chemical|Family Medical History|3033,3036|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|3033,3036|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|3033,3036|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Family Medical History|3033,3036|false|false|false|||air
Finding|Finding|Family Medical History|3033,3036|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|3033,3036|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|3033,3036|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Family Medical History|3038,3046|false|false|false|||movement
Finding|Organism Function|Family Medical History|3038,3046|false|false|false|C0026649|Movement|movement
Event|Event|Family Medical History|3054,3061|true|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|3054,3061|true|false|false|C0043144|Wheezing|wheezes
Event|Event|Family Medical History|3063,3068|true|false|false|||rales
Finding|Finding|Family Medical History|3063,3068|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|Family Medical History|3070,3077|true|false|false|||rhonchi
Finding|Finding|Family Medical History|3070,3077|true|false|false|C0035508|Rhonchi|rhonchi
Event|Activity|Family Medical History|3106,3110|false|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|3106,3110|false|false|false|||rate
Finding|Idea or Concept|Family Medical History|3106,3110|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|3115,3121|false|false|false|||rhythm
Finding|Finding|Family Medical History|3115,3121|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|3115,3121|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Organ or Tissue Function|Family Medical History|3142,3150|true|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|3142,3157|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|3151,3157|true|false|false|||murmur
Finding|Finding|Family Medical History|3151,3157|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|3158,3163|true|false|false|||heard
Event|Event|Family Medical History|3181,3185|true|false|false|||rubs
Finding|Finding|Family Medical History|3181,3185|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|3189,3196|true|false|false|||gallops
Anatomy|Body Location or Region|Family Medical History|3199,3202|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|Family Medical History|3199,3202|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|Family Medical History|3199,3202|true|false|false|||ABD
Disorder|Disease or Syndrome|Family Medical History|3204,3208|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|3204,3208|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3237,3242|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|3237,3249|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|3243,3249|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3243,3249|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3250,3257|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|3250,3257|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|Family Medical History|3263,3281|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|Family Medical History|3271,3281|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|3271,3281|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|3271,3281|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Family Medical History|3285,3293|true|false|false|||guarding
Finding|Finding|Family Medical History|3285,3293|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|Family Medical History|3298,3310|true|false|false|||organomegaly
Finding|Finding|Family Medical History|3298,3310|true|false|false|C4054315|Organomegaly|organomegaly
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3312,3318|true|false|false|C0034896;C4482211|Pelvis>Rectum;Rectum|Rectum
Disorder|Disease or Syndrome|Family Medical History|3312,3318|true|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|Rectum
Disorder|Neoplastic Process|Family Medical History|3312,3318|true|false|false|C0034882;C0154062;C0496867;C0496908|Benign neoplasm of rectum;Carcinoma in situ of rectum;Neoplasm of uncertain or unknown behavior of rectum;Rectal Diseases|Rectum
Event|Event|Family Medical History|3312,3318|true|false|false|||Rectum
Procedure|Health Care Activity|Family Medical History|3312,3318|true|false|false|C0869814|Procedure on rectum|Rectum
Disorder|Disease or Syndrome|Family Medical History|3331,3342|true|false|false|C0019112|Hemorrhoids|hemorrhoids
Event|Event|Family Medical History|3331,3342|true|false|false|||hemorrhoids
Disorder|Congenital Abnormality|Family Medical History|3345,3348|true|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|Family Medical History|3345,3348|true|false|false|||EXT
Finding|Gene or Genome|Family Medical History|3345,3348|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|Family Medical History|3350,3354|false|false|false|||Warm
Finding|Finding|Family Medical History|3350,3354|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3350,3354|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|3356,3360|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3361,3369|true|false|false|||perfused
Drug|Food|Family Medical History|3374,3380|true|false|false|C5890763||pulses
Event|Event|Family Medical History|3374,3380|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|3374,3380|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|3374,3380|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|3385,3393|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|3385,3393|true|false|false|||clubbing
Event|Event|Family Medical History|3395,3403|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|3395,3403|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|3408,3413|true|false|false|C1717255||edema
Event|Event|Family Medical History|3408,3413|true|false|false|||edema
Finding|Pathologic Function|Family Medical History|3408,3413|true|false|false|C0013604|Edema|edema
Anatomy|Body System|Family Medical History|3416,3420|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|Family Medical History|3416,3420|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|Family Medical History|3416,3420|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|Family Medical History|3416,3420|false|false|false|||SKIN
Finding|Body Substance|Family Medical History|3416,3420|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|Family Medical History|3416,3420|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|Family Medical History|3422,3427|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|3422,3427|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Family Medical History|3444,3452|true|false|false|||deficits
Finding|Body Substance|Family Medical History|3455,3464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|3455,3464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|3455,3464|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|3455,3464|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|Family Medical History|3465,3473|false|false|false|||PHYSICAL
Finding|Finding|Family Medical History|3465,3473|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|3465,3473|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|3465,3473|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|3465,3478|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|3465,3478|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|Family Medical History|3474,3478|false|false|false|||EXAM
Finding|Functional Concept|Family Medical History|3474,3478|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|3474,3478|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|Family Medical History|3541,3548|false|false|false|||GENERAL
Finding|Classification|Family Medical History|3541,3548|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|3541,3548|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|Family Medical History|3550,3554|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|Family Medical History|3555,3564|false|false|false|||nourished
Finding|Finding|Family Medical History|3566,3570|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3571,3580|false|false|false|||appearing
Event|Event|Family Medical History|3582,3589|false|false|false|||sitting
Disorder|Disease or Syndrome|Family Medical History|3596,3599|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|Family Medical History|3596,3599|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|Family Medical History|3601,3604|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|3601,3604|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|3601,3604|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|3601,3604|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|3601,3604|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|3601,3604|false|false|false|||NAD
Finding|Finding|Family Medical History|3601,3604|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|3605,3610|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3612,3618|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|3612,3618|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|Family Medical History|3612,3618|false|false|false|||Sclera
Procedure|Health Care Activity|Family Medical History|3612,3618|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|Family Medical History|3619,3628|false|false|false|||anicteric
Finding|Finding|Family Medical History|3619,3628|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3630,3633|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|3630,3633|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|Family Medical History|3635,3645|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|Family Medical History|3646,3651|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|3646,3651|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|Family Medical History|3654,3658|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Family Medical History|3654,3658|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Family Medical History|3654,3658|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|Family Medical History|3660,3666|true|false|false|||supple
Finding|Functional Concept|Family Medical History|3660,3666|true|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|3668,3671|true|false|false|||JVP
Finding|Finding|Family Medical History|3668,3671|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|Family Medical History|3676,3684|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3689,3692|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|3689,3692|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|3689,3692|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|3689,3692|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3695,3700|true|false|false|C0024109|Lung|LUNGS
Event|Event|Family Medical History|3712,3719|false|false|false|||wheezes
Finding|Sign or Symptom|Family Medical History|3712,3719|false|false|false|C0043144|Wheezing|wheezes
Attribute|Clinical Attribute|Family Medical History|3739,3743|true|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|Family Medical History|3739,3743|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|Family Medical History|3744,3752|true|false|false|||distress
Finding|Finding|Family Medical History|3744,3752|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|3744,3752|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Activity|Family Medical History|3780,3784|false|false|false|C0871208|Rating (action)|rate
Event|Event|Family Medical History|3780,3784|false|false|false|||rate
Finding|Idea or Concept|Family Medical History|3780,3784|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Family Medical History|3789,3795|false|false|false|||rhythm
Finding|Finding|Family Medical History|3789,3795|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|3789,3795|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Organ or Tissue Function|Family Medical History|3816,3824|true|false|false|C0039155|Systole|systolic
Finding|Finding|Family Medical History|3816,3831|true|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|Family Medical History|3825,3831|true|false|false|||murmur
Finding|Finding|Family Medical History|3825,3831|true|false|false|C0018808|Heart murmur|murmur
Event|Event|Family Medical History|3832,3837|true|false|false|||heard
Event|Event|Family Medical History|3855,3859|true|false|false|||rubs
Finding|Finding|Family Medical History|3855,3859|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|3863,3870|true|false|false|||gallops
Anatomy|Body Location or Region|Family Medical History|3871,3874|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|Family Medical History|3871,3874|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|Family Medical History|3871,3874|true|false|false|||ABD
Disorder|Disease or Syndrome|Family Medical History|3876,3880|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|3876,3880|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3909,3914|true|false|false|C0021853|Intestines|bowel
Finding|Finding|Family Medical History|3909,3921|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|Family Medical History|3915,3921|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3915,3921|true|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3922,3929|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|3922,3929|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|Family Medical History|3935,3953|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|Family Medical History|3943,3953|true|false|false|||tenderness
Finding|Mental Process|Family Medical History|3943,3953|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|3943,3953|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Family Medical History|3957,3965|true|false|false|||guarding
Finding|Finding|Family Medical History|3957,3965|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|Family Medical History|3970,3982|true|false|false|||organomegaly
Finding|Finding|Family Medical History|3970,3982|true|false|false|C4054315|Organomegaly|organomegaly
Disorder|Congenital Abnormality|Family Medical History|3983,3986|true|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|Family Medical History|3983,3986|true|false|false|||EXT
Finding|Gene or Genome|Family Medical History|3983,3986|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|Family Medical History|3988,3992|false|false|false|||Warm
Finding|Finding|Family Medical History|3988,3992|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3988,3992|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|3994,3998|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3999,4007|true|false|false|||perfused
Drug|Food|Family Medical History|4012,4018|true|false|false|C5890763||pulses
Event|Event|Family Medical History|4012,4018|true|false|false|||pulses
Finding|Physiologic Function|Family Medical History|4012,4018|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Family Medical History|4012,4018|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|Family Medical History|4023,4031|true|false|false|C0149651|Clubbing|clubbing
Event|Event|Family Medical History|4023,4031|true|false|false|||clubbing
Event|Event|Family Medical History|4033,4041|true|false|false|||cyanosis
Finding|Sign or Symptom|Family Medical History|4033,4041|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|Family Medical History|4046,4051|true|false|false|C1717255||edema
Event|Event|Family Medical History|4046,4051|true|false|false|||edema
Finding|Pathologic Function|Family Medical History|4046,4051|true|false|false|C0013604|Edema|edema
Anatomy|Body System|Family Medical History|4054,4058|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|Family Medical History|4054,4058|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|Family Medical History|4054,4058|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|Family Medical History|4054,4058|false|false|false|||SKIN
Finding|Body Substance|Family Medical History|4054,4058|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|Family Medical History|4054,4058|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|Family Medical History|4060,4065|false|false|false|||clear
Finding|Idea or Concept|Family Medical History|4060,4065|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|Family Medical History|4082,4090|true|false|false|||deficits
Procedure|Health Care Activity|Family Medical History|4114,4123|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|Family Medical History|4124,4128|false|false|false|||LABS
Lab|Laboratory or Test Result|Family Medical History|4124,4128|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|4159,4164|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4159,4164|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4159,4164|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|4165,4168|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|4173,4176|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4173,4176|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4173,4176|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4183,4186|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4183,4186|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|4183,4186|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4183,4186|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|4192,4195|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4192,4195|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|4203,4206|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|4203,4206|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|4203,4206|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|4203,4206|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4203,4206|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|4210,4213|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|4210,4213|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|4210,4213|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|4210,4213|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|4210,4213|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|4210,4213|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|4219,4223|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|4219,4223|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|4252,4255|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4272,4277|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4272,4277|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4272,4277|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|4282,4285|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|4282,4285|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|4282,4285|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Family Medical History|4308,4313|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4308,4313|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4308,4313|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|4308,4321|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|4308,4321|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|4308,4321|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|4314,4321|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4314,4321|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4314,4321|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4314,4321|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4314,4321|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4314,4321|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|4364,4368|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|4364,4368|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|4364,4368|false|false|false|C0202059|Bicarbonate measurement|HCO3
Attribute|Clinical Attribute|Family Medical History|4392,4400|false|false|false|C2926606||FINDINGS
Event|Event|Family Medical History|4392,4400|false|false|false|||FINDINGS
Finding|Functional Concept|Family Medical History|4392,4400|false|false|false|C2607943|findings aspects|FINDINGS
Event|Event|Family Medical History|4423,4426|true|false|false|||EGD
Procedure|Diagnostic Procedure|Family Medical History|4423,4426|true|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Family Medical History|4427,4435|false|false|false|||negative
Finding|Classification|Family Medical History|4427,4435|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Family Medical History|4427,4435|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Family Medical History|4427,4435|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Family Medical History|4427,4439|false|false|false|C0205160|Negative|negative for
Event|Event|Family Medical History|4440,4448|true|false|false|||evidence
Finding|Idea or Concept|Family Medical History|4440,4448|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Family Medical History|4440,4451|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Family Medical History|4452,4460|true|false|false|||bleeding
Finding|Pathologic Function|Family Medical History|4452,4460|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Body Substance|Family Medical History|4462,4471|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|4462,4471|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|4462,4471|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|4462,4471|true|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|Family Medical History|4472,4476|false|false|false|||LABS
Lab|Laboratory or Test Result|Family Medical History|4472,4476|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|4507,4512|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4507,4512|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4507,4512|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|4513,4516|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|4521,4524|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4521,4524|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4521,4524|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4531,4534|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4531,4534|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|4531,4534|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4531,4534|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|4540,4543|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4540,4543|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|4551,4554|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|4551,4554|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|4551,4554|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|4551,4554|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4551,4554|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|4558,4561|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|4558,4561|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|4558,4561|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|4558,4561|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|4558,4561|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|4558,4561|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|4567,4571|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|4567,4571|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|4600,4603|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|4620,4625|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4620,4625|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4620,4625|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|4630,4633|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|4630,4633|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|4630,4633|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Family Medical History|4656,4661|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4656,4661|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4656,4661|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|4656,4669|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|4656,4669|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|4656,4669|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|4662,4669|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4662,4669|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4662,4669|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4662,4669|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4662,4669|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4662,4669|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|4712,4716|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|4712,4716|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|4712,4716|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|4741,4746|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|4741,4746|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|4741,4746|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|4741,4754|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|4747,4754|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|4747,4754|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|4747,4754|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|4747,4754|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|4747,4754|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Family Medical History|4747,4754|false|false|false|||Calcium
Finding|Physiologic Function|Family Medical History|4747,4754|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|4747,4754|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4768,4772|false|false|false|C1431987|MCOLN1 protein, human|Mg-2
Drug|Biologically Active Substance|Family Medical History|4768,4772|false|false|false|C1431987|MCOLN1 protein, human|Mg-2
Finding|Gene or Genome|Family Medical History|4768,4772|false|false|false|C5890919|MCOLN1 wt Allele|Mg-2
Event|Event|Family Medical History|4777,4780|false|false|false|||PMH
Finding|Finding|Family Medical History|4777,4780|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|Family Medical History|4784,4787|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4784,4787|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|4784,4787|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|4784,4787|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|4784,4787|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|4784,4787|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|4784,4787|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4784,4787|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Family Medical History|4789,4792|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|Family Medical History|4789,4792|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4789,4792|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Disorder|Disease or Syndrome|Family Medical History|4798,4802|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Family Medical History|4798,4802|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Family Medical History|4798,4802|false|false|false|||COPD
Finding|Gene or Genome|Family Medical History|4798,4802|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Family Medical History|4807,4814|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|4807,4814|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4807,4814|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|4807,4814|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|4807,4817|false|false|false|C0262926|Medical History|history of
Event|Event|Family Medical History|4818,4827|false|false|false|||recurrent
Anatomy|Body Location or Region|Family Medical History|4828,4833|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|4828,4833|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Family Medical History|4835,4839|false|false|false|C2598155||pain
Event|Event|Family Medical History|4835,4839|false|false|false|||pain
Finding|Functional Concept|Family Medical History|4835,4839|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|4835,4839|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Family Medical History|4840,4847|false|false|false|||present
Finding|Finding|Family Medical History|4840,4847|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Family Medical History|4840,4847|false|false|false|C0150312;C0449450|Present;Presentation|present
Drug|Biomedical or Dental Material|Family Medical History|4853,4857|false|false|false|C0991568|Drops - Drug Form|drop
Event|Activity|Family Medical History|4853,4857|false|false|false|C1705648|Dropping|drop
Event|Event|Family Medical History|4853,4857|false|false|false|||drop
Event|Event|Family Medical History|4861,4864|false|false|false|||HCT
Procedure|Laboratory Procedure|Family Medical History|4861,4864|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4861,4864|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Finding|Functional Concept|Family Medical History|4869,4880|false|false|false|C0205329|Progressive|progressive
Event|Event|Family Medical History|4881,4884|false|false|false|||SOB
Finding|Sign or Symptom|Family Medical History|4881,4884|false|false|false|C0013404|Dyspnea|SOB
Event|Event|Family Medical History|4895,4903|false|false|false|||PROBLEMS
Finding|Idea or Concept|Family Medical History|4895,4903|false|false|false|C1546466|Problems - What subject filter|PROBLEMS
Finding|Pathologic Function|Family Medical History|4905,4913|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleed
Event|Event|Family Medical History|4908,4913|false|false|false|||Bleed
Finding|Pathologic Function|Family Medical History|4908,4913|false|false|false|C0019080|Hemorrhage|Bleed
Event|Event|Family Medical History|4915,4924|false|false|false|||Presented
Finding|Idea or Concept|Family Medical History|4915,4924|false|false|false|C0449450|Presentation|Presented
Disorder|Disease or Syndrome|Family Medical History|4928,4931|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Family Medical History|4928,4931|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Family Medical History|4928,4931|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4928,4931|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Family Medical History|4928,4931|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Family Medical History|4928,4931|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Family Medical History|4928,4931|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Family Medical History|4928,4931|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Family Medical History|4928,4931|false|false|false|||PCP
Finding|Gene or Genome|Family Medical History|4928,4931|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Family Medical History|4928,4931|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Family Medical History|4937,4943|false|false|false|||melena
Finding|Pathologic Function|Family Medical History|4937,4943|false|false|false|C0025222|Melena|melena
Event|Event|Family Medical History|4948,4954|false|false|false|||wiping
Disorder|Disease or Syndrome|Family Medical History|4955,4960|false|false|false|C0018932|Hematochezia|BRBPR
Event|Event|Family Medical History|4955,4960|false|false|false|||BRBPR
Anatomy|Cell Component|Family Medical History|4962,4965|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Family Medical History|4962,4965|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|Family Medical History|4971,4976|false|false|false|||taken
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4981,4984|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|4981,4984|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|Family Medical History|4981,4984|false|false|false|||Hgb
Finding|Gene or Genome|Family Medical History|4981,4984|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|4981,4984|false|false|false|C0019029|Hemoglobin concentration|Hgb
Event|Event|Family Medical History|4985,4990|false|false|false|||found
Event|Event|Family Medical History|4994,4998|false|false|false|||drop
Finding|Gene or Genome|Family Medical History|5019,5024|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|Family Medical History|5025,5029|false|false|false|||bore
Event|Event|Family Medical History|5031,5034|false|false|false|||IVs
Event|Event|Family Medical History|5040,5046|false|false|false|||placed
Event|Event|Family Medical History|5048,5055|false|false|false|||started
Finding|Finding|Family Medical History|5056,5061|false|false|false|C3714655|On IV|on IV
Drug|Pharmacologic Substance|Family Medical History|5062,5065|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|Family Medical History|5062,5065|false|false|false|||PPI
Finding|Physiologic Function|Family Medical History|5062,5065|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|Family Medical History|5079,5083|false|false|false|||type
Finding|Gene or Genome|Family Medical History|5079,5083|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Family Medical History|5079,5083|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Event|Event|Family Medical History|5089,5097|false|false|false|||screened
Event|Event|Family Medical History|5099,5105|false|false|false|||Vitals
Event|Event|Family Medical History|5115,5121|false|false|false|||stable
Finding|Intellectual Product|Family Medical History|5115,5121|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Body Substance|Family Medical History|5126,5133|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Family Medical History|5126,5133|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Family Medical History|5126,5133|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Family Medical History|5138,5147|false|false|false|||continued
Finding|Idea or Concept|Family Medical History|5152,5156|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|5152,5156|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|5152,5156|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|5157,5168|false|false|false|C1739768|rivaroxaban|rivaroxaban
Drug|Pharmacologic Substance|Family Medical History|5157,5168|false|false|false|C1739768|rivaroxaban|rivaroxaban
Event|Event|Family Medical History|5157,5168|false|false|false|||rivaroxaban
Event|Event|Family Medical History|5178,5187|false|false|false|||evaluated
Event|Event|Family Medical History|5198,5209|false|false|false|||recommended
Event|Event|Family Medical History|5220,5229|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|Family Medical History|5220,5229|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|Family Medical History|5237,5243|true|false|false|||showed
Event|Event|Family Medical History|5247,5255|true|false|false|||evidence
Finding|Idea or Concept|Family Medical History|5247,5255|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Family Medical History|5247,5258|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Family Medical History|5259,5267|true|false|false|||bleeding
Finding|Pathologic Function|Family Medical History|5259,5267|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Family Medical History|5273,5281|false|false|false|||remained
Finding|Finding|Family Medical History|5283,5305|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|Family Medical History|5299,5305|false|false|false|||stable
Finding|Intellectual Product|Family Medical History|5299,5305|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Family Medical History|5321,5330|false|false|false|||admission
Procedure|Health Care Activity|Family Medical History|5321,5330|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5332,5335|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|5332,5335|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|Family Medical History|5332,5335|false|false|false|||Hgb
Finding|Gene or Genome|Family Medical History|5332,5335|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|5332,5335|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Idea or Concept|Family Medical History|5343,5346|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Family Medical History|5343,5346|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Family Medical History|5351,5360|false|false|false|||discharge
Finding|Body Substance|Family Medical History|5351,5360|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Family Medical History|5351,5360|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Family Medical History|5351,5360|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Family Medical History|5351,5360|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Family Medical History|5370,5380|false|false|false|||discharged
Event|Event|Family Medical History|5381,5385|false|false|false|||home
Finding|Idea or Concept|Family Medical History|5381,5385|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|5381,5385|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|5381,5385|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|5398,5405|false|false|false|C3159309|Xarelto|Xarelto
Drug|Pharmacologic Substance|Family Medical History|5398,5405|false|false|false|C3159309|Xarelto|Xarelto
Drug|Amino Acid, Peptide, or Protein|Family Medical History|5411,5414|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Family Medical History|5411,5414|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Family Medical History|5411,5414|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Family Medical History|5411,5414|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Family Medical History|5411,5414|false|false|false|||ASA
Finding|Gene or Genome|Family Medical History|5411,5414|false|false|false|C1412553|ARSA gene|ASA
Event|Event|Family Medical History|5418,5421|false|false|false|||SOB
Finding|Sign or Symptom|Family Medical History|5418,5421|false|false|false|C0013404|Dyspnea|SOB
Event|Event|Family Medical History|5437,5444|false|false|false|||history
Finding|Conceptual Entity|Family Medical History|5437,5444|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|5437,5444|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|5437,5444|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|5437,5447|false|false|false|C0262926|Medical History|history of
Event|Event|Family Medical History|5448,5455|false|false|false|||smoking
Finding|Individual Behavior|Family Medical History|5448,5455|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|Family Medical History|5448,5455|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Disorder|Disease or Syndrome|Family Medical History|5460,5464|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Family Medical History|5460,5464|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Family Medical History|5460,5464|false|false|false|||COPD
Finding|Gene or Genome|Family Medical History|5460,5464|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Functional Concept|Family Medical History|5466,5477|false|false|false|C0205329|Progressive|Progressive
Finding|Sign or Symptom|Family Medical History|5479,5489|false|false|false|C0239313|exercise induced|exertional
Finding|Sign or Symptom|Family Medical History|5479,5497|false|true|false|C0231807|Dyspnea on exertion|exertional dyspnea
Event|Event|Family Medical History|5490,5497|false|false|false|||dyspnea
Finding|Finding|Family Medical History|5490,5497|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Family Medical History|5490,5497|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|Family Medical History|5506,5509|false|false|false|||use
Finding|Functional Concept|Family Medical History|5506,5509|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|5506,5509|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|Family Medical History|5506,5512|false|false|false|C1524063|Use of|use of
Drug|Organic Chemical|Family Medical History|5513,5520|false|false|false|C0905678|Spiriva|Spiriva
Drug|Pharmacologic Substance|Family Medical History|5513,5520|false|false|false|C0905678|Spiriva|Spiriva
Event|Event|Family Medical History|5513,5520|false|false|false|||Spiriva
Drug|Organic Chemical|Family Medical History|5522,5528|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|Family Medical History|5522,5528|false|false|false|C0965130|Advair|advair
Event|Event|Family Medical History|5522,5528|false|false|false|||advair
Drug|Organic Chemical|Family Medical History|5530,5541|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Family Medical History|5530,5541|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Family Medical History|5530,5541|false|false|false|||fluticasone
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|5543,5548|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Family Medical History|5543,5548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Family Medical History|5543,5548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Family Medical History|5543,5548|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Family Medical History|5543,5548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Family Medical History|5543,5548|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Pharmacologic Substance|Family Medical History|5543,5554|false|false|false|C2608294|Nasal Spray brand of phenylephrine|nasal spray
Drug|Biomedical or Dental Material|Family Medical History|5549,5554|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Family Medical History|5549,5554|false|false|false|C2003858|Spray (action)|spray
Event|Event|Family Medical History|5549,5554|false|false|false|||spray
Finding|Functional Concept|Family Medical History|5549,5554|false|false|false|C4521772|Spray (administration method)|spray
Drug|Organic Chemical|Family Medical History|5556,5568|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Family Medical History|5556,5568|false|false|false|C0039771|theophylline|theophylline
Event|Event|Family Medical History|5556,5568|false|false|false|||theophylline
Procedure|Laboratory Procedure|Family Medical History|5556,5568|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Family Medical History|5574,5583|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Family Medical History|5574,5583|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Family Medical History|5584,5594|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Family Medical History|5584,5594|false|false|false|||nebulizers
Finding|Functional Concept|Family Medical History|5618,5625|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Event|Event|Family Medical History|5626,5629|false|false|false|||use
Finding|Functional Concept|Family Medical History|5626,5629|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|5626,5629|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Conceptual Entity|Family Medical History|5632,5640|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|Family Medical History|5632,5640|true|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Event|Event|Family Medical History|5659,5665|true|false|false|||appear
Disorder|Disease or Syndrome|Family Medical History|5673,5683|true|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Family Medical History|5673,5683|true|false|false|||infectious
Event|Event|Family Medical History|5690,5700|true|false|false|||chronicity
Finding|Idea or Concept|Family Medical History|5702,5713|false|false|false|C0750501|most likely|Most likely
Finding|Finding|Family Medical History|5707,5713|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Family Medical History|5707,5713|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Family Medical History|5717,5728|false|false|false|||progression
Finding|Functional Concept|Family Medical History|5717,5728|false|true|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Family Medical History|5717,5728|false|true|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Family Medical History|5744,5748|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Family Medical History|5744,5748|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Family Medical History|5744,5748|false|false|false|||COPD
Finding|Gene or Genome|Family Medical History|5744,5748|false|false|false|C1412502|ARCN1 gene|COPD
Anatomy|Body Location or Region|Family Medical History|5750,5753|false|false|false|C5239891|area PFt|PFT
Drug|Indicator, Reagent, or Diagnostic Aid|Family Medical History|5750,5753|false|false|false|C0053122|bentiromide|PFT
Drug|Pharmacologic Substance|Family Medical History|5750,5753|false|false|false|C0053122|bentiromide|PFT
Event|Event|Family Medical History|5750,5753|false|false|false|||PFT
Procedure|Diagnostic Procedure|Family Medical History|5750,5753|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5750,5753|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Event|Event|Family Medical History|5761,5769|false|false|false|||obtained
Finding|Idea or Concept|Family Medical History|5776,5784|false|false|false|C4288901|In-House|in-house
Finding|Individual Behavior|Family Medical History|5786,5793|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Intellectual Product|Family Medical History|5786,5793|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Event|Activity|Family Medical History|5795,5804|false|false|true|C1880019|Cessation|cessation
Event|Event|Family Medical History|5795,5804|false|false|false|||cessation
Event|Event|Family Medical History|5814,5823|false|false|false|||discussed
Event|Event|Family Medical History|5830,5834|false|false|false|||need
Event|Event|Family Medical History|5835,5844|false|false|false|||continued
Event|Event|Family Medical History|5845,5855|false|false|false|||outpatient
Finding|Classification|Family Medical History|5845,5855|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Family Medical History|5845,5855|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Family Medical History|5869,5873|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Family Medical History|5869,5873|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Family Medical History|5869,5873|false|false|false|||COPD
Finding|Gene or Genome|Family Medical History|5869,5873|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Intellectual Product|Family Medical History|5876,5883|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Family Medical History|5876,5883|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Idea or Concept|Family Medical History|5884,5892|false|false|false|C1546466|Problems - What subject filter|PROBLEMS
Disorder|Disease or Syndrome|Family Medical History|5894,5898|false|false|false|C0004238|Atrial Fibrillation|Afib
Event|Event|Family Medical History|5894,5898|false|false|false|||Afib
Lab|Laboratory or Test Result|Family Medical History|5894,5898|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Event|Event|Family Medical History|5900,5909|false|false|false|||Continued
Finding|Idea or Concept|Family Medical History|5910,5914|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|5910,5914|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|5910,5914|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|5915,5925|false|false|false|C0002598|amiodarone|amiodarone
Drug|Pharmacologic Substance|Family Medical History|5915,5925|false|false|false|C0002598|amiodarone|amiodarone
Event|Event|Family Medical History|5915,5925|false|false|false|||amiodarone
Procedure|Laboratory Procedure|Family Medical History|5915,5925|false|false|false|C5399868|Drug assay amiodarone|amiodarone
Drug|Organic Chemical|Family Medical History|5930,5939|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Family Medical History|5930,5939|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Family Medical History|5930,5939|false|false|false|||diltiazem
Event|Event|Family Medical History|5941,5950|false|false|false|||Continued
Drug|Organic Chemical|Family Medical History|5952,5963|false|false|false|C1739768|rivaroxaban|rivaroxaban
Drug|Pharmacologic Substance|Family Medical History|5952,5963|false|false|false|C1739768|rivaroxaban|rivaroxaban
Event|Event|Family Medical History|5952,5963|false|false|false|||rivaroxaban
Event|Event|Family Medical History|5968,5983|false|false|false|||anticoagulation
Finding|Finding|Family Medical History|5968,5983|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Family Medical History|5968,5983|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Family Medical History|5968,5983|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Family Medical History|5988,5997|false|false|false|||discussed
Finding|Idea or Concept|Family Medical History|5998,6003|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|Family Medical History|6007,6010|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|6007,6010|false|false|false|||HTN
Event|Event|Family Medical History|6012,6018|false|false|false|||Stable
Finding|Intellectual Product|Family Medical History|6012,6018|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|Family Medical History|6020,6029|false|false|false|||continued
Finding|Idea or Concept|Family Medical History|6033,6037|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|6033,6037|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|6033,6037|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|6038,6047|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Family Medical History|6038,6047|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Family Medical History|6038,6047|false|false|false|||diltiazem
Drug|Organic Chemical|Family Medical History|6049,6054|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|Family Medical History|6049,6054|false|false|false|C0590690|Imdur|Imdur
Event|Event|Family Medical History|6049,6054|false|false|false|||Imdur
Drug|Organic Chemical|Family Medical History|6056,6060|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Family Medical History|6056,6060|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|Family Medical History|6056,6060|false|false|false|||HCTZ
Disorder|Mental or Behavioral Dysfunction|Family Medical History|6063,6070|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Family Medical History|6063,6070|false|false|false|||Anxiety
Finding|Sign or Symptom|Family Medical History|6063,6070|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Pharmacologic Substance|Family Medical History|6071,6079|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Family Medical History|6071,6079|false|false|false|||insomnia
Finding|Sign or Symptom|Family Medical History|6071,6079|false|false|false|C0917801|Sleeplessness|insomnia
Event|Event|Family Medical History|6081,6087|false|false|false|||stable
Finding|Intellectual Product|Family Medical History|6081,6087|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Family Medical History|6089,6098|false|false|false|||continued
Finding|Idea or Concept|Family Medical History|6099,6103|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|6099,6103|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|6099,6103|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|6104,6113|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Family Medical History|6104,6113|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Family Medical History|6114,6117|false|false|false|||QHS
Finding|Gene or Genome|Family Medical History|6118,6121|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Family Medical History|6127,6135|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Family Medical History|6127,6135|false|false|false|||insomnia
Finding|Sign or Symptom|Family Medical History|6127,6135|false|false|false|C0917801|Sleeplessness|insomnia
Disorder|Mental or Behavioral Dysfunction|Family Medical History|6136,6143|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Family Medical History|6136,6143|false|false|false|||anxiety
Finding|Sign or Symptom|Family Medical History|6136,6143|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Disease or Syndrome|Family Medical History|6147,6155|false|false|false|C0013238;C0022575|Dry Eye Syndromes;Keratoconjunctivitis Sicca|Dry eyes
Drug|Pharmacologic Substance|Family Medical History|6147,6155|false|false|false|C0720056|Dry Eyes brand of ocular lubricant|Dry eyes
Finding|Sign or Symptom|Family Medical History|6147,6155|false|false|false|C0314719|Dryness of eye|Dry eyes
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6151,6155|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|Family Medical History|6151,6155|false|false|false|C5848506||eyes
Event|Event|Family Medical History|6151,6155|false|false|false|||eyes
Event|Event|Family Medical History|6157,6164|false|false|false|||History
Finding|Conceptual Entity|Family Medical History|6157,6164|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Family Medical History|6157,6164|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Family Medical History|6157,6164|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Family Medical History|6157,6167|false|false|false|C0262926|Medical History|History of
Finding|Finding|Family Medical History|6157,6176|false|false|false|C0455517||History of glaucoma
Disorder|Disease or Syndrome|Family Medical History|6168,6176|false|false|false|C0017601|Glaucoma|glaucoma
Event|Event|Family Medical History|6168,6176|false|false|false|||glaucoma
Event|Event|Family Medical History|6178,6187|false|false|false|||Continued
Finding|Idea or Concept|Family Medical History|6188,6192|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|6188,6192|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|6188,6192|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|6193,6204|false|false|false|C0090306|latanoprost|latanoprost
Drug|Pharmacologic Substance|Family Medical History|6193,6204|false|false|false|C0090306|latanoprost|latanoprost
Event|Event|Family Medical History|6193,6204|false|false|false|||latanoprost
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6206,6216|false|false|false|C0015392|Eye|ophthalmic
Drug|Biomedical or Dental Material|Family Medical History|6206,6216|false|false|false|C2347396|Ophthalmic Dosage Form|ophthalmic
Finding|Functional Concept|Family Medical History|6206,6216|false|false|false|C1522230|Ophthalmic Route of Administration|ophthalmic
Drug|Biomedical or Dental Material|Family Medical History|6206,6222|false|false|false|C0015399|Eye Drops|ophthalmic drops
Drug|Biomedical or Dental Material|Family Medical History|6217,6222|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|Family Medical History|6217,6222|false|false|false|||drops
Anatomy|Anatomical Structure|Family Medical History|6226,6229|false|false|false|C3669270|Strucure of thick cushion of skin|PAD
Disorder|Disease or Syndrome|Family Medical History|6226,6229|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Disorder|Neoplastic Process|Family Medical History|6226,6229|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|PAD
Drug|Biomedical or Dental Material|Family Medical History|6226,6229|false|false|false|C2347441|Pad Dosage Form|PAD
Event|Event|Family Medical History|6226,6229|false|false|false|||PAD
Finding|Gene or Genome|Family Medical History|6226,6229|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|PAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|6226,6229|false|false|false|C3814046|PAD Regimen|PAD
Event|Event|Family Medical History|6231,6237|false|false|false|||Stable
Finding|Intellectual Product|Family Medical History|6231,6237|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|Family Medical History|6239,6248|false|false|false|||continued
Finding|Idea or Concept|Family Medical History|6252,6256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|6252,6256|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|6252,6256|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|6257,6269|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Family Medical History|6257,6269|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Family Medical History|6257,6269|false|false|false|||atorvastatin
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|6275,6280|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Family Medical History|6275,6286|false|false|false|C0850459|iliac stents|iliac stent
Event|Event|Family Medical History|6281,6286|false|false|false|||stent
Event|Event|Family Medical History|6295,6303|false|false|false|||continue
Drug|Organic Chemical|Family Medical History|6304,6311|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Family Medical History|6304,6311|false|false|false|C0004057|aspirin|aspirin
Event|Event|Family Medical History|6304,6311|false|false|false|||aspirin
Finding|Finding|Family Medical History|6315,6319|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|Family Medical History|6322,6334|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Family Medical History|6335,6341|false|false|false|||ISSUES
Event|Event|Family Medical History|6352,6360|true|false|false|||consider
Finding|Classification|Family Medical History|6361,6371|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Family Medical History|6361,6371|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Family Medical History|6372,6383|true|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Family Medical History|6372,6383|true|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Family Medical History|6372,6383|true|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|Family Medical History|6399,6407|true|false|false|||identify
Event|Event|Family Medical History|6413,6419|true|false|false|||source
Finding|Finding|Family Medical History|6413,6419|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|Family Medical History|6413,6419|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|Family Medical History|6413,6419|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Anatomy|Body Location or Region|Family Medical History|6423,6428|true|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Family Medical History|6423,6428|true|false|false|C2003888|Lower (action)|lower
Finding|Pathologic Function|Family Medical History|6423,6437|true|false|false|C0024050|Lower gastrointestinal hemorrhage|lower GI Bleed
Finding|Pathologic Function|Family Medical History|6429,6437|true|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleed
Event|Event|Family Medical History|6432,6437|true|false|false|||Bleed
Finding|Pathologic Function|Family Medical History|6432,6437|true|false|false|C0019080|Hemorrhage|Bleed
Event|Event|Family Medical History|6447,6453|false|false|false|||stable
Finding|Intellectual Product|Family Medical History|6447,6453|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|Family Medical History|6447,6464|false|false|false|C1370135|Hemoglobin.stable|stable hemoglobin
Drug|Amino Acid, Peptide, or Protein|Family Medical History|6454,6464|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Family Medical History|6454,6464|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Family Medical History|6454,6464|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Family Medical History|6454,6464|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|Family Medical History|6454,6464|false|false|false|||hemoglobin
Finding|Finding|Family Medical History|6454,6464|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Family Medical History|6454,6464|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Attribute|Clinical Attribute|Family Medical History|6465,6475|false|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|Family Medical History|6465,6475|false|false|false|||hematocrit
Finding|Finding|Family Medical History|6465,6475|false|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|Family Medical History|6465,6475|false|false|false|C0018935|Hematocrit Measurement|hematocrit
Event|Event|Family Medical History|6482,6491|true|false|false|||inpatient
Finding|Idea or Concept|Family Medical History|6482,6491|true|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Family Medical History|6482,6491|true|false|false|C1555324|inpatient encounter|inpatient
Finding|Finding|Family Medical History|6495,6499|true|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|6507,6515|true|false|false|||evidence
Finding|Idea or Concept|Family Medical History|6507,6515|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Family Medical History|6507,6518|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Family Medical History|6519,6527|true|false|false|||bleeding
Finding|Pathologic Function|Family Medical History|6519,6527|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Family Medical History|6531,6534|true|false|false|||EGD
Procedure|Diagnostic Procedure|Family Medical History|6531,6534|true|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Drug|Organic Chemical|Family Medical History|6540,6547|false|false|false|C3159309|Xarelto|Xarelto
Drug|Pharmacologic Substance|Family Medical History|6540,6547|false|false|false|C3159309|Xarelto|Xarelto
Drug|Organic Chemical|Family Medical History|6552,6559|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Family Medical History|6552,6559|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Family Medical History|6566,6575|false|false|false|||continued
Event|Event|Family Medical History|6579,6588|false|false|false|||discharge
Finding|Body Substance|Family Medical History|6579,6588|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Family Medical History|6579,6588|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Family Medical History|6579,6588|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Family Medical History|6579,6588|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Family Medical History|6595,6602|false|false|false|||treated
Drug|Pharmacologic Substance|Family Medical History|6611,6614|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|Family Medical History|6611,6614|false|false|false|||PPI
Finding|Physiologic Function|Family Medical History|6611,6614|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|Family Medical History|6621,6630|false|false|false|||inpatient
Finding|Idea or Concept|Family Medical History|6621,6630|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Family Medical History|6621,6630|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|Family Medical History|6645,6653|true|false|false|||evidence
Finding|Idea or Concept|Family Medical History|6645,6653|true|false|false|C3887511|Evidence|evidence
Event|Event|Family Medical History|6665,6673|true|false|false|||bleeding
Finding|Pathologic Function|Family Medical History|6665,6673|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Family Medical History|6679,6689|false|false|false|||discharged
Finding|Idea or Concept|Family Medical History|6693,6697|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Family Medical History|6693,6697|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Family Medical History|6693,6697|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Family Medical History|6698,6708|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Family Medical History|6698,6708|false|false|false|C0034665|ranitidine|Ranitidine
Event|Event|Family Medical History|6709,6714|false|false|false|||300mg
Event|Event|Family Medical History|6727,6735|false|false|false|||Continue
Finding|Idea or Concept|Family Medical History|6727,6735|false|false|false|C0549178|Continuous|Continue
Event|Event|Family Medical History|6739,6748|false|false|false|||encourage
Procedure|Health Care Activity|Family Medical History|6739,6766|false|false|false|C0510865|Encourage smoking cessation|encourage smoking cessation
Event|Event|Family Medical History|6749,6756|false|false|false|||smoking
Finding|Individual Behavior|Family Medical History|6749,6766|false|false|false|C0085134|Cessation of smoking|smoking cessation
Procedure|Therapeutic or Preventive Procedure|Family Medical History|6749,6766|false|false|false|C1095963|Smoking cessation therapy|smoking cessation
Event|Activity|Family Medical History|6757,6766|false|false|true|C1880019|Cessation|cessation
Event|Event|Family Medical History|6757,6766|false|false|false|||cessation
Attribute|Clinical Attribute|Family Medical History|6770,6781|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Family Medical History|6770,6781|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Family Medical History|6770,6781|false|false|false|||Medications
Finding|Intellectual Product|Family Medical History|6770,6781|false|false|false|C4284232|Medications|Medications
Finding|Finding|Family Medical History|6770,6794|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Family Medical History|6785,6794|false|false|false|||Admission
Procedure|Health Care Activity|Family Medical History|6785,6794|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Family Medical History|6813,6823|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Family Medical History|6813,6823|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Family Medical History|6813,6828|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Family Medical History|6824,6828|false|false|false|||list
Finding|Intellectual Product|Family Medical History|6824,6828|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Family Medical History|6832,6840|false|false|false|||accurate
Drug|Organic Chemical|Family Medical History|6845,6853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Family Medical History|6845,6853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Family Medical History|6845,6853|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Family Medical History|6845,6853|false|false|false|||complete
Finding|Functional Concept|Family Medical History|6845,6853|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Family Medical History|6845,6853|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Family Medical History|6858,6869|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Family Medical History|6858,6869|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Family Medical History|6879,6882|false|false|false|||QPM
Drug|Organic Chemical|Family Medical History|6887,6900|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Family Medical History|6887,6900|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Family Medical History|6887,6900|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Family Medical History|6887,6900|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Family Medical History|6915,6918|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Family Medical History|6919,6923|false|false|false|C2598155||pain
Event|Event|Family Medical History|6919,6923|false|false|false|||pain
Finding|Functional Concept|Family Medical History|6919,6923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|6919,6923|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Family Medical History|6928,6937|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Family Medical History|6928,6937|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Family Medical History|6945,6948|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Family Medical History|6945,6948|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Family Medical History|6945,6948|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Family Medical History|6945,6948|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Family Medical History|6945,6948|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Family Medical History|6956,6959|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Family Medical History|6956,6959|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Family Medical History|6956,6959|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Family Medical History|6956,6959|false|false|false|||NEB
Finding|Cell Function|Family Medical History|6956,6959|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Family Medical History|6956,6959|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Family Medical History|6967,6970|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Family Medical History|6971,6974|false|false|false|||SOB
Finding|Sign or Symptom|Family Medical History|6971,6974|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Family Medical History|6979,6986|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Family Medical History|6979,6986|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Family Medical History|7006,7018|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Family Medical History|7006,7018|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Family Medical History|7036,7045|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Family Medical History|7036,7045|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Family Medical History|7046,7054|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Family Medical History|7046,7054|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Family Medical History|7055,7062|false|false|false|||Release
Finding|Functional Concept|Family Medical History|7055,7062|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Family Medical History|7055,7062|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Family Medical History|7055,7062|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7073,7076|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7073,7076|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7073,7076|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7073,7076|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7073,7076|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|7081,7092|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|7081,7092|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Family Medical History|7081,7092|false|false|false|||Fluticasone
Drug|Organic Chemical|Family Medical History|7081,7103|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Family Medical History|7081,7103|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Family Medical History|7093,7103|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7104,7109|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Family Medical History|7104,7109|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Family Medical History|7104,7109|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Family Medical History|7104,7109|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Family Medical History|7104,7109|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Family Medical History|7104,7109|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Family Medical History|7112,7116|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7120,7123|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7120,7123|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7120,7123|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7120,7123|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7120,7123|false|false|false|C1332410|BID gene|BID
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7124,7129|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Family Medical History|7124,7129|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Family Medical History|7124,7129|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Family Medical History|7124,7129|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Family Medical History|7124,7129|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Family Medical History|7124,7129|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Family Medical History|7124,7140|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|Family Medical History|7130,7140|false|false|false|||congestion
Finding|Pathologic Function|Family Medical History|7130,7140|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Family Medical History|7145,7156|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|7145,7156|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|7145,7167|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Family Medical History|7145,7174|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Family Medical History|7145,7174|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Family Medical History|7157,7167|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Family Medical History|7157,7167|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Family Medical History|7168,7174|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Family Medical History|7187,7190|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Family Medical History|7187,7190|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Family Medical History|7187,7190|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Family Medical History|7187,7190|false|false|false|||INH
Finding|Functional Concept|Family Medical History|7187,7190|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7194,7197|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7194,7197|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7194,7197|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7194,7197|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7194,7197|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|7202,7221|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Family Medical History|7202,7221|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Family Medical History|7242,7252|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Family Medical History|7242,7252|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Family Medical History|7242,7264|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Family Medical History|7242,7264|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Family Medical History|7253,7264|false|false|false|||Mononitrate
Finding|Finding|Family Medical History|7266,7274|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Family Medical History|7266,7274|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Family Medical History|7275,7282|false|false|false|||Release
Finding|Functional Concept|Family Medical History|7275,7282|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Family Medical History|7275,7282|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Family Medical History|7275,7282|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Family Medical History|7305,7316|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Family Medical History|7305,7316|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Family Medical History|7324,7329|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Family Medical History|7339,7343|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Family Medical History|7339,7343|false|false|false|C1705648|Dropping|DROP
Event|Event|Family Medical History|7344,7348|false|false|false|||LEFT
Finding|Functional Concept|Family Medical History|7344,7348|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7344,7352|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Family Medical History|7344,7352|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Family Medical History|7349,7352|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7349,7352|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Family Medical History|7349,7352|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Family Medical History|7349,7352|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Family Medical History|7349,7352|false|false|false|||EYE
Finding|Body Substance|Family Medical History|7349,7352|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Family Medical History|7349,7352|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Family Medical History|7349,7352|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|Family Medical History|7353,7356|false|false|false|||QHS
Drug|Organic Chemical|Family Medical History|7362,7371|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Family Medical History|7362,7371|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Family Medical History|7382,7385|false|false|false|||QHS
Finding|Gene or Genome|Family Medical History|7386,7389|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Family Medical History|7390,7398|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Family Medical History|7390,7398|false|false|false|||insomnia
Finding|Sign or Symptom|Family Medical History|7390,7398|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Family Medical History|7404,7417|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Family Medical History|7404,7417|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Family Medical History|7404,7417|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Family Medical History|7404,7417|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Family Medical History|7420,7428|false|false|false|C0026162|Minerals|minerals
Event|Event|Family Medical History|7420,7428|false|false|false|||minerals
Drug|Biomedical or Dental Material|Family Medical History|7431,7434|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Family Medical History|7431,7434|false|false|false|||TAB
Drug|Organic Chemical|Family Medical History|7449,7459|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Family Medical History|7449,7459|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Family Medical History|7481,7493|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Family Medical History|7481,7493|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Family Medical History|7481,7493|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Family Medical History|7481,7493|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Family Medical History|7481,7496|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Family Medical History|7481,7496|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|Family Medical History|7494,7496|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7507,7510|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7507,7510|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7507,7510|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7507,7510|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7507,7510|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|7516,7526|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Family Medical History|7516,7526|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Family Medical History|7516,7526|false|false|false|||Tiotropium
Drug|Organic Chemical|Family Medical History|7516,7534|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Family Medical History|7516,7534|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Family Medical History|7527,7534|false|false|false|C0006222|Bromides|Bromide
Event|Event|Family Medical History|7527,7534|false|false|false|||Bromide
Procedure|Laboratory Procedure|Family Medical History|7527,7534|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Family Medical History|7537,7540|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Family Medical History|7537,7540|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Family Medical History|7537,7540|false|false|false|||CAP
Finding|Gene or Genome|Family Medical History|7537,7540|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Family Medical History|7537,7540|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7544,7547|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7544,7547|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7544,7547|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7544,7547|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7544,7547|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|7553,7561|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|Family Medical History|7553,7561|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|Family Medical History|7553,7561|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|Family Medical History|7553,7561|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|Family Medical History|7563,7569|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|Family Medical History|7563,7569|false|false|false|C0724054|Ultram|Ultram
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7580,7583|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7580,7583|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7580,7583|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7580,7583|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7580,7583|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|Family Medical History|7584,7588|false|false|false|C2598155||pain
Event|Event|Family Medical History|7584,7588|false|false|false|||pain
Finding|Functional Concept|Family Medical History|7584,7588|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|7584,7588|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Family Medical History|7594,7610|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Family Medical History|7605,7610|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Family Medical History|7605,7610|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Event|Event|Family Medical History|7611,7618|false|false|false|||Preserv
Finding|Functional Concept|Family Medical History|7611,7618|false|false|false|C0728887|Preserving|Preserv
Procedure|Laboratory Procedure|Family Medical History|7611,7618|false|false|false|C0033085|Biologic Preservation|Preserv
Finding|Functional Concept|Family Medical History|7620,7624|false|false|false|C0332296|Free of (attribute)|Free
Drug|Biomedical or Dental Material|Family Medical History|7629,7633|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Family Medical History|7629,7633|false|false|false|C1705648|Dropping|DROP
Event|Event|Family Medical History|7629,7633|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7634,7643|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7639,7643|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Family Medical History|7639,7643|false|false|false|C5848506||EYES
Event|Event|Family Medical History|7644,7647|false|false|false|||PRN
Finding|Gene or Genome|Family Medical History|7644,7647|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Family Medical History|7649,7659|false|false|false|||irritation
Finding|Intellectual Product|Family Medical History|7649,7659|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Family Medical History|7649,7659|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Family Medical History|7649,7659|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Family Medical History|7649,7659|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Family Medical History|7665,7675|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Family Medical History|7665,7675|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Family Medical History|7665,7675|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Family Medical History|7665,7675|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Event|Event|Family Medical History|7696,7705|false|false|false|||Discharge
Finding|Body Substance|Family Medical History|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Family Medical History|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Family Medical History|7696,7705|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Family Medical History|7696,7705|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Family Medical History|7696,7717|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Family Medical History|7706,7717|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Family Medical History|7706,7717|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Family Medical History|7706,7717|false|false|false|||Medications
Finding|Intellectual Product|Family Medical History|7706,7717|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Family Medical History|7722,7735|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Family Medical History|7722,7735|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Family Medical History|7722,7735|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Family Medical History|7722,7735|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Family Medical History|7750,7753|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Family Medical History|7754,7758|false|false|false|C2598155||pain
Event|Event|Family Medical History|7754,7758|false|false|false|||pain
Finding|Functional Concept|Family Medical History|7754,7758|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|7754,7758|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Family Medical History|7763,7772|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Family Medical History|7763,7772|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7780,7783|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Family Medical History|7780,7783|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Family Medical History|7780,7783|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Family Medical History|7780,7783|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Family Medical History|7780,7783|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7791,7794|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Family Medical History|7791,7794|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Family Medical History|7791,7794|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Family Medical History|7791,7794|false|false|false|||NEB
Finding|Cell Function|Family Medical History|7791,7794|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Family Medical History|7791,7794|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Family Medical History|7802,7805|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Family Medical History|7806,7809|false|false|false|||SOB
Finding|Sign or Symptom|Family Medical History|7806,7809|false|false|false|C0013404|Dyspnea|SOB
Drug|Organic Chemical|Family Medical History|7814,7824|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Family Medical History|7814,7824|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Family Medical History|7814,7824|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Family Medical History|7814,7824|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Family Medical History|7845,7857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Family Medical History|7845,7857|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Family Medical History|7875,7891|false|false|false|C0003921;C2608262;C3853661|Artificial Tears;Lubricant Eye Drops;artificial tears (medication)|Artificial Tears
Finding|Body Substance|Family Medical History|7886,7891|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Finding|Intellectual Product|Family Medical History|7886,7891|false|false|false|C0039409;C1547924;C1611838|Tears (substance);Tears specimen|Tears
Event|Event|Family Medical History|7892,7899|false|false|false|||Preserv
Finding|Functional Concept|Family Medical History|7892,7899|false|false|false|C0728887|Preserving|Preserv
Procedure|Laboratory Procedure|Family Medical History|7892,7899|false|false|false|C0033085|Biologic Preservation|Preserv
Finding|Functional Concept|Family Medical History|7901,7905|false|false|false|C0332296|Free of (attribute)|Free
Drug|Biomedical or Dental Material|Family Medical History|7910,7914|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Family Medical History|7910,7914|false|false|false|C1705648|Dropping|DROP
Event|Event|Family Medical History|7910,7914|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7915,7924|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|7920,7924|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Family Medical History|7920,7924|false|false|false|C5848506||EYES
Event|Event|Family Medical History|7925,7928|false|false|false|||PRN
Finding|Gene or Genome|Family Medical History|7925,7928|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Family Medical History|7930,7940|false|false|false|||irritation
Finding|Intellectual Product|Family Medical History|7930,7940|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Mental Process|Family Medical History|7930,7940|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Finding|Pathologic Function|Family Medical History|7930,7940|false|false|false|C1706307;C2700617;C5575347|Have Vulvar Irritation question;Irritability - emotion;Irritation (finding)|irritation
Phenomenon|Phenomenon or Process|Family Medical History|7930,7940|false|false|false|C0441723|Irritation|irritation
Drug|Organic Chemical|Family Medical History|7945,7954|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Family Medical History|7945,7954|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Family Medical History|7955,7963|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Family Medical History|7955,7963|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Family Medical History|7964,7971|false|false|false|||Release
Finding|Functional Concept|Family Medical History|7964,7971|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Family Medical History|7964,7971|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Family Medical History|7964,7971|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Family Medical History|7982,7985|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|7982,7985|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|7982,7985|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|7982,7985|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|7982,7985|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|7990,8001|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|7990,8001|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Family Medical History|7990,8001|false|false|false|||Fluticasone
Drug|Organic Chemical|Family Medical History|7990,8012|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Family Medical History|7990,8012|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Family Medical History|8002,8012|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|8013,8018|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Family Medical History|8013,8018|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Family Medical History|8013,8018|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Family Medical History|8013,8018|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Family Medical History|8013,8018|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Family Medical History|8013,8018|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Family Medical History|8021,8025|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|Family Medical History|8029,8032|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8029,8032|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|8029,8032|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|8029,8032|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|8029,8032|false|false|false|C1332410|BID gene|BID
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|8033,8038|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Family Medical History|8033,8038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Family Medical History|8033,8038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Family Medical History|8033,8038|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Family Medical History|8033,8038|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Family Medical History|8033,8038|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|Family Medical History|8033,8049|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|Family Medical History|8039,8049|false|false|false|||congestion
Finding|Pathologic Function|Family Medical History|8039,8049|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Family Medical History|8054,8065|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|8054,8065|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Family Medical History|8054,8076|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Family Medical History|8054,8083|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Family Medical History|8054,8083|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Family Medical History|8066,8076|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Family Medical History|8066,8076|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Family Medical History|8077,8083|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Family Medical History|8096,8099|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Family Medical History|8096,8099|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Family Medical History|8096,8099|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Family Medical History|8096,8099|false|false|false|||INH
Finding|Functional Concept|Family Medical History|8096,8099|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Family Medical History|8103,8106|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8103,8106|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|8103,8106|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|8103,8106|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|8103,8106|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|8111,8130|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Family Medical History|8111,8130|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Family Medical History|8151,8161|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Family Medical History|8151,8161|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Family Medical History|8151,8173|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Family Medical History|8151,8173|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Family Medical History|8162,8173|false|false|false|||Mononitrate
Finding|Finding|Family Medical History|8175,8183|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Family Medical History|8175,8183|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Family Medical History|8184,8191|false|false|false|||Release
Finding|Functional Concept|Family Medical History|8184,8191|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Family Medical History|8184,8191|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Family Medical History|8184,8191|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Family Medical History|8214,8225|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Family Medical History|8214,8225|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Family Medical History|8233,8238|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Family Medical History|8248,8252|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Family Medical History|8248,8252|false|false|false|C1705648|Dropping|DROP
Event|Event|Family Medical History|8253,8257|false|false|false|||LEFT
Finding|Functional Concept|Family Medical History|8253,8257|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|8253,8261|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Family Medical History|8253,8261|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Family Medical History|8258,8261|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|8258,8261|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Family Medical History|8258,8261|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Family Medical History|8258,8261|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Family Medical History|8258,8261|false|false|false|||EYE
Finding|Body Substance|Family Medical History|8258,8261|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Family Medical History|8258,8261|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Family Medical History|8258,8261|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Event|Event|Family Medical History|8262,8265|false|false|false|||QHS
Drug|Organic Chemical|Family Medical History|8271,8280|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Family Medical History|8271,8280|false|false|false|C0024002|lorazepam|Lorazepam
Event|Event|Family Medical History|8291,8294|false|false|false|||QHS
Finding|Gene or Genome|Family Medical History|8295,8298|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Pharmacologic Substance|Family Medical History|8299,8307|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Family Medical History|8299,8307|false|false|false|||insomnia
Finding|Sign or Symptom|Family Medical History|8299,8307|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Family Medical History|8313,8324|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Drug|Pharmacologic Substance|Family Medical History|8313,8324|false|false|false|C1739768|rivaroxaban|Rivaroxaban
Event|Event|Family Medical History|8334,8337|false|false|false|||QPM
Drug|Organic Chemical|Family Medical History|8343,8355|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Family Medical History|8343,8355|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Family Medical History|8343,8355|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Family Medical History|8343,8355|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Family Medical History|8343,8358|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Family Medical History|8343,8358|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|Family Medical History|8356,8358|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|Family Medical History|8369,8372|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8369,8372|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|8369,8372|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|8369,8372|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|8369,8372|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|8378,8388|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Family Medical History|8378,8388|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Family Medical History|8410,8418|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|Family Medical History|8410,8418|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|Family Medical History|8410,8418|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|Family Medical History|8410,8418|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|Family Medical History|8420,8426|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|Family Medical History|8420,8426|false|false|false|C0724054|Ultram|Ultram
Disorder|Mental or Behavioral Dysfunction|Family Medical History|8437,8440|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8437,8440|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|8437,8440|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|8437,8440|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|8437,8440|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|Family Medical History|8441,8445|false|false|false|C2598155||pain
Event|Event|Family Medical History|8441,8445|false|false|false|||pain
Finding|Functional Concept|Family Medical History|8441,8445|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Family Medical History|8441,8445|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Family Medical History|8451,8461|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Family Medical History|8451,8461|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Family Medical History|8451,8461|false|false|false|||Tiotropium
Drug|Organic Chemical|Family Medical History|8451,8469|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Family Medical History|8451,8469|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Family Medical History|8462,8469|false|false|false|C0006222|Bromides|Bromide
Event|Event|Family Medical History|8462,8469|false|false|false|||Bromide
Procedure|Laboratory Procedure|Family Medical History|8462,8469|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Family Medical History|8472,8475|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Family Medical History|8472,8475|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Family Medical History|8472,8475|false|false|false|||CAP
Finding|Gene or Genome|Family Medical History|8472,8475|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Family Medical History|8472,8475|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Disorder|Mental or Behavioral Dysfunction|Family Medical History|8479,8482|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8479,8482|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Family Medical History|8479,8482|false|false|false|C1530795|BID protein, human|BID
Event|Event|Family Medical History|8479,8482|false|false|false|||BID
Finding|Gene or Genome|Family Medical History|8479,8482|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Family Medical History|8488,8501|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Family Medical History|8488,8501|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Family Medical History|8488,8501|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Family Medical History|8488,8501|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Family Medical History|8504,8512|false|false|false|C0026162|Minerals|minerals
Event|Event|Family Medical History|8504,8512|false|false|false|||minerals
Drug|Biomedical or Dental Material|Family Medical History|8515,8518|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Family Medical History|8515,8518|false|false|false|||TAB
Drug|Organic Chemical|Family Medical History|8533,8540|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Family Medical History|8533,8540|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Family Medical History|8560,8569|false|false|false|||Discharge
Finding|Body Substance|Family Medical History|8560,8569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Family Medical History|8560,8569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Family Medical History|8560,8569|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Family Medical History|8560,8569|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Family Medical History|8560,8581|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Family Medical History|8560,8581|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Family Medical History|8570,8581|false|false|false|C2926604||Disposition
Event|Event|Family Medical History|8570,8581|false|false|false|||Disposition
Procedure|Health Care Activity|Family Medical History|8570,8581|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Family Medical History|8583,8587|false|false|false|||Home
Finding|Idea or Concept|Family Medical History|8583,8587|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Family Medical History|8583,8587|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Family Medical History|8583,8587|false|false|false|C1553498|home health encounter|Home
Event|Event|Family Medical History|8590,8599|false|false|false|||Discharge
Finding|Body Substance|Family Medical History|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Family Medical History|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Family Medical History|8590,8599|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Family Medical History|8590,8599|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Family Medical History|8590,8609|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Family Medical History|8600,8609|false|false|false|C0945731||Diagnosis
Event|Event|Family Medical History|8600,8609|false|false|false|||Diagnosis
Finding|Classification|Family Medical History|8600,8609|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Family Medical History|8600,8609|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Family Medical History|8600,8609|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Family Medical History|8622,8628|false|false|false|C0002871|Anemia|Anemia
Event|Event|Family Medical History|8622,8628|false|false|false|||Anemia
Disorder|Neoplastic Process|Family Medical History|8630,8639|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Family Medical History|8630,8639|false|false|false|||Secondary
Finding|Functional Concept|Family Medical History|8630,8639|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|Family Medical History|8643,8647|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|Family Medical History|8643,8647|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Disorder|Disease or Syndrome|Family Medical History|8650,8653|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|8650,8653|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|8650,8653|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|8650,8653|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|8650,8653|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|8650,8653|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|8650,8653|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|8650,8653|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Family Medical History|8656,8659|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|8656,8659|false|false|false|||HTN
Disorder|Disease or Syndrome|Family Medical History|8662,8666|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Family Medical History|8662,8666|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Family Medical History|8662,8666|false|false|false|||COPD
Finding|Gene or Genome|Family Medical History|8662,8666|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Mental Process|Discharge Condition|8691,8697|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8691,8704|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8691,8704|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8698,8704|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8698,8704|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8706,8711|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|8706,8711|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|8716,8724|false|false|false|||coherent
Finding|Finding|Discharge Condition|8716,8724|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|8726,8731|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8726,8748|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8726,8748|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8735,8748|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8735,8748|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8735,8748|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8750,8755|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8750,8755|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8750,8755|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8750,8755|false|false|false|||Alert
Finding|Finding|Discharge Condition|8750,8755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8750,8755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8750,8755|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8760,8771|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8760,8771|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8773,8781|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8773,8781|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8773,8781|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8782,8788|false|false|false|C5889824||Status
Event|Event|Discharge Condition|8782,8788|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|8782,8788|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8790,8800|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|8790,8800|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8790,8800|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8790,8800|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8790,8800|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|8803,8814|false|false|false|||Independent
Finding|Finding|Discharge Condition|8803,8814|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8803,8814|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|8862,8870|false|false|false|||admitted
Event|Event|Discharge Instructions|8888,8896|false|false|false|||decrease
Finding|Finding|Discharge Instructions|8888,8896|false|false|false|C0392756|Reduced|decrease
Finding|Body Substance|Discharge Instructions|8897,8905|false|false|false|C0005768|In Blood|in blood
Disorder|Disease or Syndrome|Discharge Instructions|8900,8905|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|8900,8905|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|8900,8905|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|8900,8911|false|false|false|C0005771|Blood Cell Count|blood count
Event|Event|Discharge Instructions|8906,8911|false|false|false|||count
Attribute|Clinical Attribute|Discharge Instructions|8915,8925|false|false|false|C2598148||laboratory
Finding|Functional Concept|Discharge Instructions|8915,8925|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Finding|Intellectual Product|Discharge Instructions|8915,8925|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Lab|Laboratory or Test Result|Discharge Instructions|8915,8925|false|false|false|C4283904|Laboratory observation|laboratory
Procedure|Laboratory Procedure|Discharge Instructions|8915,8933|false|false|false|C0022885|Laboratory Procedures|laboratory testing
Event|Event|Discharge Instructions|8926,8933|false|false|false|||testing
Finding|Functional Concept|Discharge Instructions|8926,8933|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|Discharge Instructions|8926,8933|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Event|Event|Discharge Instructions|8952,8961|false|false|false|||concerned
Event|Event|Discharge Instructions|8968,8973|false|false|false|||bleed
Finding|Pathologic Function|Discharge Instructions|8968,8973|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body System|Discharge Instructions|8982,8990|false|false|false|C0017189|Gastrointestinal tract structure|GI tract
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8985,8990|false|false|false|C1185740|Tract|tract
Event|Event|Discharge Instructions|8996,9005|false|false|false|||underwent
Event|Event|Discharge Instructions|9016,9025|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|Discharge Instructions|9016,9025|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|Discharge Instructions|9053,9057|true|false|false|||show
Event|Event|Discharge Instructions|9062,9070|true|false|false|||evidence
Finding|Idea or Concept|Discharge Instructions|9062,9070|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|9062,9073|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Discharge Instructions|9075,9083|true|false|false|||bleeding
Finding|Pathologic Function|Discharge Instructions|9075,9083|true|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|Discharge Instructions|9090,9095|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|9090,9095|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|9090,9095|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|9096,9102|false|false|false|||counts
Event|Event|Discharge Instructions|9112,9118|false|false|false|||stable
Finding|Intellectual Product|Discharge Instructions|9112,9118|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|9133,9141|false|false|false|||hospital
Finding|Idea or Concept|Discharge Instructions|9133,9141|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|9152,9162|false|false|false|||discharged
Disorder|Disease or Syndrome|Discharge Instructions|9168,9172|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Discharge Instructions|9168,9172|false|false|false|||plan
Finding|Functional Concept|Discharge Instructions|9168,9172|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Discharge Instructions|9168,9172|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Discharge Instructions|9168,9172|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|Discharge Instructions|9177,9187|false|false|false|||outpatient
Finding|Classification|Discharge Instructions|9177,9187|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|9177,9187|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|Discharge Instructions|9188,9194|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Discharge Instructions|9188,9194|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Discharge Instructions|9188,9197|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Discharge Instructions|9188,9197|false|false|false|C1522577|follow-up|follow up
Event|Event|Discharge Instructions|9195,9197|false|false|false|||up
Event|Event|Discharge Instructions|9211,9222|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|Discharge Instructions|9211,9222|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Discharge Instructions|9211,9222|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9238,9247|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Discharge Instructions|9238,9247|false|false|false|C2707265||Pulmonary
Finding|Finding|Discharge Instructions|9238,9247|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Finding|Discharge Instructions|9238,9256|false|false|false|C0231921;C1547996;C3160731|Diagnostic Service Section ID - Pulmonary Function;Pulmonary function;Pulmonary function (finding)|Pulmonary function
Finding|Intellectual Product|Discharge Instructions|9238,9256|false|false|false|C0231921;C1547996;C3160731|Diagnostic Service Section ID - Pulmonary Function;Pulmonary function;Pulmonary function (finding)|Pulmonary function
Finding|Organ or Tissue Function|Discharge Instructions|9238,9256|false|false|false|C0231921;C1547996;C3160731|Diagnostic Service Section ID - Pulmonary Function;Pulmonary function;Pulmonary function (finding)|Pulmonary function
Event|Event|Discharge Instructions|9248,9256|false|false|false|||function
Finding|Finding|Discharge Instructions|9248,9256|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Discharge Instructions|9248,9256|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Discharge Instructions|9248,9256|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Discharge Instructions|9248,9256|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|Discharge Instructions|9258,9265|false|false|false|||testing
Finding|Functional Concept|Discharge Instructions|9258,9265|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|Discharge Instructions|9258,9265|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Finding|Discharge Instructions|9278,9282|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|9319,9325|false|false|false|||follow
Event|Event|Discharge Instructions|9367,9375|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|9367,9375|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9367,9375|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|9383,9387|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|9383,9387|false|false|false|||care
Finding|Finding|Discharge Instructions|9383,9387|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9383,9387|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9383,9390|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|9421,9430|true|false|false|||questions
Event|Activity|Discharge Instructions|9441,9445|true|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|9441,9445|true|false|false|||care
Finding|Finding|Discharge Instructions|9441,9445|true|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9441,9445|true|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|9474,9482|true|false|false|||hesitate
Event|Event|Discharge Instructions|9487,9490|true|false|false|||ask
Event|Event|Discharge Instructions|9509,9518|false|false|false|||Inpatient
Finding|Idea or Concept|Discharge Instructions|9509,9518|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|Inpatient
Procedure|Health Care Activity|Discharge Instructions|9509,9518|false|false|false|C1555324|inpatient encounter|Inpatient
Event|Activity|Discharge Instructions|9523,9527|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|9523,9527|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|9523,9527|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|9523,9532|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|9523,9532|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|9536,9544|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9545,9557|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9545,9557|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9545,9557|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

