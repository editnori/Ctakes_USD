CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Plastics|Drug|false|false||PLASTICnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Paxil|Drug|false|false||Paxil
null|Paxil|Drug|false|false||Paxilnull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Craniotomy|Procedure|false|false||craniotomynull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - right|Finding|false|false|C0440857|Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Scalp flap|Anatomy|false|false|C1546653;C1534709;C0423756;C0178298;C0496955;C1546781;C0444099;C2240390;C1552823;C1412362;C1961139;C3683798;C0439061;C3263723;C0043251;C0043250;C0181078;C0037297|scalp flapnull|Scalp structure|Anatomy|false|false|C0037297;C0439061;C1412362|scalpnull|ALOX5AP gene|Finding|false|false|C0038925;C0440857;C0036270|flapnull|Surgical Flaps|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955;C1412362;C0037297;C0423756;C0439061;C1546653;C2240390;C1961139;C3683798|flapnull|Split thickness graft of skin (substance)|Drug|false|false|C1123023;C4520765;C0040748;C0332835|split thickness skin graftnull|Split thickness skin graft (procedure)|Procedure|false|false|C0332835;C1123023;C4520765;C0038925;C0036270;C0440857;C0040748|split thickness skin graftnull|Splitting|Finding|false|false|C0440857|splitnull|Thickness of skin|Finding|false|false|C0440857;C1123023;C4520765;C0038925;C0040748|thickness skinnull|Thick|Modifier|false|false||thicknessnull|Skin graft material|Drug|false|false|C1123023;C4520765;C0332835;C0040748;C0440857|skin graftnull|skin graft (physical finding)|Finding|false|false|C1123023;C4520765;C0440857;C0040748;C0332835;C0038925|skin graftnull|Skin Transplantation|Procedure|false|false|C0040748;C1123023;C4520765;C0038925;C0036270;C0332835;C0440857|skin graftnull|Transplanted skin|Anatomy|false|false|C0037297;C1961139;C3683798;C1546781;C0444099;C2240390;C4545112;C0423756;C0178298;C0496955;C0181078;C0439061;C1546653|skin graftnull|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765;C0038925;C0440857;C0332835;C0040748|skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765;C0038925;C0440857;C0332835;C0040748|skinnull|Skin Specimen Source Code|Finding|false|false|C0038925;C0440857;C0040748;C0332835;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0038925;C0440857;C0040748;C0332835;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C2240390;C0181078;C0037297;C4545112;C0423756;C0439061;C1546781;C0444099;C1961139;C3683798;C1546653|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C2240390;C0181078;C0037297;C4545112;C0423756;C0439061;C1546781;C0444099;C1961139;C3683798;C1546653|skinnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0440857;C0332835;C0038925;C1123023;C4520765;C0040748|graftnull|Graft Procedures on the Head|Procedure|false|false|C0332835;C0040748;C1123023;C4520765;C0038925;C0440857|graft
null|Grafting procedure|Procedure|false|false|C0332835;C0040748;C1123023;C4520765;C0038925;C0440857|graftnull|Transplanted tissue|Anatomy|false|false|C1961139;C3683798;C0178298;C0496955;C0439061;C1546781;C0444099;C0037297;C0181074;C1705210;C1546653;C4545112;C2240390;C0181078|graftnull|Wounds and Injuries|Disorder|false|false|C0440857|wound
null|Traumatic Wound|Disorder|false|false|C0440857|wound
null|Traumatic injury|Disorder|false|false|C0440857|woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||VACnull|VAC Regimen (Vincristine-Dactinomycin-Cyclophosphamide)|Procedure|false|false||VAC
null|cyclophosphamide/doxorubicin/vinblastine protocol|Procedure|false|false||VAC
null|cyclophosphamide/dactinomycin/vinblastine protocol|Procedure|false|false||VAC
null|VAC protocol|Procedure|false|false||VACnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Numerous|LabModifier|false|false||multiplenull|null|Time|false|false||priornull|Operative Surgical Procedures|Procedure|false|false||surgeriesnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Chemotherapy Regimen|Procedure|false|false||chemo
null|Chemotherapy|Procedure|false|false||chemonull|Radiation Ionizing Radiotherapy|Procedure|false|false||radiation
null|Radiotherapy Research|Procedure|false|false||radiation
null|Radiation therapy (procedure)|Procedure|false|false||radiationnull|Electromagnetic Radiation|Phenomenon|false|false||radiation
null|Radiation|Phenomenon|false|false||radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Transaction counts and value totals - month|Finding|false|false|C0018670;C0152336|month
null|Precision - month|Finding|false|false|C0018670;C0152336|monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Medical History|Finding|false|false|C0018670;C0152336|history ofnull|History of present illness (finding)|Finding|false|false|C0018670;C0152336|history
null|History of previous events|Finding|false|false|C0018670;C0152336|history
null|Historical aspects qualifier|Finding|false|false|C0018670;C0152336|history
null|Medical History|Finding|false|false|C0018670;C0152336|history
null|Concept History|Finding|false|false|C0018670;C0152336|historynull|History|Subject|false|false||historynull|Pruritus|Finding|false|false|C0018670;C0152336|pruritusnull|sensory perception of itch|Modifier|false|false||pruritusnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0033774;C0876917;C0262926;C1705255;C0019665;C0262512;C2004062;C1561541;C1561542;C0362076;C0262926|head
null|Head|Anatomy|false|false|C0033774;C0876917;C0262926;C1705255;C0019665;C0262512;C2004062;C1561541;C1561542;C0362076;C0262926|headnull|Head Device|Device|false|false||headnull|husband|Subject|false|false||husbandnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Metals|Drug|false|false||metalnull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardware
null|Computer Hardware Device|Device|false|false||hardwarenull|History of surgery|Finding|false|false||prior surgerynull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Metals|Drug|false|false||metalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Bone flap|Anatomy|false|false|C1412362|bone flapnull|Specimen Type - Bone|Finding|true|false|C0038925;C1442209;C0262950|bone
null|null|Finding|true|false|C0038925;C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1412362;C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1412362;C1546560;C1550616|bonenull|ALOX5AP gene|Finding|true|false|C1442209;C0262950;C0038925;C1266913|flapnull|Surgical Flaps|Anatomy|false|false|C1546560;C1550616;C1412362|flapnull|Rotational|Modifier|false|false||rotationalnull|ALOX5AP gene|Finding|false|false|C0038925|flapnull|Surgical Flaps|Anatomy|false|false|C0178298;C0496955;C1546653;C1546781;C0444099;C3263723;C0043251;C0043250;C2240390;C1412362;C1961139;C3683798;C0037297|flapnull|Skin graft material|Drug|false|false|C0332835;C0040748;C1123023;C4520765|skin graftnull|skin graft (physical finding)|Finding|false|false|C0040748;C1123023;C4520765;C0332835;C0038925|skin graftnull|Skin Transplantation|Procedure|false|false|C0040748;C0332835;C1123023;C4520765;C0038925|skin graftnull|Transplanted skin|Anatomy|false|false|C2240390;C1546653;C0037297;C3263723;C0043251;C0043250;C1546781;C0444099;C1961139;C3683798;C0178298;C0496955;C0181078|skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0332835;C0038925;C1123023;C4520765;C0040748|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C0332835;C0038925;C1123023;C4520765;C0040748|skinnull|Skin Specimen Source Code|Finding|false|false|C0038925;C0332835;C0040748;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0038925;C0332835;C0040748;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C2240390;C1961139;C3683798;C1546653;C0178298;C0496955;C1546781;C0444099;C0037297;C0181078|skin
null|Skin|Anatomy|false|false|C2240390;C1961139;C3683798;C1546653;C0178298;C0496955;C1546781;C0444099;C0037297;C0181078|skinnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0038925;C0040748;C1123023;C4520765;C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C1123023;C4520765;C0040748;C0332835;C0038925|graft
null|Grafting procedure|Procedure|false|false|C1123023;C4520765;C0040748;C0332835;C0038925|graftnull|Transplanted tissue|Anatomy|false|false|C0178298;C0496955;C0181078;C1546781;C0444099;C0181074;C1705210;C3263723;C0043251;C0043250;C1961139;C3683798;C1546653;C2240390;C0037297|graftnull|coverage - HL7PublishingDomain|Finding|false|false||coverage
null|null|Finding|false|false||coverage
null|coverage - financial contract|Finding|false|false||coveragenull|Wounds and Injuries|Disorder|false|false|C0038925;C0040748;C0332835|wound
null|Traumatic Wound|Disorder|false|false|C0038925;C0040748;C0332835|wound
null|Traumatic injury|Disorder|false|false|C0038925;C0040748;C0332835|woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Parietal|Modifier|false|false||parietalnull|Anaplastic astrocytoma|Disorder|false|false||anaplastic astrocytomanull|Undifferentiated|Modifier|false|false||anaplasticnull|Astrocytoma|Disorder|false|false||astrocytomanull|Craniotomy|Procedure|false|false||Craniotomynull|Radiation therapy (procedure)|Procedure|false|false||irradiationnull|Irradiation (physical force)|Phenomenon|false|false||irradiation
null|Radiation|Phenomenon|false|false||irradiationnull|cGy|LabModifier|false|false||cGynull|event cycle|Time|false|false||cyclesnull|Temodar|Drug|false|false||Temodar
null|Temodar|Drug|false|false||Temodarnull|Craniotomy|Procedure|false|false||craniotomynull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Revision procedure|Procedure|false|false||revision
null|Surgical revision|Procedure|false|false||revisionnull|Revision|Time|false|false||revisionnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|Accutane|Drug|false|false||Accutane
null|Accutane|Drug|false|false||Accutanenull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Disease|Disorder|false|false||diseasenull|Tubal Ligation|Procedure|false|false||tubal ligationnull|Ligation|Procedure|false|false||ligationnull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Acute bronchitis|Disorder|false|false||bronchitis
null|Bronchitis|Disorder|false|false||bronchitisnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Seizures|Finding|false|false||seizuresnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Apyrexial|Finding|false|false||Afebrilenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Table Cell Horizontal Align - right|Finding|false|false|C0036270|Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Scalp structure|Anatomy|false|false|C0332803;C1552823;C0184898|scalpnull|Surgical wound|Disorder|false|false|C2338258;C0036270|incisionnull|Surgical incisions|Procedure|false|false|C2338258;C0036270|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Cleaning (activity)|Event|false|false||cleannull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Table Cell Horizontal Align - right|Finding|false|false|C1515974|Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C1552823|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Body Substance Discharge|Finding|true|false||drainage
null|Body Fluid Discharge|Finding|true|false||drainagenull|Drainage procedure|Procedure|true|false||drainagenull|Hemorrhage|Finding|true|false||bleedingnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Plastic surgery service|Entity|false|false||plastic surgery servicenull|Plastic Surgical Procedures|Procedure|false|false||plastic surgerynull|Plastic Surgery Specialty|Title|false|false||plastic surgerynull|Plastics|Drug|false|false||plasticnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|ALOX5AP gene|Finding|false|false|C0038925|flapnull|Surgical Flaps|Anatomy|false|false|C1412362;C1546781;C0444099;C0037297;C2240390;C0178298;C0496955|flapnull|Skin graft material|Drug|false|false|C0040748;C0332835;C1123023;C4520765|skin graftnull|skin graft (physical finding)|Finding|false|false|C1123023;C4520765;C0332835;C0038925;C0040748|skin graftnull|Skin Transplantation|Procedure|false|false|C0038925;C0332835;C1123023;C4520765;C0040748;C0036270|skin graftnull|Transplanted skin|Anatomy|false|false|C1961139;C3683798;C4048801;C0181078;C0178298;C0496955;C1546781;C0444099;C0037297;C2240390;C1546653;C1861101|skin graftnull|Skin and subcutaneous tissue disorders|Disorder|false|false|C0040748;C1123023;C4520765;C0332835;C0038925|skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0040748;C1123023;C4520765;C0332835;C0038925|skinnull|Skin Specimen Source Code|Finding|false|false|C0332835;C0038925;C1123023;C4520765;C0040748|skin
null|Skin Specimen|Finding|false|false|C0332835;C0038925;C1123023;C4520765;C0040748|skinnull|Skin, Human|Anatomy|false|false|C2240390;C1961139;C3683798;C1546653;C1546781;C0444099;C0037297;C0178298;C0496955;C0181078|skin
null|Skin|Anatomy|false|false|C2240390;C1961139;C3683798;C1546653;C1546781;C0444099;C0037297;C0178298;C0496955;C0181078|skinnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C1123023;C4520765;C0332835;C0040748|graftnull|Graft Procedures on the Head|Procedure|false|false|C1123023;C4520765;C0040748;C0332835|graft
null|Grafting procedure|Procedure|false|false|C1123023;C4520765;C0040748;C0332835|graftnull|Transplanted tissue|Anatomy|false|false|C1546781;C0444099;C2240390;C0037297;C1546653;C0181078;C1861101;C4048801;C0181074;C1705210;C0178298;C0496955;C1961139;C3683798|graftnull|Scalp defect|Disorder|false|false|C0040748;C0332835;C0036270|scalp defectnull|Scalp structure|Anatomy|false|false|C1861101;C1457869;C4048801;C0037297|scalpnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|false|false|C0036270;C0332835;C0040748|defectnull|Defect|Finding|false|false|C0036270|defectnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Pain Relief brand of acetaminophen|Drug|false|false||pain relief
null|Pain Relief brand of acetaminophen|Drug|false|false||pain reliefnull|Pain relief|Procedure|false|false||pain reliefnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Cardiovascular system|Anatomy|false|false||cardiovascular
null|Cardiovascular|Anatomy|false|false||cardiovascularnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Pulmonary (intended site)|Finding|false|false|C0024109|Pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268|Pulmonarynull|null|Attribute|false|false|C0024109|Pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||Pulmonarynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C4522268;C2707265|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Oral intake|Finding|false|false|C0226896|oral intakenull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C2137071;C1512806;C1527415;C4521986;C4521161;C3251814|oralnull|Oral|Modifier|false|false||oralnull|Intake|Finding|false|false|C0226896|intakenull|Measurement of fluid intake|Procedure|false|false|C0226896|intake
null|Intake (treatment)|Procedure|false|false|C0226896|intakenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Appropriate|Modifier|false|false||appropriatenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Intestines|Anatomy|false|false||bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Defecation|Finding|false|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementnull|Measuring intake and output|Procedure|false|false||Intake and outputnull|Intake|Finding|false|false||Intakenull|Measurement of fluid intake|Procedure|false|false||Intake
null|Intake (treatment)|Procedure|false|false||Intakenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|On IV|Finding|false|false||on IVnull|cefazolin|Drug|false|false||cefazolin
null|cefazolin|Drug|false|false||cefazolinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|cefadroxil|Drug|false|false||cefadroxil
null|cefadroxil|Drug|false|false||cefadroxilnull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Prophylactic treatment|Procedure|false|false||Prophylaxisnull|prevention & control|Modifier|false|false||Prophylaxisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|subcutaneous heparin|Drug|false|false||subcutaneous heparin
null|subcutaneous heparin|Drug|false|false||subcutaneous heparinnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Ambulate|Finding|false|false||ambulatenull|Early|Time|false|false||earlynull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Urination|Finding|false|false||voiding
null|Voids|Finding|false|false||voidingnull|Helping Behavior|Finding|true|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Scalp structure|Anatomy|false|false|C1546653;C1961139;C3683798|scalpnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0036270;C1515974;C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C0332835;C0036270;C1515974|graft
null|Grafting procedure|Procedure|false|false|C0332835;C0036270;C1515974|graftnull|Transplanted tissue|Anatomy|false|false|C1961139;C3683798;C0181074;C1705210;C1546653|graftnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546653;C1961139;C3683798;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Cleaning (activity)|Event|false|false||cleannull|Pink color|Modifier|false|false||pinknull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Entity|Entity|false|false||thingnull|Donor graft|Drug|false|false|C1515974;C0332835|graft donornull|Graft Dosage Form|Drug|false|false|C1444716;C0332835|graft
null|Graft material|Drug|false|false|C1444716;C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C1444716;C1515974;C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C1444716;C0332835;C1515974|graft
null|Grafting procedure|Procedure|false|false|C1444716;C0332835;C1515974|graftnull|Transplanted tissue|Anatomy|false|false|C1546778;C0730393;C1546653;C1961139;C3683798;C0181074;C1705210|graftnull|Donor site|Anatomy|false|false|C1546653;C1961139;C3683798;C0181074;C1705210;C1546778|donor sitenull|null|Attribute|false|false|C1515974|donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false|C0332835;C1444716;C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0730393;C3263710;C1546653;C1961139;C3683798;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Original|Modifier|false|false||originalnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|Ability to dress|Finding|false|false||dressing
null|null|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Pentasa|Drug|false|false||Pentasa
null|Pentasa|Drug|false|false||Pentasanull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|zolpidem|Drug|false|false||zolpidem
null|zolpidem|Drug|false|false||zolpidemnull|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl er
null|Venlafaxine Hydrochloride ER|Drug|false|false||venlafaxine hcl ernull|venlafaxine hydrochloride|Drug|false|false||venlafaxine hcl
null|venlafaxine hydrochloride|Drug|false|false||venlafaxine hclnull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|Flinders medical centre-7 marker|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hcl
null|hydrochloride|Drug|false|false||hclnull|Hairy Cell Leukemia|Disorder|false|false||hclnull|promethazine|Drug|false|false||promethazine
null|promethazine|Drug|false|false||promethazinenull|Keflex|Drug|false|false||keflex
null|Keflex|Drug|false|false||keflexnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprine
null|azathioprine|Drug|false|false||azathioprinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|dicyclomine|Drug|false|false||dicyclomine
null|dicyclomine|Drug|false|false||dicyclominenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C1720374;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C1720374;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Every eight hours|Time|false|false||Q8Hnull|Every - dosing instruction fragment|Finding|false|false|C0524463;C1325531|everynull|Every (qualifier)|Modifier|false|false||everynull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|fluticasone / salmeterol|Drug|false|false||fluticasone-salmeterolnull|fluticasone|Drug|false|false||fluticasone
null|fluticasone|Drug|false|false||fluticasonenull|salmeterol|Drug|false|false||salmeterol
null|salmeterol|Drug|false|false||salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C0993608;C1550509;C0034789|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329;C1556138|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C4035627;C0993608;C0004048;C0205535;C1561538;C1561539;C4546282;C1550509;C1332410|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false|C1556138|Inhalation
null|Inspiration (function)|Finding|false|false|C1556138|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C1556138|BIDnull|BID gene|Finding|false|false|C1556138|BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false|C1556138|2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false|C1556138|day
null|Precision - day|Finding|false|false|C1556138|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|mesalamine|Drug|false|false||mesalamine
null|mesalamine|Drug|false|false||mesalaminenull|Extended Release Oral Capsule|Drug|false|false|C0524463;C1325531|Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0231448;C5781021;C0006935;C0991505|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0231448;C5781021;C0006935;C0991505|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false|C0524463;C1325531|Extended
null|Extension|Finding|false|false|C0524463;C1325531|Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Extended Release Oral Capsule|Drug|false|false|C0524463;C1325531|Capsule, Extended Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0231448;C5781021;C0991505;C0006935;C5975557;C4264481;C1561538;C1561539|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0231448;C5781021;C0991505;C0006935;C5975557;C4264481;C1561538;C1561539|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Extended (finding)|Finding|false|false|C0524463;C1325531|Extended
null|Extension|Finding|false|false|C0524463;C1325531|Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Four times daily|Time|false|false||QIDnull|4 times|Finding|false|false|C0524463;C1325531|4 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false|C0524463;C1325531|timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false|C0524463;C1325531|day
null|Precision - day|Finding|false|false|C0524463;C1325531|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|topiramate|Drug|false|false||topiramate
null|topiramate|Drug|false|false||topiramatenull|Topiramate measurement|Procedure|false|false||topiramatenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|venlafaxine|Drug|false|false||venlafaxine
null|venlafaxine|Drug|false|false||venlafaxinenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false|C0524463;C1325531|Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C1707871;C0694878;C0015306;C1283071;C0391871;C1337463;C0030685;C0680255;C1963578;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C1707871;C0694878;C0015306;C1283071;C0391871;C1337463;C0030685;C0680255;C1963578;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false|C0524463;C1325531|Extnull|EXT1 wt Allele|Finding|false|false|C0524463;C1325531|Ext
null|EXT1 gene|Finding|false|false|C0524463;C1325531|Extnull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|CAPSULE, EXT RELEASE 24 HR|Drug|false|false|C0524463;C1325531|Capsule, Ext Release 24 hrnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C1707871;C0694878;C1337463;C0006935;C0015306|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0030685;C0680255;C1963578;C1283071;C0391871;C1707871;C0694878;C1337463;C0006935;C0015306|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Hereditary Multiple Exostoses|Disorder|false|false|C0524463;C1325531|Extnull|EXT1 wt Allele|Finding|false|false|C0524463;C1325531|Ext
null|EXT1 gene|Finding|false|false|C0524463;C1325531|Extnull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|propylthiouracil|Drug|false|false||propylthiouracil
null|propylthiouracil|Drug|false|false||propylthiouracilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every eight hours|Time|false|false||Q8Hnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|bacitracin zinc|Drug|false|false||bacitracin zinc
null|bacitracin zinc|Drug|false|false||bacitracin zincnull|bacitracin|Drug|false|false||bacitracin
null|bacitracin|Drug|false|false||bacitracinnull|Zinc Supplements|Drug|false|false||zinc
null|Zinc Drug Class|Drug|false|false||zinc
null|Dietary Zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zinc
null|zinc|Drug|false|false||zincnull|Zinc measurement|Procedure|false|false||zincnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Ointments|Drug|false|false||Ointmentnull|APPL1 gene|Finding|false|false||Applnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|refill|Finding|false|false||Refillsnull|cefadroxil|Drug|false|false||cefadroxil
null|cefadroxil|Drug|false|false||cefadroxilnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|7 days|Time|false|false||7 daysnull|day|Time|false|false||daysnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|MAX protein, human|Drug|false|false||Max
null|MAX protein, human|Drug|false|false||Maxnull|Max (cigarettes)|Finding|false|false||Max
null|Oncogene MAX|Finding|false|false||Max
null|MAX gene|Finding|false|false||Maxnull|Maximum|LabModifier|false|false||Maxnull|per day|Time|false|false||/daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|alprazolam|Drug|false|false||alprazolam
null|alprazolam|Drug|false|false||alprazolamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Craniotomy|Procedure|false|false||craniotomynull|Wound status|Finding|false|false||wound Statusnull|null|Attribute|false|false||wound Statusnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Hardware Removal|Procedure|false|false||hardware removalnull|Computer Hardware Device|Device|false|false||hardware
null|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||hardwarenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Splitting|Finding|false|false||splitnull|Thickness of skin|Finding|false|false|C0332835;C1123023;C4520765;C0040748|thickness skinnull|Thick|Modifier|false|false||thicknessnull|Skin graft material|Drug|false|false|C0332835;C1123023;C4520765;C0040748|skin graftnull|skin graft (physical finding)|Finding|false|false|C0040748;C0332835;C1123023;C4520765|skin graftnull|Skin Transplantation|Procedure|false|false|C0332835;C1123023;C4520765;C0040748|skin graftnull|Transplanted skin|Anatomy|false|false|C2240390;C1961139;C3683798;C0870325;C4048755;C2347934;C1947919;C1547755;C1546653;C0423756;C0185125;C0178298;C0496955;C1546781;C0444099;C0181078;C0037297|skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765;C0040748;C0332835|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765;C0040748;C0332835|skinnull|Skin Specimen Source Code|Finding|false|false|C0332835;C1123023;C4520765;C0040748|skin
null|Skin Specimen|Finding|false|false|C0332835;C1123023;C4520765;C0040748|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0185125;C2240390;C0423756;C0178298;C0496955;C0037297;C1546653;C1961139;C3683798;C0870325;C4048755;C2347934;C1947919;C1547755;C0181078|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0185125;C2240390;C0423756;C0178298;C0496955;C0037297;C1546653;C1961139;C3683798;C0870325;C4048755;C2347934;C1947919;C1547755;C0181078|skinnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0040748;C0332835;C1123023;C4520765|graftnull|Graft Procedures on the Head|Procedure|false|false|C0040748;C0332835;C1123023;C4520765|graft
null|Grafting procedure|Procedure|false|false|C0040748;C0332835;C1123023;C4520765|graftnull|Transplanted tissue|Anatomy|false|false|C0037297;C1546781;C0444099;C0181078;C0423756;C0185125;C2240390;C1961139;C3683798;C1546653;C0181074;C1705210;C0178298;C0496955;C0870325;C4048755;C2347934;C1947919;C1547755|graftnull|HL7 Version 2.5 - Application|Finding|false|false|C0036270;C0040748;C1123023;C4520765;C0332835|application
null|Application Document|Finding|false|false|C0036270;C0040748;C1123023;C4520765;C0332835|application
null|Computer Application|Finding|false|false|C0036270;C0040748;C1123023;C4520765;C0332835|application
null|Regulatory Application|Finding|false|false|C0036270;C0040748;C1123023;C4520765;C0332835|application
null|Apply|Finding|false|false|C0036270;C0040748;C1123023;C4520765;C0332835|applicationnull|Application procedure|Procedure|false|false|C0332835;C1123023;C4520765;C1444716;C0040748;C0036270|applicationnull|Application - unit of product usage|LabModifier|false|false||applicationnull|Scalp structure|Anatomy|false|false|C0870325;C4048755;C2347934;C1947919;C1547755;C0185125|scalpnull|Donor site|Anatomy|false|false|C1546778;C0185125|donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false|C1515974;C1444716|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Always - AcknowledgementCondition|Finding|false|false||always
null|All of the Time|Finding|false|false||alwaysnull|Always (frequency)|Time|false|false||alwaysnull|Apply (administration method)|Finding|false|false||apply
null|Apply (instruction)|Finding|false|false||apply
null|null|Finding|false|false||apply
null|Apply|Finding|false|false||applynull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Suction drainage|Procedure|false|false||suctionnull|Location Equipment - Suction|Modifier|false|false||suctionnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Suction drainage|Procedure|false|false||suctionnull|Location Equipment - Suction|Modifier|false|false||suctionnull|Skin graft material|Drug|false|false|C0332835;C1123023;C4520765;C0040748|skin graftnull|skin graft (physical finding)|Finding|false|false|C1515974;C0040748;C1123023;C4520765;C0332835|skin graftnull|Skin Transplantation|Procedure|false|false|C0040748;C1515974;C1123023;C4520765;C0332835|skin graftnull|Transplanted skin|Anatomy|false|false|C1961139;C3683798;C0181074;C1705210;C0037297;C0178298;C0496955;C1546781;C0444099;C1546653;C2240390;C1546778;C0181078|skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765;C0040748;C1515974;C0332835|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765;C0040748;C1515974;C0332835|skinnull|Skin Specimen Source Code|Finding|false|false|C0332835;C0040748;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0332835;C0040748;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546653;C0037297;C2240390;C1961139;C3683798;C0181078;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546653;C0037297;C2240390;C1961139;C3683798;C0181078;C1546781;C0444099|skinnull|Graft Dosage Form|Drug|false|false|C0040748;C1515974;C0332835|graft
null|Graft material|Drug|false|false|C0040748;C1515974;C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0040748;C1123023;C4520765;C0332835;C1515974|graftnull|Graft Procedures on the Head|Procedure|false|false|C0040748;C1515974;C0332835;C1123023;C4520765|graft
null|Grafting procedure|Procedure|false|false|C0040748;C1515974;C0332835;C1123023;C4520765|graftnull|Transplanted tissue|Anatomy|false|false|C1546781;C0444099;C1546653;C1961139;C3683798;C0178298;C0496955;C2240390;C0181074;C1705210;C0181078;C1546778;C0037297|graftnull|null|Finding|false|false|C1515974;C0040748;C0332835|sitenull|Anatomic Site|Anatomy|false|false|C2240390;C1961139;C3683798;C0037297;C1546653;C0178298;C0496955;C0181074;C1705210;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Scalp structure|Anatomy|false|false||scalpnull|Xeroform|Drug|false|false||Xeroform
null|Xeroform|Drug|false|false||Xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|null|Drug|false|false||bacitracin ointmentnull|bacitracin|Drug|false|false||bacitracin
null|bacitracin|Drug|false|false||bacitracinnull|Ointments|Drug|false|false||ointmentnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Warning - AcknowledgementDetailType|Finding|false|false||WARNING
null|Cautionary Warning|Finding|false|false||WARNING
null|System Alert|Finding|false|false||WARNING
null|Warning - Error severity|Finding|false|false||WARNING
null|Warning - EquipmentAlertLevel|Finding|false|false||WARNINGnull|Warning - Alert level|Modifier|false|false||WARNINGnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Skin graft material|Drug|false|false|C0332835;C1123023;C4520765;C0040748|skin graftnull|skin graft (physical finding)|Finding|false|false|C0332835;C1515974;C0040748;C1123023;C4520765|skin graftnull|Skin Transplantation|Procedure|false|false|C0332835;C1515974;C0040748;C1123023;C4520765|skin graftnull|Transplanted skin|Anatomy|false|false|C1546778;C1546653;C1961139;C3683798;C2240390;C1546781;C0444099;C0037297;C0181078;C0178298;C0496955|skin graftnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0332835;C1123023;C4520765;C0040748|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C0332835;C1123023;C4520765;C0040748|skinnull|Skin Specimen Source Code|Finding|false|false|C0332835;C0040748;C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C0332835;C0040748;C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C0181078;C2240390;C1961139;C3683798;C1546778;C0037297;C1546781;C0444099;C1546653|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C0181078;C2240390;C1961139;C3683798;C1546778;C0037297;C1546781;C0444099;C1546653|skinnull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C1515974;C0040748;C0332835;C1123023;C4520765|graftnull|Graft Procedures on the Head|Procedure|false|false|C0040748;C1515974;C0332835;C1123023;C4520765|graft
null|Grafting procedure|Procedure|false|false|C0040748;C1515974;C0332835;C1123023;C4520765|graftnull|Transplanted tissue|Anatomy|false|false|C0178298;C0496955;C0181074;C1705210;C1546781;C0444099;C2240390;C0181078;C0037297;C1546653;C1961139;C3683798;C1546778|graftnull|null|Finding|false|false|C0040748;C0332835;C1515974;C1123023;C4520765|sitenull|Anatomic Site|Anatomy|false|false|C1546653;C2240390;C1961139;C3683798;C0037297;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Free of (attribute)|Finding|false|false||free ofnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Pressure (finding)|Finding|true|false||pressure
null|null|Finding|true|false||pressure
null|Baresthesia|Finding|true|false||pressurenull|null|Phenomenon|true|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Temperature extreme|Phenomenon|false|false||extreme temperaturesnull|Extreme Response|Finding|false|false||extremenull|Extreme|Modifier|false|false||extremenull|Temperature|LabModifier|false|false||temperaturesnull|null|Finding|false|false||covernull|Cover (physical object)|Device|false|false||cover
null|Cover Device|Device|false|false||covernull|Loose|Modifier|false|false||loosenull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C1515974;C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C1515974;C0332835|graft
null|Grafting procedure|Procedure|false|false|C1515974;C0332835|graftnull|Transplanted tissue|Anatomy|false|false|C1961139;C3683798;C0181074;C1705210;C1546778;C1546653|graftnull|null|Finding|false|false|C0332835;C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546653;C1961139;C3683798;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Water running|Procedure|false|false||water runnull|Running water|Phenomenon|false|false||water runnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Does run (finding)|Finding|false|false||run
null|Running (physical activity)|Finding|false|false||run
null|Go Jogging or Running Question|Finding|false|false||run
null|Run action|Finding|false|false||runnull|Rundi language|Entity|false|false||runnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917|head
null|Head|Anatomy|false|false|C0362076;C0876917|headnull|Head Device|Device|false|false||headnull|Scalp structure|Anatomy|false|false||scalpnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0812434;C0684335|necknull|Lower extremity>Thigh|Anatomy|false|false|C1546778;C2681903;C1140091;C1866503|thigh
null|Thigh structure|Anatomy|false|false|C1546778;C2681903;C1140091;C1866503|thighnull|Donor site|Anatomy|false|false|C1546778;C1552822;C2681903;C1140091;C1866503|donor sitenull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false|C0039866;C4299091;C1444716;C1515974|sitenull|Anatomic Site|Anatomy|false|false|C2681903;C1140091;C1866503;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Table Cell Horizontal Align - left|Finding|false|false|C1444716|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C1515974;C1444716;C0039866;C4299091|air
null|AIRN gene|Finding|false|false|C1515974;C1444716;C0039866;C4299091|air
null|AI/RHEUM|Finding|false|false|C1515974;C1444716;C0039866;C4299091|airnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Old|Time|false|false||oldnull|Xeroform|Drug|false|false||xeroform
null|Xeroform|Drug|false|false||xeroformnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Own|Finding|false|false||ownnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|null|Attribute|false|false||donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0332296;C0020311;C1547961;C0332296|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Plastics|Drug|false|false||Plasticnull|Free of (attribute)|Finding|false|false|C1515974|free ofnull|Free of (attribute)|Finding|false|false|C1515974|freenull|Empty (qualifier)|Modifier|false|false||freenull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false|C1515974|waternull|Hydrotherapy|Procedure|false|false|C1515974|waternull|Shower (physical object)|Device|false|false||showernull|Plastics|Drug|false|false||plasticnull|Leave from Employment|Finding|false|false||leavenull|null|Event|false|false||leavenull|Donor site|Anatomy|false|false|C2681903;C1140091;C1866503;C1546778|donor sitenull|null|Attribute|false|false|C1515974|donornull|Participation Type - donor|Subject|false|false||donor
null|Tissue Donors|Subject|false|false||donor
null|Donor person|Subject|false|false||donornull|null|Finding|false|false|C1515974;C1444716|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C3263710;C2681903;C1140091;C1866503|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false|C1444716;C1515974|air
null|AIRN gene|Finding|false|false|C1444716;C1515974|air
null|AI/RHEUM|Finding|false|false|C1444716;C1515974|airnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Decompression Sickness|Disorder|false|false||bendnull|Does bend|Finding|false|false||bendnull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|false|false||liftingnull|Strenuous Exercise|Finding|false|false||strenuous activitynull|Strenuous|Modifier|false|false||strenuousnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Regular|Modifier|false|false||regularnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenol
null|Tylenol Extra Strength|Drug|false|false||Extra Strength Tylenolnull|Strength (attribute)|Finding|false|false||Strengthnull|Pharmaceutical Strength|LabModifier|false|false||Strength
null|Physical Strength|LabModifier|false|false||Strengthnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Mild pain|Finding|false|false||mild pain
null|Neck Pain Score 2|Finding|false|false||mild painnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Packaging Materials|Device|false|false||packaging
null|Drug Packaging|Device|false|false||packagingnull|Packaging|Phenomenon|false|false||packagingnull|Packing (action)|Event|false|false||packagingnull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|Vicodin|Drug|false|false||Vicodin
null|Vicodin|Drug|false|false||Vicodinnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Active ingredient|Drug|false|false||active ingredientnull|Has active ingredient|Modifier|false|false||active ingredientnull|Ingredient|Drug|false|false||ingredientnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|true|false||medsnull|Medications|Finding|true|false||medsnull|Additional|Finding|false|false||additionalnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||tylenol
null|Tylenol|Drug|false|false||tylenolnull|Antibiotics|Drug|false|false||antibioticnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C3844164;C5975557;C4035627|mouth
null|Oral region|Anatomy|false|false|C1527415;C3844164;C5975557;C4035627|mouthnull|2 times per day|Finding|false|false|C0230028;C0226896|2 times per daynull|2 times|Finding|false|false|C0230028;C0226896|2 timesnull|times/day|LabModifier|false|false||times per daynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false|C0230028;C0226896|timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Different|Modifier|false|false||differentnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Have Constipation|Finding|false|false||have constipationnull|Constipation|Finding|false|false||constipationnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Vicodin|Drug|false|false||vicodin
null|Vicodin|Drug|false|false||vicodinnull|hydrocodone|Drug|false|false||hydrocodone
null|hydrocodone|Drug|false|false||hydrocodonenull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Etc.|Finding|false|false||etcnull|Drinking (function)|Finding|false|false||drinking
null|Alcohol consumption|Finding|false|false||drinkingnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Stool Softener|Drug|false|false||stool softenersnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Food|Drug|false|false||foodsnull|Message Waiting Priority - High|Finding|false|false|C1304649|high
null|high - ActExposureLevelCode|Finding|false|false|C1304649|high
null|IPSS Risk Category High|Finding|false|false|C1304649|high
null|IPSS-R Risk Category High|Finding|false|false|C1304649|high
null|High (finding)|Finding|false|false|C1304649|highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|fiber|Drug|false|false|C1304649|fiber
null|Fiber brand of calcium polycarbophil|Drug|false|false|C1304649|fibernull|Tissue fiber|Anatomy|false|false|C3887512;C5200928;C1561958;C4522209;C5202936;C0225326;C1321801|fibernull|Fiber Device|Device|false|false||fibernull|Animal in fiber production|Entity|false|false||fiber
null|Plant fiber|Entity|false|false||fibernull|Pharmaceutical Preparations|Drug|true|false||medicinesnull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Etc.|Finding|false|false||etcnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Stat (do immediately)|Time|false|false||IMMEDIATELYnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Fever with chills|Finding|false|false||fever with chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Physiologic warmth|Finding|false|false|C1515974|warmth
null|Social warmth|Finding|false|false|C1515974|warmthnull|Emotional tenderness|Finding|false|false|C1515974|tenderness
null|Sore to touch|Finding|false|false|C1515974|tendernessnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0684239;C0234233;C0543467;C0587668;C0518610;C0392197|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Unusual|Modifier|false|false||unusualnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false|C2338258|drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0013103;C0184898;C0332803|incisionnull|Large amount|LabModifier|false|false||large amountnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Amount class - Amount|Finding|false|false|C2338258|amountnull|Quantity|LabModifier|false|false||amountnull|Hemorrhage|Finding|false|false|C2338258|bleedingnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C1561574;C0019080;C0184898|incisionnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Severe Extremity Pain|Finding|false|false||Severe pain
null|Severe pain|Finding|false|false||Severe pain
null|Neck Pain Score 6|Finding|false|false||Severe painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false|C2338258|dischargenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0030685;C0332803|incisionnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C2926613|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Else|Finding|false|false||elsenull|Equipment Alert Level - Serious|Finding|false|false||serious
null|Device Alert Level - Serious|Finding|false|false||serious
null|Alert level - Serious|Finding|false|false||seriousnull|Serious|Modifier|false|false||seriousnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Concern|Finding|false|false||concernnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions