CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Low Back Pain|Finding|false|false|C1140621;C0023216|Low back painnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Back Pain with Radiation|Finding|false|false|C1140621;C0023216;C0230442;C0230415|back pain with radiationnull|Back Pain|Finding|false|false|C0230442;C0230415;C1140621;C0023216|back painnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216;C0230442;C0230415|pain
null|Pain|Finding|false|false|C1140621;C0023216;C0230442;C0230415|painnull|null|Attribute|false|false||painnull|Radiation Ionizing Radiotherapy|Procedure|false|false|C0230442;C0230415;C1140621;C0023216|radiation
null|Radiotherapy Research|Procedure|false|false|C0230442;C0230415;C1140621;C0023216|radiation
null|Radiation therapy (procedure)|Procedure|false|false|C0230442;C0230415;C1140621;C0023216|radiationnull|Electromagnetic Radiation|Phenomenon|false|false|C0230442;C0230415;C1140621;C0023216|radiation
null|Radiation|Phenomenon|false|false|C0230442;C0230415;C1140621;C0023216|radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Structure of right lower leg|Anatomy|false|false|C0034519;C0851346;C0004604;C1522449;C1524020;C1524021;C1552823;C1549543;C0030193;C0740363|right leg
null|Right lower extremity|Anatomy|false|false|C0034519;C0851346;C0004604;C1522449;C1524020;C1524021;C1552823;C1549543;C0030193;C0740363|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C1140621;C0023216;C0230442;C0230415|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false|C1549543;C0030193;C0024031;C0740363;C1522449;C1524020;C1524021;C1552823;C0004604;C0034519;C0851346|leg
null|Lower Extremity|Anatomy|false|false|C1549543;C0030193;C0024031;C0740363;C1522449;C1524020;C1524021;C1552823;C0004604;C0034519;C0851346|legnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Decompression - action (qualifier value)|Finding|false|false||DECOMPRESSIONnull|Decompression|Procedure|false|false||DECOMPRESSION
null|Decompressive incision|Procedure|false|false||DECOMPRESSIONnull|external decompression|Phenomenon|false|false||DECOMPRESSIONnull|Fused structure|Finding|false|false||FUSIONnull|Fusion procedure|Procedure|false|false||FUSIONnull|Duraplasty|Procedure|false|false||DURAPLASTYnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Cerebral Aneurysm|Disorder|false|false|C0228174;C0006104|cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0002940;C0162871;C0917996|cerebral
null|Brain|Anatomy|false|false|C0002940;C0162871;C0917996|cerebralnull|Aortic Aneurysm, Abdominal|Disorder|false|false|C0003483;C0000726;C0228174;C0006104|aneurysm, abdominal aorticnull|Aneurysm|Finding|false|false|C0228174;C0006104|aneurysmnull|Abdomen|Anatomy|false|false|C0162871|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Aorta|Anatomy|false|false|C0162871|aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Pallister W syndrome|Disorder|false|false||syndrome wnull|Syndrome|Disorder|false|false||syndromenull|Numerous|LabModifier|false|false||multiplenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Event|Event|false|false|C1690938;C3853547;C0687080;C0016504|eventnull|Bilateral|Modifier|false|false||bilateralnull|LARGE1 wt Allele|Finding|false|false|C1690938;C3853547;C0687080;C0016504|large
null|LARGE1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|largenull|Large|LabModifier|false|false||largenull|Personal Experience Scales|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEs
null|PES1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false|C0441471;C0851145;C5890938;C1416798;C1418467;C0687136|PEs
null|Hindfoot of quadruped|Anatomy|false|false|C0441471;C0851145;C5890938;C1416798;C1418467;C0687136|PEs
null|Paw|Anatomy|false|false|C0441471;C0851145;C5890938;C1416798;C1418467;C0687136|PEs
null|Foot|Anatomy|false|false|C0441471;C0851145;C5890938;C1416798;C1418467;C0687136|PEsnull|Iranian Persian language|Entity|false|false||PEsnull|on warfarin|Procedure|false|false|C1690938;C3853547;C0687080;C0016504|on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|BRCA1 gene mutation|Disorder|false|false||BRCA1 mutationnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||mutationnull|Mutation|Finding|false|false||mutationnull|Malignant neoplasm of breast|Disorder|false|false|C0006141|breast cancer
null|Breast Carcinoma|Disorder|false|false|C0006141|breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0191838;C0496956;C0006826;C0006142;C0678222;C0567499|breastnull|Malignant Neoplasms|Disorder|false|false|C0006141|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Transaction counts and value totals - month|Finding|false|false|C1548802;C0230102;C2939142|month
null|Precision - month|Finding|false|false|C1548802;C0230102;C2939142|monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|right-sided low back pain|Finding|false|false|C0230102;C2939142;C1548802|right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false|C0230102;C2939142;C1548802|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false|C0230102;C2939142;C1548802|lower back painnull|Lower back (surface region)|Anatomy|false|false|C1552823;C2219286;C2598155;C1561541;C1561542;C0004604;C0024031;C1549543;C0030193|lower back
null|Lower back structure|Anatomy|false|false|C1552823;C2219286;C2598155;C1561541;C1561542;C0004604;C0024031;C1549543;C0030193|lower backnull|Body Site Modifier - Lower|Anatomy|false|false|C1561541;C1561542;C1549543;C0030193;C2598155;C2003888;C2219286;C1552823;C0024031;C0004604|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false|C0230102;C2939142;C1548802|back painnull|Administration Method - Pain|Finding|false|false|C1548802;C0230102;C2939142|pain
null|Pain|Finding|false|false|C1548802;C0230102;C2939142|painnull|null|Attribute|false|false|C0230102;C2939142;C1548802|painnull|Radicular pain|Finding|false|false||radicular painnull|Dermatomal|Modifier|false|false||radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in right leg|Finding|false|false|C1140621;C0023216;C0230442;C0230415|right leg painnull|Structure of right lower leg|Anatomy|false|false|C2598155;C0023222;C5848135;C1552823;C1549543;C0030193|right leg
null|Right lower extremity|Anatomy|false|false|C2598155;C0023222;C5848135;C1552823;C1549543;C0030193|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C1140621;C0023216;C0230442;C0230415|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false|C0230442;C0230415;C1140621;C0023216|leg painnull|Leg|Anatomy|false|false|C5848135;C1549543;C0030193;C2598155;C1552823;C0023222|leg
null|Lower Extremity|Anatomy|false|false|C5848135;C1549543;C0030193;C2598155;C1552823;C0023222|legnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216;C0230442;C0230415|pain
null|Pain|Finding|false|false|C1140621;C0023216;C0230442;C0230415|painnull|null|Attribute|false|false|C0230442;C0230415;C1140621;C0023216|painnull|Recent|Time|false|false||recentnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Background|Finding|false|false||backgroundnull|month|Time|false|false||monthsnull|Pain in right leg|Finding|false|false|C1140621;C0023216;C0230442;C0230415|right leg painnull|Structure of right lower leg|Anatomy|false|false|C1552823;C2598155;C1549543;C0030193;C5848135;C0023222|right leg
null|Right lower extremity|Anatomy|false|false|C1552823;C2598155;C1549543;C0030193;C5848135;C0023222|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C0230442;C0230415|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false|C1140621;C0023216;C0230442;C0230415|leg painnull|Leg|Anatomy|false|false|C5848135;C0023222;C1549543;C0030193|leg
null|Lower Extremity|Anatomy|false|false|C5848135;C0023222;C1549543;C0030193|legnull|Administration Method - Pain|Finding|false|false|C0230442;C0230415;C1140621;C0023216|pain
null|Pain|Finding|false|false|C0230442;C0230415;C1140621;C0023216|painnull|null|Attribute|false|false|C0230442;C0230415|painnull|Evidence of (contextual qualifier)|Finding|false|false|C5239664|evidence ofnull|Evidence|Finding|false|false|C5239664|evidencenull|Deep thrombophlebitis|Disorder|true|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|true|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C3887511;C2926618;C0149871;C0151950;C0332120|DVTnull|null|Attribute|true|false|C5239664|DVTnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|right trochanteric bursitis|Disorder|false|false||right trochanteric bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Injection of steroid|Procedure|false|false||steroid injectionnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Right tibia|Anatomy|false|false|C0740426;C1552823;C2598155;C1549543;C0030193|right tibianull|Table Cell Horizontal Align - right|Finding|false|false|C0040184;C0817321|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Tibia pain|Finding|false|false|C0817321;C0040184|tibia painnull|Bone structure of tibia|Anatomy|false|false|C1552823;C0740426;C1549543;C0030193|tibianull|Tibia <Rostellariidae>|Entity|false|false||tibianull|Administration Method - Pain|Finding|false|false|C0040184;C0817321|pain
null|Pain|Finding|false|false|C0040184;C0817321|painnull|null|Attribute|false|false|C0817321|painnull|Varicosity|Disorder|false|false|C0042449|varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0398102;C0042345|veinsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT A
null|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT Anull|Nephrolithiasis|Disorder|false|false||nephrolithiasisnull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920|spine
null|Vertebral column|Anatomy|false|false|C0150920|spinenull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C1621443;C1556138|disc
null|Discontinued|Finding|false|false|C1621443;C1556138|discnull|Disc - Body Part|Anatomy|false|false|C0038999;C0993608;C1696131;C1444662|disc
null|death-inducing signaling complex location|Anatomy|false|false|C0038999;C0993608;C1696131;C1444662|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Swelling|Finding|false|false|C1621443;C1556138|bulgenull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Narrow|Modifier|false|false||narrowing ofnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Spinal Canal|Anatomy|false|false|C0040433;C0010383;C0017589;C0349017|spinal canalnull|Spinal|Modifier|false|false||spinalnull|canal [body parts]|Anatomy|false|false|C0040433;C0010383;C0017589;C0349017|canal
null|Pulp Canals|Anatomy|false|false|C0040433;C0010383;C0017589;C0349017|canalnull|Geographic canal|Entity|false|false||canalnull|Tooth Crowding|Finding|false|false|C0007458;C0037922;C0086881;C1550227|crowding
null|Crowding|Finding|false|false|C0007458;C0037922;C0086881;C1550227|crowdingnull|Malignant neoplasm of cauda equina|Disorder|false|false|C0037922;C0007458;C0086881;C1550227|cauda equinanull|Cauda Equina|Anatomy|false|false|C0040433;C0010383;C0017589;C0349017|cauda equinanull|Glanders|Disorder|false|false|C0037922;C0007458;C0086881;C1550227|equinanull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false|C0042449|Varicose veinsnull|Varicose|Modifier|false|false||Varicosenull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0042345;C0398102|veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEs
null|PES1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false|C1418467;C0687136|PEs
null|Hindfoot of quadruped|Anatomy|false|false|C1418467;C0687136|PEs
null|Paw|Anatomy|false|false|C1418467;C0687136|PEs
null|Foot|Anatomy|false|false|C1418467;C0687136|PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false|C1167408;C3665580|antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false|C1167408;C3665580|antiphospholipid antibodynull|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibodynull|Antibody (immunoassay)|Procedure|false|false|C1167408;C3665580|antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false|C0162595;C4019436;C0039082;C0085278;C4551530;C0003241;C0021027|antibody
null|immunoglobulin complex location|Anatomy|false|false|C0162595;C4019436;C0039082;C0085278;C4551530;C0003241;C0021027|antibodynull|Syndrome|Disorder|false|false|C1167408;C3665580|syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false||A1Cnull|Cerebral Aneurysm|Disorder|false|false|C0228174;C0006104|cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0917996;C0002940|cerebral
null|Brain|Anatomy|false|false|C0917996;C0002940|cerebralnull|Aneurysm|Finding|false|false|C0228174;C0006104|aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|false|false|C0009368;C4071907|colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|false|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0009376|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0750873;C0009376|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|polyps|Disorder|false|false||polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false|C0392905;C1269611;C0022417;C3890599|CMC
null|Capillary malformation (disorder)|Disorder|false|false|C0392905;C1269611;C0022417;C3890599|CMCnull|MCC protocol|Procedure|false|false|C3890599;C0392905;C1269611;C0022417|CMCnull|Circulating Melanoma Cell|Anatomy|false|false|C0065772;C0006845;C0340803;C0575044|CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false|C0392905;C1269611;C0022417|joint arthroplastynull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417;C3890599|jointnull|null|Anatomy|false|false|C0575044;C0006845;C0340803;C0065772;C0003893|joint
null|Joints|Anatomy|false|false|C0575044;C0006845;C0340803;C0065772;C0003893|joint
null|Articular system|Anatomy|false|false|C0575044;C0006845;C0340803;C0065772;C0003893|jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false||arthroplasty
null|Arthroplasty|Procedure|false|false||arthroplasty
null|Reconstruction of joint|Procedure|false|false||arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false|C0085515;C1550244|rotator cuff repairnull|Rotator Cuff|Anatomy|false|false|C0186666;C3668885|rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false|C1550244;C0085515|cuffnull|Cuff - body part|Anatomy|false|false|C3668885;C0186666|cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Excision|Procedure|false|false||excision
null|removal technique|Procedure|false|false||excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false|C0582802|digitnull|Digit structure|Anatomy|false|false|C4761764|digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false|C4482304;C0030288;C0687028;C1550227;C0030274|pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic duct
null|Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic ductnull|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreaticnull|Pancreas|Anatomy|false|false|C0030292;C0153461|pancreaticnull|Duct (organ) structure|Anatomy|false|false|C0153461|duct
null|canal [body parts]|Anatomy|false|false|C0153461|ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false|C4482304;C0030288|explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|ovarian neoplasm|Disorder|false|false|C0205065|OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false|C0205065|OVARIAN CANCERnull|Ovarian|Anatomy|false|false|C0006826;C0919267;C1140680|OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false|C0205065|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Malignant neoplasm of brain|Disorder|false|false|C4266577;C0006104|BRAIN CANCER
null|Brain Neoplasms|Disorder|false|false|C4266577;C0006104|BRAIN CANCERnull|Brain Diseases|Disorder|false|false|C4266577;C0006104|BRAINnull|Head>Brain|Anatomy|false|false|C0006111;C0006826;C0153633;C0006118|BRAIN
null|Brain|Anatomy|false|false|C0006111;C0006826;C0153633;C0006118|BRAINnull|Malignant Neoplasms|Disorder|false|false|C4266577;C0006104|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Platinum-Group Metal|Drug|false|false|C0205065|PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false|C0205065|PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false|C0205065|PGMnull|phosphoglycerate mutase activity|Finding|false|false|C0205065|PGMnull|ovarian neoplasm|Disorder|false|false|C0205065|OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false|C0205065|OVARIAN CANCERnull|Ovarian|Anatomy|false|false|C0006826;C1150365;C0919267;C1140680;C3815181;C0031653|OVARIANnull|Malignant Neoplasms|Disorder|false|false|C0205065|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Aunt|Subject|false|false||Auntnull|ovarian neoplasm|Disorder|false|true|C0205065|OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|true|C0205065|OVARIAN CANCERnull|Ovarian|Anatomy|false|false|C0006826;C0919267;C1140680|OVARIANnull|Malignant Neoplasms|Disorder|false|true|C0205065|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|true||CANCERnull|Paternal aunt|Subject|false|false||paternal auntnull|Paternal Relative|Subject|false|false||paternalnull|Paternal (qualifier value)|Modifier|false|false||paternalnull|Aunt|Subject|false|false||auntnull|Endometrial Carcinoma|Disorder|false|false||ENDOMETRIAL CANCER
null|Malignant neoplasm of endometrium|Disorder|false|false||ENDOMETRIAL CANCERnull|Endometrial|Modifier|false|false||ENDOMETRIALnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|STAT5A protein, human|Drug|false|false|C0033572;C4266527|MGF
null|IGF1 protein, human|Drug|false|false|C0033572;C4266527|MGF
null|IGF1 protein, human|Drug|false|false|C0033572;C4266527|MGF
null|STAT5A protein, human|Drug|false|false|C0033572;C4266527|MGF
null|Kit Ligand, human|Drug|false|false|C0033572;C4266527|MGF
null|Kit Ligand, human|Drug|false|false|C0033572;C4266527|MGFnull|STAT5A wt Allele|Finding|false|false|C0033572;C4266527|MGF
null|KITLG gene|Finding|false|false|C0033572;C4266527|MGF
null|STAT5A gene|Finding|false|false|C0033572;C4266527|MGF
null|KITLG wt Allele|Finding|false|false|C0033572;C4266527|MGFnull|Malignant neoplasm of prostate|Disorder|false|false|C0033572;C4266527|PROSTATE CANCER
null|Prostate carcinoma|Disorder|false|false|C0033572;C4266527|PROSTATE CANCERnull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false|C0033572;C4266527|PROSTATE
null|Prostatic Diseases|Disorder|false|false|C0033572;C4266527|PROSTATE
null|Carcinoma in situ of prostate|Disorder|false|false|C0033572;C4266527|PROSTATE
null|Benign neoplasm of prostate|Disorder|false|false|C0033572;C4266527|PROSTATEnull|Structure of prostate (body structure)|Anatomy|false|false|C1366394;C3887684;C3712803;C0006826;C0376358;C0600139;C1335875;C1705050;C1704887;C1366480;C0496923;C0154088;C0033575;C0154009|PROSTATE
null|Prostate|Anatomy|false|false|C1366394;C3887684;C3712803;C0006826;C0376358;C0600139;C1335875;C1705050;C1704887;C1366480;C0496923;C0154088;C0033575;C0154009|PROSTATEnull|Malignant Neoplasms|Disorder|false|false|C0033572;C4266527|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Malignant neoplasm of kidney|Disorder|false|false|C0227665;C0022646|KIDNEY CANCER
null|Renal carcinoma|Disorder|false|false|C0227665;C0022646|KIDNEY CANCERnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|KIDNEY
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|KIDNEYnull|Kidney problem|Finding|false|false|C0227665;C0022646|KIDNEYnull|examination of kidney|Procedure|false|false|C0227665;C0022646|KIDNEY
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|KIDNEYnull|Kidney|Anatomy|false|false|C0006826;C0496927;C0496892;C4554465;C0869841;C0740457;C1378703;C0812426|KIDNEY
null|Both kidneys|Anatomy|false|false|C0006826;C0496927;C0496892;C4554465;C0869841;C0740457;C1378703;C0812426|KIDNEYnull|Malignant Neoplasms|Disorder|false|false|C0227665;C0022646|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Kidney Failure|Disorder|false|false|C0022646|RENAL FAILUREnull|Urologic Diseases|Disorder|false|false|C0022646|RENALnull|Kidney|Anatomy|false|false|C0035078;C0680095;C0231174;C5200924;C0042075|RENALnull|Failure (biologic function)|Finding|false|false|C0022646|FAILURE
null|Failure|Finding|false|false|C0022646|FAILURE
null|Personal failure|Finding|false|false|C0022646|FAILUREnull|Congestive|Modifier|false|false||CONGESTIVEnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|HEART
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|HEARTnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Diabetes Mellitus|Disorder|false|false||DIABETES MELLITUSnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||DIABETES
null|Diabetes|Disorder|false|false||DIABETES
null|Diabetes Mellitus|Disorder|false|false||DIABETESnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Alcohol abuse|Disorder|false|false||ALCOHOL ABUSEnull|Alcohols|Drug|false|false||ALCOHOL
null|Alcohols|Drug|false|false||ALCOHOL
null|ethanol|Drug|false|false||ALCOHOL
null|ethanol|Drug|false|false||ALCOHOLnull|Alcohol - Recreational Drug Use Code|Finding|false|false||ALCOHOLnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Sister - courtesy title|Finding|false|false||Sister
null|Relationship - Sister|Finding|false|false||Sisternull|Sister|Subject|false|false||Sisternull|ovarian neoplasm|Disorder|false|false|C0205065|OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false|C0205065|OVARIAN CANCERnull|Ovarian|Anatomy|false|false|C0006826;C0919267;C1140680|OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false|C0205065|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|true||age
null|Glycation End Products, Advanced|Drug|false|true||agenull|null|Attribute|false|true||agenull|Age|Subject|false|false||agenull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Throat cancer|Disorder|false|false|C0230069;C3665375;C0031354|THROAT CANCERnull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|THROATnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|THROAT
null|null|Finding|false|false|C0230069;C3665375;C0031354|THROATnull|Throat|Anatomy|false|false|C0740339;C1550663;C1547926;C0006826;C1950455|THROAT
null|Anterior portion of neck|Anatomy|false|false|C0740339;C1550663;C1547926;C0006826;C1950455|THROAT
null|Pharyngeal structure|Anatomy|false|false|C0740339;C1550663;C1547926;C0006826;C1950455|THROATnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false|C0230069;C3665375;C0031354|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Sister - courtesy title|Finding|false|false|C0006141|Sister
null|Relationship - Sister|Finding|false|false|C0006141|Sisternull|Sister|Subject|false|false||Sisternull|BRCA1 gene mutation|Disorder|false|false||BRCA1 MUTATIONnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||MUTATIONnull|Mutation|Finding|false|false||MUTATIONnull|Malignant neoplasm of breast|Disorder|false|true|C0006141|BREAST CANCER
null|Breast Carcinoma|Disorder|false|true|C0006141|BREAST CANCERnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|BREASTnull|Breast problem|Finding|false|false|C0006141|BREASTnull|Procedures on breast|Procedure|false|false|C0006141|BREASTnull|Breast|Anatomy|false|false|C0191838;C0567499;C0006142;C0678222;C0496956;C0006826;C1546515;C1704647|BREASTnull|Malignant Neoplasms|Disorder|false|false|C0006141|CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Daughter|Subject|false|false||Daughternull|Abnormal cervical smear|Finding|false|true|C3496568|ABNORMAL PAP SMEARnull|Observation Interpretation - Abnormal|Finding|false|false||ABNORMAL
null|Abnormal|Finding|false|false||ABNORMALnull|Pap smear|Procedure|false|false|C3496568|PAP SMEAR
null|Papanicolaou Test|Procedure|false|false|C3496568|PAP SMEARnull|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false|C3496568|PAP
null|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false|C3496568|PAP
null|ACPP protein, human|Drug|false|false|C3496568|PAP
null|ACPP protein, human|Drug|false|false|C3496568|PAPnull|null|Finding|false|false|C3496568|PAP
null|PAPOLA wt Allele|Finding|false|false|C3496568|PAP
null|PDAP1 gene|Finding|false|false|C3496568|PAP
null|TUSC2 wt Allele|Finding|false|false|C3496568|PAP
null|ASAP1 wt Allele|Finding|false|false|C3496568|PAP
null|ACP3 wt Allele|Finding|false|false|C3496568|PAP
null|Pulmonary artery pressure|Finding|false|false|C3496568|PAP
null|TUSC2 gene|Finding|false|false|C3496568|PAP
null|ASAP2 gene|Finding|false|false|C3496568|PAP
null|ASAP1 gene|Finding|false|false|C3496568|PAP
null|REG3A gene|Finding|false|false|C3496568|PAP
null|PITUITARY ADENOMA PREDISPOSITION|Finding|false|false|C3496568|PAP
null|PAPOLA gene|Finding|false|false|C3496568|PAP
null|ACP3 gene|Finding|false|false|C3496568|PAP
null|REG3A wt Allele|Finding|false|false|C3496568|PAP
null|MRPS30 gene|Finding|false|false|C3496568|PAPnull|pars anterior of the paramedian lobule|Anatomy|false|false|C0444186;C1740167;C0760170;C0079104;C3541459;C3872789;C0476427;C1422804;C3889402;C1423108;C1863340;C3538851;C1418410;C1705531;C1705530;C1413945;C1538823;C1367456;C0428642;C1413944;C1705529;C1424700;C2266415|PAPnull|Papiamento language|Entity|false|false||PAPnull|Smearing technique|Finding|false|false|C3496568|SMEARnull|Smear test|Procedure|false|false|C3496568|SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|Substance Abuse Problems|Disorder|false|false||SUBSTANCE ABUSE
null|Harmful pattern of substance use|Disorder|false|false||SUBSTANCE ABUSEnull|Substance|Drug|false|false||SUBSTANCEnull|administrative information regarding test substance|Finding|false|false||SUBSTANCEnull|null|Attribute|false|false||SUBSTANCEnull|Substance (attribute)|Modifier|false|false||SUBSTANCEnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|SON gene|Finding|false|false||Sonnull|Son (person)|Subject|false|false||Sonnull|Songhay Languages|Entity|false|false||Sonnull|Substance Abuse Problems|Disorder|false|false||SUBSTANCE ABUSE
null|Harmful pattern of substance use|Disorder|false|false||SUBSTANCE ABUSEnull|Substance|Drug|false|false||SUBSTANCEnull|administrative information regarding test substance|Finding|false|false||SUBSTANCEnull|null|Attribute|false|false||SUBSTANCEnull|Substance (attribute)|Modifier|false|false||SUBSTANCEnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Heroin overdose|Disorder|false|false||heroin overdosenull|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroinnull|Poisoning by heroin|Disorder|false|false||heroinnull|Drug Overdose|Disorder|false|false||overdosenull|Event Qualification - Overdose|Finding|false|false||overdose
null|Overdose|Finding|false|false||overdosenull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Weepiness|Finding|false|false||Tearfulnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false|C1140621;C0023216|leg painnull|Leg|Anatomy|false|false|C0023222;C1549543;C0030193|leg
null|Lower Extremity|Anatomy|false|false|C0023222;C1549543;C0030193|legnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216|pain
null|Pain|Finding|false|false|C1140621;C0023216|painnull|null|Attribute|false|false||painnull|Spasm|Finding|false|false||spasmsnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0741025|Chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|Chestnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0496956;C0191838;C5575035;C0567499;C0205249;C0184898|breastnull|Surgical incisions|Procedure|false|false|C0006141|incisionsnull|Well (answer to question)|Finding|false|false|C0006141|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Healed|Finding|false|false|C0006141|healednull|Axilla|Anatomy|false|false|C0543467;C0587668|axillanull|Operative Surgical Procedures|Procedure|false|false|C0004454|surgical
null|Surgical service|Procedure|false|false|C0004454|surgicalnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false|C0230415;C0023216|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Right lower extremity|Anatomy|false|false|C1552823;C5575035;C2003888|right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false|C0230415;C0023216;C0015385|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false|C2003888;C1552823;C5575035|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0023216;C0015385;C0230415|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false|C1552823;C2003888|extremitynull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Movement|Finding|false|false||movementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||Swelling
null|Edema|Finding|false|false||Swellingnull|Palpable|Modifier|false|false||Palpablenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skinnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Varicosity|Disorder|false|false|C0023216;C0278454;C0015385;C0042449|varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false|C0023216;C0278454;C0015385;C0042449|veinsnull|Veins|Anatomy|false|false|C0042345;C0398102|veinsnull|Lower Extremity|Anatomy|false|false|C0398102;C2003888;C0042345|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0023216;C0278454;C0015385|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C0398102;C0042345;C2003888|extremities
null|Limb structure|Anatomy|false|false|C0398102;C0042345;C2003888|extremitiesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Medullary sponge kidney|Disorder|false|false||MSK
null|Medullary sponge kidney|Disorder|false|false||MSKnull|SIK1 gene|Finding|false|false||MSKnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|SI joint|Anatomy|false|false|C0684239;C0234233;C0240094;C0575044|SI Jointnull|Joint tenderness|Finding|false|false|C5453012;C0392905;C1269611;C0022417|Joint tendernessnull|Joint problem|Finding|false|false|C5453012;C0392905;C1269611;C0022417|Jointnull|null|Anatomy|false|false|C0684239;C0234233;C0575044;C0240094|Joint
null|Joints|Anatomy|false|false|C0684239;C0234233;C0575044;C0240094|Joint
null|Articular system|Anatomy|false|false|C0684239;C0234233;C0575044;C0240094|Jointnull|Joint Device|Device|false|false||Jointnull|Emotional tenderness|Finding|false|false|C5453012;C0392905;C1269611;C0022417|tenderness
null|Sore to touch|Finding|false|false|C5453012;C0392905;C1269611;C0022417|tendernessnull|Radicular pain|Finding|false|false||Radicular painnull|Dermatomal|Modifier|false|false||Radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Hip flexion|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip flexionnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1292890;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2237371|hip
null|Hip structure|Anatomy|false|false|C1292890;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2237371|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1292890;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2237371|hip
null|Bone structure of ischium|Anatomy|false|false|C1292890;C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C2237371|hipnull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Knee flexion|Finding|false|false|C1963703;C0022742;C4299094;C0022745|knee flexionnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C0231452;C0562271;C0240114|knee
null|Knee|Anatomy|false|false|C0231452;C0562271;C0240114|knee
null|Lower extremity>Knee|Anatomy|false|false|C0231452;C0562271;C0240114|knee
null|Knee joint|Anatomy|false|false|C0231452;C0562271;C0240114|kneenull|null|Finding|false|false|C1963703;C0022742;C4299094;C0022745|flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Foot problem|Finding|false|false|C0442036;C0230463;C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980|foot
null|Foot|Anatomy|false|false|C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Plantar (qualifier value)|Anatomy|false|false|C0555980;C2229507;C0036658;C0542538|plantar
null|Sole of Foot|Anatomy|false|false|C0555980;C2229507;C0036658;C0542538|plantarnull|Observation of Sensation|Finding|false|false|C0442036;C0230463|sensation
null|Sensory perception|Finding|false|false|C0442036;C0230463|sensationnull|sensory exam|Procedure|false|false|C0442036;C0230463|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Tact|Drug|false|false||tact
null|Tact|Drug|false|false||tact
null|Tact|Drug|false|false||tact
null|bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|Drug|false|false||tactnull|Ortho-|Finding|false|false|C2752558;C0037949|Orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||Orthonull|Spine Problem|Finding|false|false|C2752558;C0037949|Spinenull|Neuron spine|Anatomy|false|false|C0150920;C0812371|Spine
null|Vertebral column|Anatomy|false|false|C0150920;C0812371|Spinenull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|null|Attribute|false|false||resp effortnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||respnull|Respiratory rate|Attribute|false|false||respnull|Exertion|Finding|false|false||effortnull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|LAT protein, human|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|LAT protein, human|Drug|false|false||latnull|LAT gene|Finding|false|false|C0446516;C1140618;C1269078|lat
null|ORC3 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|lat
null|ORC3 gene|Finding|false|false|C0446516;C1140618;C1269078|lat
null|SPNS1 gene|Finding|false|false|C0446516;C1140618;C1269078|latnull|Latin Language|Entity|false|false||latnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044;C1705279;C1335085;C1425844;C2240043|arm
null|null|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044;C1705279;C1335085;C1425844;C2240043|arm
null|Upper Extremity|Anatomy|false|false|C1522541;C5400986;C4761640;C3495676;C1824218;C3715044;C1705279;C1335085;C1425844;C2240043|armnull|Thumb structure|Anatomy|false|false||thumbnull|Middle|Modifier|false|false||midnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Multiple Epiphyseal Dysplasia|Disorder|false|false|C0446516;C1140618;C1269078|mednull|Master of Education|Finding|false|false|C0446516;C1140618;C1269078|med
null|COMP wt Allele|Finding|false|false|C0446516;C1140618;C1269078|med
null|COL9A3 gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|SCN8A wt Allele|Finding|false|false|C0446516;C1140618;C1269078|med
null|COL9A2 gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|COMP gene|Finding|false|false|C0446516;C1140618;C1269078|med
null|SCN8A gene|Finding|false|false|C0446516;C1140618;C1269078|mednull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C1522541;C5400986;C4761640;C1824218;C3715044;C3495676;C0026760|arm
null|null|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C1522541;C5400986;C4761640;C1824218;C3715044;C3495676;C0026760|arm
null|Upper Extremity|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C1522541;C5400986;C4761640;C1824218;C3715044;C3495676;C0026760|armnull|Trunk of elephant|Anatomy|false|false||Trunk
null|Trunk structure|Anatomy|false|false||Trunk
null|dendritic shaft|Anatomy|false|false||Trunknull|Pelvis>Groin|Anatomy|false|false||Groin
null|Inguinal region|Anatomy|false|false||Groin
null|Inguinal part of abdomen|Anatomy|false|false||Groinnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|Kneenull|Knee region structure|Anatomy|false|false|C0562271|Knee
null|Knee|Anatomy|false|false|C0562271|Knee
null|Lower extremity>Knee|Anatomy|false|false|C0562271|Knee
null|Knee joint|Anatomy|false|false|C0562271|Kneenull|Multiple Epiphyseal Dysplasia|Disorder|false|false|C0230445;C1305418|Mednull|Master of Education|Finding|false|false|C0230445;C1305418|Med
null|COMP wt Allele|Finding|false|false|C0230445;C1305418|Med
null|COL9A3 gene|Finding|false|false|C0230445;C1305418|Med
null|SCN8A wt Allele|Finding|false|false|C0230445;C1305418|Med
null|COL9A2 gene|Finding|false|false|C0230445;C1305418|Med
null|COMP gene|Finding|false|false|C0230445;C1305418|Med
null|SCN8A gene|Finding|false|false|C0230445;C1305418|Mednull|Structure of calf of leg|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C0026760|Calf
null|null|Anatomy|false|false|C4321267;C1419866;C1549978;C5781216;C1456376;C1413596;C1413597;C0026760|Calfnull|Cattle calf (organism)|Entity|false|false||Calfnull|Clava structure (body structure)|Anatomy|false|false||Grtnull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Thigh|Anatomy|false|false||Thigh
null|Thigh structure|Anatomy|false|false||Thighnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|CDAN1 wt Allele|Finding|false|false||Dlt
null|CDAN1 gene|Finding|false|false||Dltnull|imidazole mustard|Drug|false|false|C3495985;C0175372|Bic
null|imidazole mustard|Drug|false|false|C3495985;C0175372|Bicnull|MIR155HG gene|Finding|false|false|C3495985;C0175372|Bic
null|MIR155 gene|Finding|false|false|C3495985;C0175372|Bicnull|BIC Regimen|Procedure|false|false|C3495985;C0175372|Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|imidazole mustard|Drug|false|false|C3495985;C0175372|Bic
null|imidazole mustard|Drug|false|false|C3495985;C0175372|Bicnull|MIR155HG gene|Finding|false|false|C3495985;C0175372|Bic
null|MIR155 gene|Finding|false|false|C3495985;C0175372|Bicnull|BIC Regimen|Procedure|false|false|C3495985;C0175372|Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false|C0063382;C1537811;C2681931;C5202575|Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Fenamole|Drug|false|false||Pat
null|Fenamole|Drug|false|false||Patnull|Paroxysmal atrial tachycardia|Disorder|false|false||Patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||Pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||Pat
null|protein acetyltransferase activity|Finding|false|false||Patnull|Thermoacoustic Computed Tomography|Procedure|false|false||Patnull|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Achnull|Achondroplasia|Disorder|false|false||Achnull|FGFR3 wt Allele|Finding|false|false||Ach
null|FGFR3 gene|Finding|false|false||Ach
null|Ache|Finding|false|false||Achnull|Acoli Language|Entity|false|false||Achnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Babinski Reflex|Finding|false|false||Babinskinull|Clonus|Finding|false|false||Clonusnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|null|Attribute|false|false|C2752558;C0037949;C0581269;C0817096|MR THORACIC SPINEnull|Thoracic spine structure|Anatomy|false|false|C0009924;C0150920;C0882557;C5779551|THORACIC SPINEnull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false|C0817096;C2752558;C0037949;C0581269|THORACICnull|Chest|Anatomy|false|false|C0150920;C5779551;C0882557|THORACICnull|Spine Problem|Finding|false|false|C0817096;C2752558;C0037949;C0581269|SPINEnull|Neuron spine|Anatomy|false|false|C0150920;C0882557;C5779551|SPINE
null|Vertebral column|Anatomy|false|false|C0150920;C0882557;C5779551|SPINEnull|Contrast Media|Drug|false|false|C0581269|CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Spine Problem|Finding|false|false|C2752558;C0037949|SPINEnull|Neuron spine|Anatomy|false|false|C0150920|SPINE
null|Vertebral column|Anatomy|false|false|C0150920|SPINEnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Central cord canal structure|Anatomy|false|false|C1879652;C3854333|central canalnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false|C0459414|centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false|C0459414|narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Level 5|Modifier|false|false||5 levelnull|Abnormal degeneration|Finding|false|false||degenerative changesnull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|LARGE1 wt Allele|Finding|false|false||Large
null|LARGE1 gene|Finding|false|false||Largenull|Large|LabModifier|false|false||Largenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Paramedian approach|Modifier|false|false||paramediannull|Upper|Modifier|false|false||superiornull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C1621443;C1556138|disc
null|Discontinued|Finding|false|false|C1621443;C1556138|discnull|Disc - Body Part|Anatomy|false|false|C0993608;C1696131;C1444662;C0443213|disc
null|death-inducing signaling complex location|Anatomy|false|false|C0993608;C1696131;C1444662;C0443213|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Extrusion|Finding|false|false|C1621443;C1556138|extrusionnull|Level 5|Modifier|false|false||5 levelnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lateral|Modifier|false|false||lateralnull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Nerve|Anatomy|false|false|C5203119;C1547231;C0205082;C1547227;C1561581;C3854333|nervesnull|Severe - Severity of Illness Code|Finding|false|false|C0027740|severe
null|Intensity and Distress 5|Finding|false|false|C0027740|severe
null|Severe - Triage Code|Finding|false|false|C0027740|severe
null|Severe (severity modifier)|Finding|false|false|C0027740|severe
null|Allergy Severity - Severe|Finding|false|false|C0027740|severenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false|C0027740|narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Advanced phase|Modifier|false|false||Advancednull|Abnormal degeneration|Finding|false|false|C0024090;C0024091;C3887615|degenerative changesnull|biologic degeneration|Finding|false|false|C0024091;C3887615;C2752558;C0037949|degenerative
null|Abnormal degeneration|Finding|false|false|C0024091;C3887615;C2752558;C0037949|degenerativenull|Changing|Finding|false|false|C0024090;C2752558;C0037949;C0024091;C3887615|changesnull|Changed status|LabModifier|false|false||changesnull|Lumbar spine structure|Anatomy|false|false|C0150920;C0011164;C0011164;C1880269;C0392747|lumbar spine
null|Bone structure of lumbar vertebra|Anatomy|false|false|C0150920;C0011164;C0011164;C1880269;C0392747|lumbar spinenull|Lumbar Region|Anatomy|false|false|C0011164;C0392747;C0150920|lumbarnull|Spine Problem|Finding|false|false|C0024091;C3887615;C2752558;C0037949;C0024090|spinenull|Neuron spine|Anatomy|false|false|C0150920;C0392747;C0011164;C1880269|spine
null|Vertebral column|Anatomy|false|false|C0150920;C0392747;C0011164;C1880269|spinenull|Moderate - Severity of Illness Code|Finding|false|false|C0459414|Moderate
null|Moderate|Finding|false|false|C0459414|Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Central cord canal structure|Anatomy|false|false|C3854333;C1879652;C5201148;C1547226|central canalnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false|C0459414;C0086881;C1550227|centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false|C3854333;C1879652|canal
null|Pulp Canals|Anatomy|false|false|C3854333;C1879652|canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false|C0459414;C0086881;C1550227|narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Moderate to severe|Modifier|false|false||moderate to severenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Levels (qualifier value)|Modifier|false|false||levelsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false|C0024091;C3887615|narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Lumbar spine structure|Anatomy|false|false|C0150920;C3854333|lumbar spine
null|Bone structure of lumbar vertebra|Anatomy|false|false|C0150920;C3854333|lumbar spinenull|Lumbar Region|Anatomy|false|false|C0150920|lumbarnull|Spine Problem|Finding|false|false|C2752558;C0037949;C0024091;C3887615;C0024090|spinenull|Neuron spine|Anatomy|false|false|C0150920|spine
null|Vertebral column|Anatomy|false|false|C0150920|spinenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Abnormal degeneration|Finding|false|false|C0581269;C0817096|Degenerative changesnull|biologic degeneration|Finding|false|false|C2752558;C0037949;C0817096;C0581269|Degenerative
null|Abnormal degeneration|Finding|false|false|C2752558;C0037949;C0817096;C0581269|Degenerativenull|Changing|Finding|false|false|C0817096;C0581269|changesnull|Changed status|LabModifier|false|false||changesnull|Thoracic spine structure|Anatomy|false|false|C0011164;C1547225;C0392747;C0150920;C0011164;C1880269;C5201148;C1547226;C5779551|thoracic spinenull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false|C0817096;C0581269|thoracicnull|Chest|Anatomy|false|false|C0392747;C0011164;C0011164;C1880269;C0150920;C5779551|thoracicnull|Spine Problem|Finding|false|false|C2752558;C0037949;C0817096;C0581269|spinenull|Neuron spine|Anatomy|false|false|C0150920;C1547225;C0011164;C1880269|spine
null|Vertebral column|Anatomy|false|false|C0150920;C1547225;C0011164;C1880269|spinenull|Mild to moderate|Modifier|false|false||mild-to-moderatenull|Mild Severity of Illness Code|Finding|false|false|C0581269;C2752558;C0037949|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Moderate - Severity of Illness Code|Finding|false|false|C0581269|moderate
null|Moderate|Finding|false|false|C0581269|moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|null|Attribute|false|false|C0449202;C0000726|CT ABDnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C0153663;C3811055;C1644645;C0812455|ABD
null|Abdomen|Anatomy|false|false|C0153663;C3811055;C1644645;C0812455|ABDnull|Malignant neoplasm of pelvis|Disorder|false|false|C0449202;C0000726;C4266535;C0030797;C0559769|PELVISnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769;C0449202;C0000726|PELVISnull|Pelvis+|Anatomy|false|false|C0153663;C0812455|PELVIS
null|Pelvic cavity structure|Anatomy|false|false|C0153663;C0812455|PELVIS
null|Pelvis|Anatomy|false|false|C0153663;C0812455|PELVISnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Admission Level of Care Code - Acute|Finding|true|false|C0230168;C0000726|acute
null|Acute - Triage Code|Finding|true|false|C0230168;C0000726|acutenull|acute|Time|false|false||acutenull|findings aspects|Finding|false|false|C0230168;C0000726|findingsnull|null|Attribute|false|false||findingsnull|Malignant neoplasm of abdomen|Disorder|true|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|true|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0941288;C0153662;C0812455;C2607943;C0153663;C1547295;C1547229|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662;C0812455;C2607943;C0153663;C1547295;C1547229|abdomennull|Malignant neoplasm of pelvis|Disorder|true|false|C4266535;C0030797;C0559769;C0230168;C0000726|pelvisnull|Pelvis problem|Finding|true|false|C4266535;C0030797;C0559769;C0230168;C0000726|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663|pelvisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Obstructed|Finding|true|false||obstructivenull|Nephrolithiasis|Disorder|false|false|C0022646|renal stonenull|Renal stone (substance)|Finding|false|false|C0022646|renal stone
null|Kidney Calculi|Finding|false|false|C0022646|renal stonenull|Urologic Diseases|Disorder|false|false|C0022646|renalnull|Kidney|Anatomy|false|false|C0392525;C0022650;C1458136;C0006736;C0042075|renalnull|Calculi|Finding|false|false|C0022646|stonenull|Pyelonephritis|Disorder|false|false||pyelonephritisnull|Diverticulosis of sigmoid colon|Disorder|false|false|C0227391|Sigmoid diverticulosisnull|Sigmoid colon|Anatomy|false|false|C0012818;C1510475|Sigmoidnull|Diverticulosis|Disorder|false|false|C0227391|diverticulosisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Diverticulitis|Disorder|false|false||diverticulitisnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||Labsnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Low Back Pain|Finding|false|false||Low Back painnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Back Pain|Finding|false|false|C1140621;C0023216|Back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in lower limb|Finding|false|false|C1140621;C0023216|Leg Painnull|Leg|Anatomy|false|false|C0023222;C1549543;C0030193;C0004604|Leg
null|Lower Extremity|Anatomy|false|false|C0023222;C1549543;C0030193;C0004604|Legnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216|Pain
null|Pain|Finding|false|false|C1140621;C0023216|Painnull|null|Attribute|false|false||Painnull|Radiculopathy|Disorder|false|false||Radiculopathynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|right-sided low back pain|Finding|false|false|C0230102;C2939142;C1548802|right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false|C1548802;C0230102;C2939142|lower back painnull|Lower back (surface region)|Anatomy|false|false|C2219286;C0024031|lower back
null|Lower back structure|Anatomy|false|false|C2219286;C0024031|lower backnull|Body Site Modifier - Lower|Anatomy|false|false|C1549543;C0030193;C2003888;C0004604;C0024031;C2219286|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false|C1548802|back painnull|Administration Method - Pain|Finding|false|false|C1548802|pain
null|Pain|Finding|false|false|C1548802|painnull|null|Attribute|false|false||painnull|Prominent|Modifier|false|false||prominentnull|Protein Component|Drug|false|false||component
null|Protein Component|Drug|false|false||componentnull|Specimen Child Role - Component|Finding|false|false||component
null|Component (part)|Finding|false|false||component
null|Component, LOINC Axis 1|Finding|false|false||componentnull|Component object|Device|false|false||componentnull|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT A
null|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT Anull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Visceral|Modifier|false|false||visceralnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Nephrolithiasis|Disorder|false|false||nephrolithiasisnull|CYREN gene|Finding|false|false|C3887615;C2752558;C0037949|MRInull|Magnetic resonance imaging service|Procedure|false|false|C3887615;C2752558;C0037949|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C3887615;C2752558;C0037949|MRInull|Maori Language|Entity|false|false||MRInull|Lumbar spine structure|Anatomy|false|false|C1824234;C0024485;C0587658;C0150920|L spinenull|Spine Problem|Finding|false|false|C3887615;C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C1824234;C0024485;C0587658;C0150920|spine
null|Vertebral column|Anatomy|false|false|C1824234;C0024485;C0587658;C0150920|spinenull|Significant|Finding|false|false|C1621443;C1556138|significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C1621443;C1556138|disc
null|Discontinued|Finding|false|false|C1621443;C1556138|discnull|Disc - Body Part|Anatomy|false|false|C1696131;C1444662;C0993608;C0750502|disc
null|death-inducing signaling complex location|Anatomy|false|false|C1696131;C1444662;C0993608;C0750502|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Swelling|Finding|false|false||bulgenull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Narrow|Modifier|false|false||narrowing ofnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Spinal|Modifier|false|false||spinalnull|canal [body parts]|Anatomy|false|false|C0750502;C0443213|canal
null|Pulp Canals|Anatomy|false|false|C0750502;C0443213|canalnull|Geographic canal|Entity|false|false||canalnull|Extrusion|Finding|false|false|C0086881;C1550227|extrusionnull|Significant|Finding|false|false|C0086881;C1550227;C0228084|significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Fourth lumbar nerve|Anatomy|false|false|C1705917|L4 nervenull|Nerve root structure|Anatomy|false|false|C0750502;C1705917|nerve rootnull|Nerve|Anatomy|false|false|C1705917|nervenull|Tree Root (hierarchy)|Finding|false|false|C0501792;C0027740;C0040452;C1318154;C0228084|rootnull|Tooth root structure|Anatomy|false|false|C1705917|root
null|Root body part|Anatomy|false|false|C1705917|rootnull|Plant Roots|Entity|false|false||rootnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Recent|Time|false|false||recentlynull|Pain in right leg|Finding|false|false|C0230442;C0230415;C1140621;C0023216|right leg painnull|Structure of right lower leg|Anatomy|false|false|C5848135;C1549543;C0030193|right leg
null|Right lower extremity|Anatomy|false|false|C5848135;C1549543;C0030193|right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false|C1140621;C0023216|leg painnull|Leg|Anatomy|false|false|C0023222;C5848135|leg
null|Lower Extremity|Anatomy|false|false|C0023222;C5848135|legnull|Administration Method - Pain|Finding|false|false|C0230442;C0230415|pain
null|Pain|Finding|false|false|C0230442;C0230415|painnull|null|Attribute|false|false||painnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Bursitis|Disorder|false|false||bursitisnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Corticosteroid [EPC]|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroidnull|Current (present time)|Time|false|false||Currentlynull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Compression of umbilical cord|Disorder|true|false|C1550235|cord compression
null|Compression of spinal cord|Disorder|true|false|C1550235|cord compressionnull|Cone-Rod Dystrophy 2|Disorder|false|false|C1550235|cordnull|Cord - Body Parts|Anatomy|false|false|C3489532;C0728907;C0332459;C4551657;C0037926;C0266798;C1257972;C0565514|cordnull|Cord Device|Device|false|false||cordnull|null|Finding|true|false|C1550235|compression
null|Compressed structure|Finding|true|false|C1550235|compressionnull|Compression Therapy|Procedure|true|false|C1550235|compression
null|Data Compression|Procedure|true|false|C1550235|compressionnull|Compression|Phenomenon|true|false|C1550235|compressionnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Ortho-|Finding|false|false|C2752558;C0037949|orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||orthonull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920;C0812371|spine
null|Vertebral column|Anatomy|false|false|C0150920;C0812371|spinenull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|Decompression - action (qualifier value)|Finding|false|false||DECOMPRESSIONnull|Decompression|Procedure|false|false||DECOMPRESSION
null|Decompressive incision|Procedure|false|false||DECOMPRESSIONnull|external decompression|Phenomenon|false|false||DECOMPRESSIONnull|Fused structure|Finding|false|false||FUSIONnull|Fusion procedure|Procedure|false|false||FUSIONnull|Duraplasty|Procedure|false|false||DURAPLASTYnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Dysuria|Finding|false|false||Dysurianull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Recent|Time|false|false||recentlynull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|abdomennull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Specimen Type - Leukocytes|Finding|false|false|C0023516|leukocytes
null|null|Finding|false|false|C0023516|leukocytesnull|Leukocytes|Anatomy|false|false|C1550647;C1547962|leukocytesnull|Leukocytes|Anatomy|false|false||WBCnull|Urine culture|Procedure|false|false||urine culturenull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Bacterial|Modifier|false|false||bacterialnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Contamination|Finding|false|false||contaminationnull|adulteration|Phenomenon|false|false||contaminationnull|Specimen Reject Reason - Contamination|Modifier|false|false||contaminationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Abdominal Pain|Finding|false|false|C0000726|Abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Constipation|Finding|false|false||constipationnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|opioid use|Disorder|false|false||opioid usenull|Opioids|Drug|false|false||opioid
null|Opioids|Drug|false|false||opioid
null|Opioids|Drug|false|false||opioidnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Report (document)|Finding|false|false||Reportsnull|Reporting|Procedure|false|false||Reportsnull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Bactrim DS|Drug|false|false||bactrim DS
null|Bactrim DS|Drug|false|false||bactrim DSnull|Bactrim|Drug|false|false||bactrim
null|Bactrim|Drug|false|false||bactrimnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Medical History|Finding|false|false|C5239664|History ofnull|History of present illness (finding)|Finding|false|false|C5239664|History
null|History of previous events|Finding|false|false|C5239664|History
null|Historical aspects qualifier|Finding|false|false|C5239664|History
null|Medical History|Finding|false|false|C5239664|History
null|Concept History|Finding|false|false|C5239664|Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0262926;C0262926;C1705255;C0019665;C0262512;C2004062;C0149871;C0151950;C2926618|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Antiphospholipid Syndrome|Disorder|false|false|C1167408;C3665580|Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false|C1167408;C3665580|Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibodynull|Antibody (immunoassay)|Procedure|false|false|C1167408;C3665580|antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false|C4551530;C4019436;C0003241;C0021027;C0085278;C0162595|antibody
null|immunoglobulin complex location|Anatomy|false|false|C4551530;C4019436;C0003241;C0021027;C0085278;C0162595|antibodynull|Syndrome|Disorder|false|false||syndromenull|Lupus anticoagulant positive|Lab|false|false||Lupus anticoagulant positivenull|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulant
null|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulantnull|Lupus anticoagulant disorder|Disorder|false|false||Lupus anticoagulantnull|null|Finding|false|false||Lupus anticoagulantnull|Lupus anticoagulant assay|Procedure|false|false||Lupus anticoagulantnull|Chronic discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus|Disorder|false|false||Lupus
null|Lupus Vulgaris|Disorder|false|false||Lupus
null|Discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus, Systemic|Disorder|false|false||Lupusnull|Anti-coagulant [EPC]|Drug|false|false||anticoagulant
null|Anticoagulants|Drug|false|false||anticoagulantnull|Bilateral|Modifier|false|false||bilateralnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|day|Time|false|false||daysnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Charts (publication)|Finding|false|false||chartnull|chart [medical device]|Device|false|false||chartnull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|null|Attribute|false|false|C0449202;C0000726|CT abdnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|abdnull|ABD (body structure)|Anatomy|false|false|C0153663;C1644645;C3811055|abd
null|Abdomen|Anatomy|false|false|C0153663;C1644645;C3811055|abdnull|Malignant neoplasm of pelvis|Disorder|false|false|C0449202;C0000726;C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0812455;C0153663|pelvis
null|Pelvis|Anatomy|false|false|C0812455;C0153663|pelvisnull|Aortic Aneurysm, Abdominal|Disorder|false|false|C0003483;C0000726|abdominal aortic aneurysmnull|null|Attribute|false|false|C0003483;C0000726|abdominal aortic aneurysmnull|Abdomen|Anatomy|false|false|C0002940;C2926614;C0003486;C0340629;C0162871|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|null|Disorder|false|false|C0003483;C0000726|aortic aneurysm
null|Aortic Aneurysm|Disorder|false|false|C0003483;C0000726|aortic aneurysmnull|Aorta|Anatomy|false|false|C0162871;C2926614;C0003486;C0340629;C0002940|aorticnull|Aneurysm|Finding|false|false|C0000726;C0003483|aneurysmnull|Vitamin D Deficiency|Disorder|false|false||Vitamin D deficiencynull|Decreased circulating vitamin D concentration|Finding|false|false||Vitamin D deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Daily|Time|false|false||dailynull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPAPnull|Continuous Positive Airway Pressure|Procedure|false|false||CPAPnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||Medsnull|Medications|Finding|false|false||Medsnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|Daily|Time|false|false||dailynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|Opioids|Drug|false|false||opioids
null|Opioids|Drug|false|false||opioids
null|Opioids|Drug|false|false||opioids
null|Analgesics, Opioid|Drug|false|false||opioids
null|Analgesics, Opioid|Drug|false|false||opioidsnull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Daily|Time|false|false||dailynull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Rare|Modifier|false|false||rarelynull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Ortho-|Finding|false|false||Orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||Orthonull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920|spine
null|Vertebral column|Anatomy|false|false|C0150920|spinenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|Cerebral Aneurysm|Disorder|false|false|C0228174;C0006104|cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0162871;C0917996;C0002940|cerebral
null|Brain|Anatomy|false|false|C0162871;C0917996;C0002940|cerebralnull|Aortic Aneurysm, Abdominal|Disorder|false|false|C0000726;C0228174;C0006104;C0003483|aneurysm, abdominal aorticnull|Aneurysm|Finding|false|false|C0228174;C0006104|aneurysmnull|Abdomen|Anatomy|false|false|C0162871|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Aorta|Anatomy|false|false|C0162871|aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Pallister W syndrome|Disorder|false|false||syndrome wnull|Syndrome|Disorder|false|false||syndromenull|Numerous|LabModifier|false|false||multiplenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Event|Event|false|false|C1690938;C3853547;C0687080;C0016504|eventnull|Bilateral|Modifier|false|false||bilateralnull|LARGE1 wt Allele|Finding|false|false|C1690938;C3853547;C0687080;C0016504|large
null|LARGE1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|largenull|Large|LabModifier|false|false||largenull|Personal Experience Scales|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEs
null|PES1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false|C1418467;C0687136;C0441471;C5890938;C1416798;C0851145|PEs
null|Hindfoot of quadruped|Anatomy|false|false|C1418467;C0687136;C0441471;C5890938;C1416798;C0851145|PEs
null|Paw|Anatomy|false|false|C1418467;C0687136;C0441471;C5890938;C1416798;C0851145|PEs
null|Foot|Anatomy|false|false|C1418467;C0687136;C0441471;C5890938;C1416798;C0851145|PEsnull|Iranian Persian language|Entity|false|false||PEsnull|on warfarin|Procedure|false|false|C1690938;C3853547;C0687080;C0016504|on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|BRCA1 gene mutation|Disorder|false|false||BRCA1 mutationnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||mutationnull|Mutation|Finding|false|false||mutationnull|Malignant neoplasm of breast|Disorder|false|false|C0006141|breast cancer
null|Breast Carcinoma|Disorder|false|false|C0006141|breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false|C0006141|breastnull|Breast problem|Finding|false|false|C0006141|breastnull|Procedures on breast|Procedure|false|false|C0006141|breastnull|Breast|Anatomy|false|false|C0567499;C0496956;C0006826;C0191838;C0006142;C0678222|breastnull|Malignant Neoplasms|Disorder|false|false|C0006141|cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Transaction counts and value totals - month|Finding|false|false|C1548802;C0230102;C2939142|month
null|Precision - month|Finding|false|false|C1548802;C0230102;C2939142|monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|right-sided low back pain|Finding|false|false|C0230102;C2939142;C1548802|right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false|C0230102;C2939142;C1548802|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false|C1548802;C0230102;C2939142|lower back painnull|Lower back (surface region)|Anatomy|false|false|C2219286;C0004604;C2598155;C1552823;C0024031;C1561541;C1561542;C1549543;C0030193|lower back
null|Lower back structure|Anatomy|false|false|C2219286;C0004604;C2598155;C1552823;C0024031;C1561541;C1561542;C1549543;C0030193|lower backnull|Body Site Modifier - Lower|Anatomy|false|false|C2598155;C0004604;C1561541;C1561542;C0024031;C2219286;C1552823;C2003888;C1549543;C0030193|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false|C0230102;C2939142;C1548802|back painnull|Administration Method - Pain|Finding|false|false|C0230102;C2939142;C1548802|pain
null|Pain|Finding|false|false|C0230102;C2939142;C1548802|painnull|null|Attribute|false|false|C1548802;C0230102;C2939142|painnull|Radicular pain|Finding|false|false||radicular painnull|Dermatomal|Modifier|false|false||radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in right leg|Finding|false|false|C1140621;C0023216;C0230442;C0230415|right leg painnull|Structure of right lower leg|Anatomy|false|false|C0023222;C0750502;C1696131;C1444662;C1552823;C1549543;C0030193;C2598155;C5848135|right leg
null|Right lower extremity|Anatomy|false|false|C0023222;C0750502;C1696131;C1444662;C1552823;C1549543;C0030193;C2598155;C5848135|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C0230442;C0230415;C1140621;C0023216|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false|C0230442;C0230415;C1140621;C0023216;C1621443;C1556138|leg painnull|Leg|Anatomy|false|false|C5848135;C2598155;C1549543;C0030193;C0023222;C1552823|leg
null|Lower Extremity|Anatomy|false|false|C5848135;C2598155;C1549543;C0030193;C0023222;C1552823|legnull|Administration Method - Pain|Finding|false|false|C1140621;C0023216;C1621443;C1556138;C0230442;C0230415|pain
null|Pain|Finding|false|false|C1140621;C0023216;C1621443;C1556138;C0230442;C0230415|painnull|null|Attribute|false|false|C1140621;C0023216;C0230442;C0230415|painnull|Significant|Finding|false|false|C0230442;C0230415|significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Intervertebral Disk Displacement|Disorder|false|false|C1621443;C1556138|disc herniationsnull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C1621443;C1556138;C0230442;C0230415|disc
null|Discontinued|Finding|false|false|C1621443;C1556138;C0230442;C0230415|discnull|Disc - Body Part|Anatomy|false|false|C1696131;C1444662;C1549543;C0030193;C0021818;C0023222;C0993608|disc
null|death-inducing signaling complex location|Anatomy|false|false|C1696131;C1444662;C1549543;C0030193;C0021818;C0023222;C0993608|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Hernia|Disorder|false|false||herniationsnull|Diskectomy|Procedure|false|false||discectomynull|Fused structure|Finding|false|false||fusionnull|Fusion procedure|Procedure|false|false||fusionnull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Course|Time|false|false||coursenull|Relationship modifier - Patient|Finding|false|false|C2752558;C0037949|Patient
null|Specimen Type - Patient|Finding|false|false|C2752558;C0037949|Patient
null|Mail Claim Party - Patient|Finding|false|false|C2752558;C0037949|Patient
null|Report source - Patient|Finding|false|false|C2752558;C0037949|Patient
null|null|Finding|false|false|C2752558;C0037949|Patient
null|Disabled Person Code - Patient|Finding|false|false|C2752558;C0037949|Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Procedure on spinal cord (procedure)|Procedure|false|false|C2752558;C0037949|Spine Surgery
null|Operation on spinal cord (procedure)|Procedure|false|false|C2752558;C0037949|Spine Surgerynull|Spine Problem|Finding|false|false|C2752558;C0037949|Spinenull|Neuron spine|Anatomy|false|false|C0543467;C3245478;C0150920;C0038895;C1457907;C1547138;C0920347;C2608059;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485|Spine
null|Vertebral column|Anatomy|false|false|C0543467;C3245478;C0150920;C0038895;C1457907;C1547138;C0920347;C2608059;C1578483;C1550655;C1578481;C1578486;C1578484;C1578485|Spinenull|Level of Care - Surgery|Finding|false|false|C2752558;C0037949|Surgery
null|Surgical procedure finding|Finding|false|false|C2752558;C0037949|Surgery
null|Surgical aspects|Finding|false|false|C2752558;C0037949|Surgerynull|Operative Surgical Procedures|Procedure|false|false|C2752558;C0037949|Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|ActInformationPrivacyReason - service|Finding|false|false|C2752558;C0037949|Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Operating Room|Device|false|false||Operating Roomnull|Operating Room|Entity|false|false||Operating Roomnull|Patient location type - Operating Room|Modifier|false|false||Operating Roomnull|Operating|Finding|false|false||Operatingnull|Room - Patient location type|Modifier|false|false||Room
null|Room|Modifier|false|false||Roomnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|null|Attribute|false|false||operative notenull|Operative|Time|false|false||operativenull|Further|Modifier|false|false||furthernull|Details|Modifier|false|false||detailsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Complication (attribute)|Finding|false|false||complication
null|Complication|Finding|false|false||complicationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Postoperative deep vein thrombosis|Disorder|false|false|C5239664|Postoperative DVTnull|Postoperative Period|Time|false|false||Postoperativenull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2926618;C0589110;C3469826;C3470073|DVTnull|null|Attribute|false|false|C5239664|DVTnull|SLC35G1 gene|Finding|false|false|C5239664|post
null|DESI1 gene|Finding|false|false|C5239664|postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Bed rest|Procedure|false|false||bedrestnull|Dural tear|Disorder|false|false||dural tearnull|Laceration|Disorder|false|false||tear
null|Rupture|Disorder|false|false||tearnull|Tears (substance)|Finding|false|false||tearnull|Tear Shape|Modifier|false|false||tearnull|Precaution|Finding|false|false||precautionsnull|Hour|Time|false|false||hoursnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|Intravenous Route of Administration|Finding|false|false||Intravenousnull|Intravenous|Modifier|false|false||Intravenousnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Postoperative Period|Time|false|false||postopnull|Type of Agreement - Standard|Finding|false|false||standard
null|Standard (document)|Finding|false|false||standardnull|Standard base excess calculation technique|Procedure|false|false||standardnull|Standard (qualifier)|Modifier|false|false||standardnull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Pain, Postoperative|Finding|false|false||postop painnull|Postoperative Period|Time|false|false||postopnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical therapynull|Physical therapy|Procedure|false|false||Physical therapynull|Physical therapy (field)|Title|false|false||Physical therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Diagnostic Service Section ID - Occupational Therapy|Finding|false|false||Occupational therapynull|Occupational therapy (procedure)|Procedure|false|false||Occupational therapynull|Occupational|Finding|false|false||Occupationalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|physical therapy mobilization (treatment)|Procedure|false|false||mobilization
null|Mobilization (procedure)|Procedure|false|false||mobilizationnull|Ambulate|Finding|false|false||ambulatenull|VISCERAL LEIOMYOPATHY, AFRICAN DEGENERATIVE|Disorder|false|false||ADLnull|Activity of daily living (function)|Finding|false|false||ADL
null|SGCA gene|Finding|false|false||ADL
null|SGCA wt Allele|Finding|false|false||ADLnull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Course|Time|false|false||coursenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||acute blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||acute blood loss anemianull|Acute hemorrhage|Finding|false|false||acute blood lossnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||blood loss anemia
null|Anemia due to blood loss|Disorder|false|false||blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||blood loss anemianull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Constipation|Finding|false|false||constipationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hypokalemia|Finding|false|false||hypokalemianull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||Acute blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||Acute blood loss anemianull|Acute hemorrhage|Finding|false|false||Acute blood lossnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||blood loss anemia
null|Anemia due to blood loss|Disorder|false|false||blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||blood loss anemianull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|Immediate Release Dosage Form|Drug|false|false||Immediate releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Valium|Drug|false|false||Valium
null|Valium|Drug|false|false||Valiumnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Drug|false|false|C0226896|Oral Potassiumnull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C4553027;C0357141;C1527415;C4521986;C0202194;C1272919|Oralnull|Oral|Modifier|false|false||Oralnull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false|C0226896|Potassiumnull|Potassium measurement|Procedure|false|false|C0226896|Potassiumnull|Hypokalemia|Finding|false|false||hypokalemianull|Laboratory test finding|Lab|false|false||labsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hospital course|Finding|false|false||Hospital coursenull|null|Attribute|false|false||Hospital coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||coursenull|null|Modifier|false|false||unremarkablenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Feeling comfortable|Finding|false|false||comfortablenull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C0221776;C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false|C0524470|Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false|C0524470|PTCH
null|PTCH1 wt Allele|Finding|false|false|C0524470|PTCH
null|PTCH1 gene|Finding|false|false|C0524470|PTCH
null|PTCH1 protein, human|Finding|false|false|C0524470|PTCHnull|Every morning|Time|false|false||QAMnull|Right hip region structure|Anatomy|false|false|C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C0332461;C1552823;C4308013;C1826732;C0694887;C1705339|right hipnull|Table Cell Horizontal Align - right|Finding|false|false|C0524470|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Hip structure|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Bone structure of ischium|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hipnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false|C1140621;C0023216|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|Leg swellingnull|Leg|Anatomy|false|false|C1422467;C0581394;C0013604;C0038999|Leg
null|Lower Extremity|Anatomy|false|false|C1422467;C0581394;C0013604;C0038999|Legnull|Swelling|Finding|false|false|C1140621;C0023216|swelling
null|Edema|Finding|false|false|C1140621;C0023216|swellingnull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|diazepam|Drug|false|false||Diazepam
null|diazepam|Drug|false|false||Diazepamnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Spasm|Finding|false|false||spasm
null|KANTR gene|Finding|false|false||spasmnull|Somnolence|Disorder|false|false||drowsinessnull|Drowsiness|Finding|false|false||drowsinessnull|diazepam|Drug|false|false||diazepam
null|diazepam|Drug|false|false||diazepamnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid Syndromenull|Syndrome|Disorder|false|false||Syndromenull|Biomaterial Treatment|Finding|false|false||Treatment
null|Treating|Finding|false|false||Treatment
null|therapeutic aspects|Finding|false|false||Treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||Treatment
null|Administration (procedure)|Procedure|false|false||Treatment
null|Therapeutic procedure|Procedure|false|false||Treatmentnull|Fixation of dental bridge|Procedure|false|false||Bridgenull|Type of bridge device|Device|false|false||Bridgenull|morphine sulfate|Drug|false|false||Morphine Sulfate
null|morphine sulfate|Drug|false|false||Morphine Sulfatenull|morphine|Drug|false|false||Morphine
null|morphine|Drug|false|false||Morphinenull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Intrinsic drive|Finding|false|false||drivenull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false|C1140621;C0023216|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|Leg swellingnull|Leg|Anatomy|false|false|C0581394;C1422467;C0013604;C0038999|Leg
null|Lower Extremity|Anatomy|false|false|C0581394;C1422467;C0013604;C0038999|Legnull|Swelling|Finding|false|false|C1140621;C0023216|swelling
null|Edema|Finding|false|false|C1140621;C0023216|swellingnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false|C0524470|Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false|C0524470|PTCH
null|PTCH1 wt Allele|Finding|false|false|C0524470|PTCH
null|PTCH1 gene|Finding|false|false|C0524470|PTCH
null|PTCH1 protein, human|Finding|false|false|C0524470|PTCHnull|Every morning|Time|false|false||QAMnull|Right hip region structure|Anatomy|false|false|C0332461;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890;C1552823;C4308013;C1826732;C0694887;C1705339|right hipnull|Table Cell Horizontal Align - right|Finding|false|false|C0524470|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0524470;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Hip structure|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hip
null|Bone structure of ischium|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1292890|hipnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Spinal stenosis of lumbar region|Disorder|false|false|C0024090|Lumbar spinal stenosisnull|Lumbar Region|Anatomy|false|false|C0037944;C1861329;C0158288;C1261287|Lumbarnull|Spinal canal stenosis|Disorder|false|false|C0024090|spinal stenosis
null|Spinal Stenosis|Disorder|false|false|C0024090|spinal stenosisnull|Spinal|Modifier|false|false||spinalnull|Stenosis|Finding|false|false|C0024090|stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Spondylolisthesis, L4-L5|Finding|false|false||Spondylolisthesis, L4-L5null|Congenital spondylolisthesis|Disorder|false|false||Spondylolisthesis
null|Spondylolisthesis|Disorder|false|false||Spondylolisthesis
null|Acquired spondylolisthesis|Disorder|false|false||Spondylolisthesisnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Constipation|Finding|false|false||Constipationnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis|Procedure|false|false||Diagnosesnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false|C5239664|History
null|History of previous events|Finding|false|false|C5239664|History
null|Historical aspects qualifier|Finding|false|false|C5239664|History
null|Medical History|Finding|false|false|C5239664|History
null|Concept History|Finding|false|false|C5239664|Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0262926;C1705255;C0019665;C0262512;C2004062;C0149871;C0151950;C2926618|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Antiphospholipid Syndrome|Disorder|false|false|C1167408;C3665580|Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false|C1167408;C3665580|Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibodynull|Antibody (immunoassay)|Procedure|false|false|C1167408;C3665580|antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false|C4019436;C0162595;C0003241;C0021027;C4551530;C0085278;C0039082|antibody
null|immunoglobulin complex location|Anatomy|false|false|C4019436;C0162595;C0003241;C0021027;C4551530;C0085278;C0039082|antibodynull|Syndrome|Disorder|false|false|C1167408;C3665580|syndromenull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPAPnull|Continuous Positive Airway Pressure|Procedure|false|false||CPAPnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false|C0230442;C0230415;C1140621;C0023216|pain
null|Pain|Finding|false|false|C0230442;C0230415;C1140621;C0023216|painnull|null|Attribute|false|false||painnull|Structure of right lower leg|Anatomy|false|false|C1549543;C0030193;C1552823|right leg
null|Right lower extremity|Anatomy|false|false|C1549543;C0030193;C1552823|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C0230442;C0230415;C1140621;C0023216|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false|C1549543;C0030193;C1552823|leg
null|Lower Extremity|Anatomy|false|false|C1549543;C0030193;C1552823|legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Difficult (qualifier value)|Finding|false|false||difficultnull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Intervertebral Disk Displacement|Disorder|false|false|C1621443;C1556138|disc herniationnull|Disk Drug Form|Drug|false|false|C1621443;C1556138|discnull|Disc (List bullets)|Finding|false|false|C1621443;C1556138|disc
null|Discontinued|Finding|false|false|C1621443;C1556138|discnull|Disc - Body Part|Anatomy|false|false|C0019270;C1696131;C1444662;C0993608;C0021818|disc
null|death-inducing signaling complex location|Anatomy|false|false|C0019270;C1696131;C1444662;C0993608;C0021818|discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Hernia|Disorder|false|false|C1621443;C1556138|herniationnull|Lower back (surface region)|Anatomy|false|false|C1549543;C0030193;C2598155;C2003888|lower back
null|Lower back structure|Anatomy|false|false|C1549543;C0030193;C2598155;C2003888|lower backnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0230102;C2939142|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Administration Method - Pain|Finding|false|false|C0230102;C2939142|pain
null|Pain|Finding|false|false|C0230102;C2939142|painnull|null|Attribute|false|false|C0230102;C2939142|painnull|Spine Problem|Finding|false|false|C2752558;C0037949|spinenull|Neuron spine|Anatomy|false|false|C0150920|spine
null|Vertebral column|Anatomy|false|false|C0150920|spinenull|Surgeon|Subject|false|false||surgeonsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Past 30 days|Time|false|false||past monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Decompression of spinal cord|Procedure|false|false||spinal decompression
null|Laminectomy|Procedure|false|false||spinal decompressionnull|Spinal|Modifier|false|false||spinalnull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Urinary tract infection|Disorder|false|false|C0042027;C1185740;C0042027;C1508753|urinary tract infectionnull|Urinary tract|Anatomy|false|false|C0042029;C0009450|urinary tract
null|Urinary system|Anatomy|false|false|C0042029;C0009450|urinary tractnull|Urinary tract|Anatomy|false|false|C0009450;C0042029|urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false|C0009450;C0042029|tractnull|Communicable Diseases|Disorder|false|false|C1185740;C0042027;C0042027;C1508753|infectionnull|Infection|Finding|false|false||infectionnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Lumbar Region|Anatomy|false|false|C0011117;C0021153;C1829459;C1965697|Lumbarnull|Decompression - action (qualifier value)|Finding|false|false|C0024090|Decompressionnull|Decompression|Procedure|false|false|C0024090|Decompression
null|Decompressive incision|Procedure|false|false|C0024090|Decompressionnull|external decompression|Phenomenon|false|false|C0024090|Decompressionnull|Fused structure|Finding|false|false||Fusionnull|Fusion procedure|Procedure|false|false||Fusionnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Lumbar Region|Anatomy|false|false|C0011117;C1965697;C0021153;C1829459|Lumbarnull|Decompression - action (qualifier value)|Finding|false|false|C0024090|Decompressionnull|Decompression|Procedure|false|false|C0024090|Decompression
null|Decompressive incision|Procedure|false|false|C0024090|Decompressionnull|external decompression|Phenomenon|false|false|C0024090|Decompressionnull|Fused structure|Finding|false|false||Fusionnull|Fusion procedure|Procedure|false|false||Fusionnull|Stat (do immediately)|Time|false|false||Immediatelynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Greater|LabModifier|false|false||greaternull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|More|LabModifier|false|false||morenull|Feeling comfortable|Finding|false|false||comfortablenull|Does sit|Finding|true|false||sit
null|Sitting position|Finding|true|false||sit
null|HHAT gene|Finding|true|false||sit
null|SIT1 gene|Finding|true|false||sitnull|Does stand|Finding|true|false||stand
null|standards characteristics|Finding|true|false||standnull|Stand (physical object)|Device|true|false||stand
null|Stand Device|Device|true|false||standnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|45 Minutes|Time|false|false||45 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Encounter due to care involving use of rehabilitation procedures|Finding|false|false||Rehabilitation
null|Rehabilitation aspects|Finding|false|false||Rehabilitationnull|Rehabilitation therapy|Procedure|false|false||Rehabilitationnull|null|Title|false|false||Rehabilitationnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Walking (function)|Finding|false|false||walknull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Much|Finding|false|false||muchnull|Terminology Kind|Finding|false|false||kindnull|null|Modifier|false|false||kindnull|Lifting|Event|false|false||liftingnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|MCL1 wt Allele|Finding|false|false||Eat
null|Eating|Finding|false|false||Eatnull|Diet, Healthy|Finding|false|false||healthy dietnull|Healthy|Modifier|false|false||healthynull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Constipation|Finding|false|false||constipationnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|Application of brace (procedure)|Procedure|false|false||Bracenull|Braces - Orthopedic appliances|Device|false|false||Brace
null|Braces - garment|Device|false|false||Bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Wound care management|Procedure|false|false|C2338258|Wound Care
null|wound care|Procedure|false|false|C2338258|Wound Carenull|Wound Care kit|Device|false|false||Wound Carenull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|In care (finding)|Finding|false|false|C2338258|Care
null|Continuity Assessment Record and Evaluation|Finding|false|false|C2338258|Carenull|care activity|Event|false|false||Carenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0886052;C1272654;C0184898;C0332803;C0580931;C2362566|incisionnull|null|Device|false|false||dry dressingnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Appointments|Event|false|false||appointmentnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Bathing|Procedure|false|false||bathnull|Pool (action)|Finding|false|false||poolnull|Sample pool|Attribute|false|false||poolnull|Pool (environment)|Entity|false|false||poolnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Moist|Modifier|false|false||wetnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Additional|Finding|false|false||Additionalnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|72 Hours|Time|false|false||72 hoursnull|Hour|Time|false|false||hoursnull|refill|Finding|false|false||refillnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Authorization Mode - Fax|Finding|false|false||fax
null|Fax Number|Finding|false|false||faxnull|Facsimile Machine|Device|false|false||fax
null|Telefacsimile|Device|false|false||faxnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Oxycontin|Drug|false|false||oxycontin
null|Oxycontin|Drug|false|false||oxycontinnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|90 days|Time|false|false||90 daysnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Follow-up status|Finding|false|false||Follow upnull|follow-up|Procedure|false|false||Follow upnull|Follow - dosing instruction imperative|Finding|false|false||Follow
null|Follow|Finding|false|false||Follownull|Followed by|Time|false|false||Follownull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Appointments|Event|false|false||appointmentnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Visit|Finding|false|false||visitnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|X-rays, Homeopathic Preparations|Drug|false|false||X-raysnull|Plain x-ray|Procedure|false|false||X-rays
null|Diagnostic radiologic examination|Procedure|false|false||X-raysnull|Roentgen Rays|Phenomenon|false|false||X-raysnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|Full|Modifier|false|false||fullnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Degrees fahrenheit|LabModifier|false|false||Fahrenheitnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|Weight-Bearing state|Subject|false|false||Weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|Bearing Device|Device|false|false||bearingnull|Gait|Finding|false|false||Gaitnull|Balance training|Procedure|false|false||balance trainingnull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|Processing ID - Training|Finding|false|false||trainingnull|Training Programs|Procedure|false|false||training
null|Training|Procedure|false|false||trainingnull|training aspects|Modifier|false|false||trainingnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Decompression Sickness|Disorder|true|false||bendingnull|Bending - Changing basic body position|Finding|true|false||bending
null|Does bend|Finding|true|false||bendingnull|Bent|Modifier|false|false||bendingnull|Musculoskeletal torsion (function)|Finding|true|false||twisting
null|Torsion (malposition)|Finding|true|false||twistingnull|Therapeutic procedure|Procedure|false|false||Treatmentsnull|Frequency|Finding|false|false||Frequency
null|How Often|Finding|false|false||Frequencynull|With frequency|Time|false|false||Frequency
null|Frequencies (time pattern)|Time|false|false||Frequencynull|Kind of quantity - Frequency|LabModifier|false|false||Frequency
null|Statistical Frequency|LabModifier|false|false||Frequency
null|Spatial Frequency|LabModifier|false|false||Frequencynull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|null|Device|false|false||dry dressingnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Bathing|Procedure|false|false||bathnull|Pool (action)|Finding|false|false|C2338258|poolnull|Sample pool|Attribute|false|false|C2338258|poolnull|Pool (environment)|Entity|false|false||poolnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C1509144;C0332803;C0184898;C2349200|incisionnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Moist|Modifier|false|false||wetnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions