 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
M|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
MEDICINE|153,161
<EOL>|161,162
<EOL>|163,164
Corgard|176,183
/|184,185
Vasotec|186,193
<EOL>|193,194
<EOL>|195,196
Attending|196,205
:|205,206
_|207,208
_|208,209
_|209,210
<EOL>|210,211
<EOL>|212,213
leg|230,233
edema|234,239
<EOL>|239,240
<EOL>|241,242
Major|242,247
Surgical|248,256
or|257,259
Invasive|260,268
Procedure|269,278
:|278,279
<EOL>|279,280
None|280,284
<EOL>|284,285
<EOL>|285,286
<EOL>|287,288
HISTORY|316,323
OF|324,326
PRESENTING|327,337
ILLNESS|338,345
:|345,346
<EOL>|348,349
Mr.|350,353
_|354,355
_|355,356
_|356,357
is|358,360
an|361,363
_|364,365
_|365,366
_|366,367
year|368,372
old|373,376
gentleman|377,386
with|387,391
history|392,399
of|400,402
CAD|403,406
<EOL>|407,408
(|408,409
s|409,410
/|410,411
p|411,412
3V|413,415
CABG|416,420
_|421,422
_|422,423
_|423,424
,|424,425
LM|426,428
PCI|429,432
_|433,434
_|434,435
_|435,436
,|436,437
pulmonary|438,447
HTN|448,451
,|451,452
AFib|453,457
on|458,460
<EOL>|461,462
anticoagulation|462,477
,|477,478
_|479,480
_|480,481
_|481,482
(|483,484
EF|484,486
50|487,489
%|489,490
)|490,491
who|492,495
presents|496,504
with|505,509
volume|510,516
overload|517,525
<EOL>|526,527
and|527,530
new|531,534
found|535,540
RV|541,543
dilation|544,552
on|553,555
office|556,562
echocardiogram|563,577
.|577,578
<EOL>|580,581
Patient|582,589
reports|590,597
he|598,600
has|601,604
had|605,608
10|609,611
days|612,616
of|617,619
waking|620,626
up|627,629
feeling|630,637
nervous|638,645
<EOL>|646,647
and|647,650
jittery|651,658
.|658,659
He|660,662
also|663,667
endorses|668,676
weight|677,683
gain|684,688
,|688,689
and|690,693
new|694,697
onset|698,703
lower|704,709
<EOL>|710,711
extremity|711,720
swelling|721,729
.|729,730
He|731,733
has|734,737
not|738,741
had|742,745
chest|746,751
pain|752,756
,|756,757
palpitations|758,770
,|770,771
<EOL>|772,773
orthopnea|773,782
,|782,783
or|784,786
PND|787,790
.|790,791
He|792,794
has|795,798
not|799,802
had|803,806
any|807,810
fevers|811,817
,|817,818
cough|819,824
,|824,825
recent|826,832
<EOL>|833,834
travel|834,840
,|840,841
medication|842,852
non|853,856
compliance|857,867
,|867,868
increased|869,878
salty|879,884
food|885,889
intake|890,896
.|896,897
<EOL>|898,899
He|899,901
also|902,906
has|907,910
not|911,914
had|915,918
dyspnea|919,926
on|927,929
exertion|930,938
and|939,942
rides|943,948
4|949,950
miles|951,956
per|957,960
<EOL>|961,962
day|962,965
on|966,968
a|969,970
stationary|971,981
bike|982,986
and|987,990
does|991,995
6|996,997
minutes|998,1005
of|1006,1008
weight|1009,1015
lifting|1016,1023
.|1023,1024
<EOL>|1026,1027
He|1028,1030
presented|1031,1040
to|1041,1043
Dr.|1044,1047
_|1048,1049
_|1049,1050
_|1050,1051
today|1052,1057
for|1058,1061
evaluation|1062,1072
.|1072,1073
There|1074,1079
<EOL>|1080,1081
he|1081,1083
had|1084,1087
a|1088,1089
TTE|1090,1093
that|1094,1098
showed|1099,1105
new|1106,1109
RV|1110,1112
dilation|1113,1121
and|1122,1125
was|1126,1129
referred|1130,1138
to|1139,1141
the|1142,1145
<EOL>|1146,1147
_|1147,1148
_|1148,1149
_|1149,1150
ED|1151,1153
for|1154,1157
further|1158,1165
evaluation|1166,1176
with|1177,1181
concern|1182,1189
for|1190,1193
pulmonary|1194,1203
<EOL>|1204,1205
embolism|1205,1213
.|1213,1214
<EOL>|1216,1217
<EOL>|1218,1219
In|1220,1222
the|1223,1226
ED|1227,1229
,|1229,1230
initial|1231,1238
vitals|1239,1245
were|1246,1250
:|1250,1251
<EOL>|1253,1254
T98|1255,1258
.|1258,1259
HR|1260,1262
70|1263,1265
,|1265,1266
BP|1267,1269
166|1270,1273
/|1273,1274
65|1274,1276
,|1276,1277
RR|1278,1280
16|1281,1283
,|1283,1284
100|1285,1288
%|1288,1289
RA|1290,1292
.|1292,1293
<EOL>|1295,1296
Exam|1297,1301
in|1302,1304
ED|1305,1307
notable|1308,1315
for|1316,1319
bilateral|1320,1329
pitting|1330,1337
edema|1338,1343
to|1344,1346
knees|1347,1352
.|1352,1353
Labs|1354,1358
<EOL>|1359,1360
notable|1360,1367
for|1368,1371
mild|1372,1376
hyponatremia|1377,1389
,|1389,1390
Cr|1391,1393
1.1|1394,1397
.|1397,1398
ALT|1399,1402
/|1402,1403
AST|1403,1406
mildly|1407,1413
elevated|1414,1422
<EOL>|1423,1424
at|1424,1426
81|1427,1429
/|1429,1430
64|1430,1432
.|1432,1433
WBC|1434,1437
4|1438,1439
,|1439,1440
Hgb|1441,1444
11.3|1445,1449
,|1449,1450
INR|1451,1454
1.3|1455,1458
.|1458,1459
DDimer|1460,1466
<|1467,1468
150|1468,1471
.|1471,1472
UA|1473,1475
<EOL>|1476,1477
unremarkable|1477,1489
.|1489,1490
<EOL>|1492,1493
CXR|1494,1497
with|1498,1502
mild|1503,1507
cardiomegaly|1508,1520
but|1521,1524
no|1525,1527
evidence|1528,1536
of|1537,1539
consolidation|1540,1553
or|1554,1556
<EOL>|1557,1558
pulmonary|1558,1567
edema|1568,1573
.|1573,1574
CTA|1575,1578
was|1579,1582
negative|1583,1591
for|1592,1595
PE|1596,1598
,|1598,1599
showed|1600,1606
severe|1607,1613
<EOL>|1614,1615
emphysema|1615,1624
and|1625,1628
dilated|1629,1636
pulmonary|1637,1646
artery|1647,1653
.|1653,1654
<EOL>|1656,1657
Patient|1658,1665
received|1666,1674
20|1675,1677
mg|1678,1680
IV|1681,1683
Lasix|1684,1689
with|1690,1694
significant|1695,1706
urine|1707,1712
output|1713,1719
<EOL>|1720,1721
per|1721,1724
patient|1725,1732
.|1732,1733
He|1734,1736
was|1737,1740
then|1741,1745
admitted|1746,1754
to|1755,1757
the|1758,1761
heart|1762,1767
failure|1768,1775
service|1776,1783
<EOL>|1784,1785
for|1785,1788
acute|1789,1794
heart|1795,1800
failure|1801,1808
exacerbation|1809,1821
and|1822,1825
further|1826,1833
workup|1834,1840
of|1841,1843
RV|1844,1846
<EOL>|1847,1848
dilation|1848,1856
.|1856,1857
<EOL>|1859,1860
Vitals|1861,1867
on|1868,1870
transfer|1871,1879
:|1879,1880
Afebrile|1881,1889
,|1889,1890
HR|1891,1893
66|1894,1896
,|1896,1897
BP|1898,1900
129|1901,1904
/|1904,1905
54|1905,1907
,|1907,1908
RR|1909,1911
19|1912,1914
,|1914,1915
95|1916,1918
%|1918,1919
RA|1919,1921
.|1921,1922
<EOL>|1924,1925
<EOL>|1926,1927
On|1928,1930
review|1931,1937
of|1938,1940
systems|1941,1948
,|1948,1949
he|1950,1952
denies|1953,1959
any|1960,1963
prior|1964,1969
history|1970,1977
of|1978,1980
stroke|1981,1987
,|1987,1988
<EOL>|1989,1990
TIA|1990,1993
,|1993,1994
deep|1995,1999
venous|2000,2006
thrombosis|2007,2017
,|2017,2018
pulmonary|2019,2028
embolism|2029,2037
,|2037,2038
bleeding|2039,2047
at|2048,2050
the|2051,2054
<EOL>|2055,2056
time|2056,2060
of|2061,2063
surgery|2064,2071
,|2071,2072
myalgias|2073,2081
,|2081,2082
joint|2083,2088
pains|2089,2094
,|2094,2095
cough|2096,2101
,|2101,2102
hemoptysis|2103,2113
,|2113,2114
black|2115,2120
<EOL>|2121,2122
stools|2122,2128
or|2129,2131
red|2132,2135
stools|2136,2142
.|2142,2143
He|2144,2146
denies|2147,2153
recent|2154,2160
fevers|2161,2167
,|2167,2168
chills|2169,2175
or|2176,2178
rigors|2179,2185
.|2185,2186
<EOL>|2187,2188
He|2188,2190
denies|2191,2197
exertional|2198,2208
buttock|2209,2216
or|2217,2219
calf|2220,2224
pain|2225,2229
.|2229,2230
All|2231,2234
of|2235,2237
the|2238,2241
other|2242,2247
<EOL>|2248,2249
review|2249,2255
of|2256,2258
systems|2259,2266
were|2267,2271
negative|2272,2280
.|2280,2281
<EOL>|2283,2284
<EOL>|2285,2286
Cardiac|2287,2294
review|2295,2301
of|2302,2304
systems|2305,2312
is|2313,2315
notable|2316,2323
for|2324,2327
absence|2328,2335
of|2336,2338
chest|2339,2344
pain|2345,2349
,|2349,2350
<EOL>|2351,2352
paroxysmal|2352,2362
nocturnal|2363,2372
dyspnea|2373,2380
,|2380,2381
orthopnea|2382,2391
,|2391,2392
palpitations|2393,2405
,|2405,2406
syncope|2407,2414
<EOL>|2415,2416
or|2416,2418
presyncope|2419,2429
.|2429,2430
<EOL>|2432,2433
<EOL>|2434,2435
<EOL>|2435,2436
<EOL>|2437,2438
<EOL>|2459,2460
BILATERAL|2482,2491
MODERATE|2492,2500
CAROTID|2501,2508
DISEASE|2509,2516
<EOL>|2517,2518
CONGESTIVE|2518,2528
HEART|2529,2534
FAILURE|2535,2542
<EOL>|2543,2544
CORONARY|2544,2552
ARTERY|2553,2559
DISEASE|2560,2567
<EOL>|2568,2569
GASTROESOPHAGEAL|2569,2585
REFLUX|2586,2592
<EOL>|2593,2594
HYPERTENSION|2594,2606
<EOL>|2607,2608
SEVERE|2608,2614
EMPHYSEMA|2615,2624
<EOL>|2625,2626
PULMONARY|2626,2635
HYPERTENSION|2636,2648
<EOL>|2649,2650
RIGHT|2650,2655
BUNDLE|2656,2662
BRANCH|2663,2669
BLOCK|2670,2675
<EOL>|2676,2677
BENIGN|2677,2683
PROSTATIC|2684,2693
HYPERTROPHY|2694,2705
<EOL>|2706,2707
HYPERLIPIDEMIA|2707,2721
<EOL>|2722,2723
PAROXYSMAL|2723,2733
ATRIAL|2734,2740
FIBRILLATION|2741,2753
<EOL>|2754,2755
H|2755,2756
/|2756,2757
O|2757,2758
HISTIOPLASMOSIS|2759,2774
<EOL>|2775,2776
<EOL>|2776,2777
CARDIOVERSION|2800,2813
_|2814,2815
_|2815,2816
_|2816,2817
<EOL>|2818,2819
RIGHT|2819,2824
LOWER|2825,2830
LOBE|2831,2835
LOBECTOMY|2836,2845
_|2846,2847
_|2847,2848
_|2848,2849
<EOL>|2850,2851
CORONARY|2851,2859
BYPASS|2860,2866
SURGERY|2867,2874
_|2875,2876
_|2876,2877
_|2877,2878
<EOL>|2879,2880
<EOL>|2880,2881
<EOL>|2882,2883
:|2897,2898
<EOL>|2898,2899
_|2899,2900
_|2900,2901
_|2901,2902
<EOL>|2902,2903
:|2917,2918
<EOL>|2918,2919
Non-contributory|2919,2935
<EOL>|2935,2936
<EOL>|2937,2938
ADMISSION|2953,2962
<EOL>|2962,2963
Vitals|2963,2969
:|2969,2970
98|2971,2973
159|2974,2977
/|2977,2978
62|2978,2980
16|2981,2983
98|2984,2986
%|2986,2987
on|2988,2990
RA|2991,2993
weight|2994,3000
143|3001,3004
lbs|3005,3008
(|3009,3010
bed|3010,3013
scale|3014,3019
)|3019,3020
<EOL>|3022,3023
General|3024,3031
:|3031,3032
very|3033,3037
pleasant|3038,3046
older|3047,3052
gentleman|3053,3062
lying|3063,3068
in|3069,3071
bed|3072,3075
speaking|3076,3084
in|3085,3087
<EOL>|3088,3089
full|3089,3093
sentences|3094,3103
in|3104,3106
NAD|3107,3110
<EOL>|3112,3113
HEENT|3114,3119
:|3119,3120
PERRL|3121,3126
,|3126,3127
EOMI|3128,3132
,|3132,3133
no|3134,3136
scleral|3137,3144
icterus|3145,3152
,|3152,3153
oropharynx|3154,3164
clear|3165,3170
<EOL>|3172,3173
Neck|3174,3178
:|3178,3179
supple|3180,3186
,|3186,3187
JVP|3188,3191
at|3192,3194
6cm|3195,3198
,|3198,3199
no|3200,3202
adenopathy|3203,3213
<EOL>|3215,3216
CV|3217,3219
:|3219,3220
regular|3221,3228
rate|3229,3233
and|3234,3237
rhythm|3238,3244
,|3244,3245
normal|3246,3252
S1|3253,3255
,|3255,3256
physiologic|3257,3268
split|3269,3274
S2|3275,3277
,|3277,3278
<EOL>|3279,3280
_|3280,3281
_|3281,3282
_|3282,3283
systolic|3284,3292
murmur|3293,3299
at|3300,3302
LLSB|3303,3307
.|3307,3308
No|3309,3311
rubs|3312,3316
or|3317,3319
gallops|3320,3327
.|3327,3328
<EOL>|3330,3331
Lungs|3332,3337
:|3337,3338
CTAB|3339,3343
,|3343,3344
no|3345,3347
crackles|3348,3356
,|3356,3357
wheezes|3358,3365
,|3365,3366
or|3367,3369
rhonchi|3370,3377
<EOL>|3379,3380
Abdomen|3381,3388
:|3388,3389
soft|3390,3394
,|3394,3395
non|3396,3399
distended|3400,3409
,|3409,3410
non|3411,3414
tender|3415,3421
to|3422,3424
deep|3425,3429
palpation|3430,3439
,|3439,3440
+|3441,3442
BS|3442,3444
<EOL>|3445,3446
<EOL>|3447,3448
GU|3449,3451
:|3451,3452
no|3453,3455
CVA|3456,3459
tenderness|3460,3470
,|3470,3471
no|3472,3474
foley|3475,3480
<EOL>|3482,3483
Extr|3484,3488
:|3488,3489
warm|3490,3494
,|3494,3495
well|3496,3500
perfused|3501,3509
,|3509,3510
2|3511,3512
+|3512,3513
pulses|3514,3520
in|3521,3523
radial|3524,3530
and|3531,3534
DP|3535,3537
,|3537,3538
2|3539,3540
+|3540,3541
edema|3542,3547
<EOL>|3548,3549
in|3549,3551
bilateral|3552,3561
lower|3562,3567
extremities|3568,3579
to|3580,3582
knees|3583,3588
<EOL>|3590,3591
Neuro|3592,3597
:|3597,3598
aoxo3|3599,3604
,|3604,3605
CN2|3606,3609
-|3609,3610
12|3610,3612
grossly|3613,3620
intact|3621,3627
,|3627,3628
moving|3629,3635
all|3636,3639
4|3640,3641
extremities|3642,3653
<EOL>|3654,3655
without|3655,3662
deficit|3663,3670
,|3670,3671
stable|3672,3678
gait|3679,3683
<EOL>|3685,3686
Skin|3687,3691
:|3691,3692
warm|3693,3697
,|3697,3698
well|3699,3703
perfused|3704,3712
,|3712,3713
dry|3714,3717
,|3717,3718
no|3719,3721
rashes|3722,3728
or|3729,3731
lesions|3732,3739
<EOL>|3741,3742
<EOL>|3742,3743
DISCHARGE|3743,3752
<EOL>|3752,3753
Vitals|3753,3759
:|3759,3760
98.3|3761,3765
100|3766,3769
-|3769,3770
121|3770,3773
/|3773,3774
49|3774,3776
-|3776,3777
59|3777,3779
54|3780,3782
-|3782,3783
62|3783,3785
18|3786,3788
96RA|3789,3793
<EOL>|3793,3794
Tele|3794,3798
:|3798,3799
no|3800,3802
tele|3803,3807
<EOL>|3807,3808
Last|3808,3812
8|3813,3814
hours|3815,3820
I|3821,3822
/|3822,3823
O|3823,3824
:|3824,3825
_|3826,3827
_|3827,3828
_|3828,3829
<EOL>|3829,3830
Last|3830,3834
24|3835,3837
hours|3838,3843
I|3844,3845
/|3845,3846
O|3846,3847
:|3847,3848
1200|3849,3853
/|3853,3854
3150|3854,3858
<EOL>|3858,3859
Weight|3859,3865
on|3866,3868
admission|3869,3878
:|3878,3879
64.3|3880,3884
<EOL>|3884,3885
Today|3885,3890
's|3890,3892
weight|3893,3899
:|3899,3900
63.1|3901,3905
<EOL>|3905,3906
<EOL>|3906,3907
General|3907,3914
:|3914,3915
elderly|3916,3923
,|3923,3924
NAD|3925,3928
<EOL>|3930,3931
Neck|3931,3935
:|3935,3936
JVP|3937,3940
at|3941,3943
base|3944,3948
of|3949,3951
clavicle|3952,3960
when|3961,3965
90|3966,3968
degrees|3969,3976
<EOL>|3976,3977
Lungs|3977,3982
:|3982,3983
CTAB|3985,3989
no|3990,3992
crackles|3993,4001
<EOL>|4001,4002
CV|4002,4004
:|4004,4005
RRR|4006,4009
,|4009,4010
split|4011,4016
S2|4017,4019
<EOL>|4019,4020
Abdomen|4020,4027
:|4027,4028
slightly|4029,4037
obese|4038,4043
,|4043,4044
soft|4045,4049
,|4049,4050
NTND|4051,4055
,|4055,4056
NABS|4057,4061
<EOL>|4061,4062
Ext|4062,4065
:|4065,4066
no|4067,4069
edema|4070,4075
<EOL>|4075,4076
<EOL>|4077,4078
Pertinent|4078,4087
Results|4088,4095
:|4095,4096
<EOL>|4096,4097
ADMISSION|4097,4106
<EOL>|4106,4107
_|4107,4108
_|4108,4109
_|4109,4110
04|4111,4113
:|4113,4114
02PM|4114,4118
BLOOD|4119,4124
WBC|4125,4128
-|4128,4129
4.0|4129,4132
RBC|4133,4136
-|4136,4137
4|4137,4138
.|4138,4139
32|4139,4141
*|4141,4142
Hgb|4143,4146
-|4146,4147
11|4147,4149
.|4149,4150
3|4150,4151
*|4151,4152
Hct|4153,4156
-|4156,4157
35|4157,4159
.|4159,4160
1|4160,4161
*|4161,4162
<EOL>|4163,4164
MCV|4164,4167
-|4167,4168
81|4168,4170
*|4170,4171
MCH|4172,4175
-|4175,4176
26.2|4176,4180
MCHC|4181,4185
-|4185,4186
32.2|4186,4190
RDW|4191,4194
-|4194,4195
16|4195,4197
.|4197,4198
3|4198,4199
*|4199,4200
RDWSD|4201,4206
-|4206,4207
48|4207,4209
.|4209,4210
3|4210,4211
*|4211,4212
Plt|4213,4216
_|4217,4218
_|4218,4219
_|4219,4220
<EOL>|4220,4221
_|4221,4222
_|4222,4223
_|4223,4224
04|4225,4227
:|4227,4228
02PM|4228,4232
BLOOD|4233,4238
_|4239,4240
_|4240,4241
_|4241,4242
PTT|4243,4246
-|4246,4247
35.8|4247,4251
_|4252,4253
_|4253,4254
_|4254,4255
<EOL>|4255,4256
_|4256,4257
_|4257,4258
_|4258,4259
04|4260,4262
:|4262,4263
02PM|4263,4267
BLOOD|4268,4273
Glucose|4274,4281
-|4281,4282
93|4282,4284
UreaN|4285,4290
-|4290,4291
17|4291,4293
Creat|4294,4299
-|4299,4300
1.1|4300,4303
Na|4304,4306
-|4306,4307
131|4307,4310
*|4310,4311
<EOL>|4312,4313
K|4313,4314
-|4314,4315
3.8|4315,4318
Cl|4319,4321
-|4321,4322
93|4322,4324
*|4324,4325
HCO3|4326,4330
-|4330,4331
27|4331,4333
AnGap|4334,4339
-|4339,4340
15|4340,4342
<EOL>|4342,4343
_|4343,4344
_|4344,4345
_|4345,4346
04|4347,4349
:|4349,4350
02PM|4350,4354
BLOOD|4355,4360
ALT|4361,4364
-|4364,4365
81|4365,4367
*|4367,4368
AST|4369,4372
-|4372,4373
64|4373,4375
*|4375,4376
AlkPhos|4377,4384
-|4384,4385
89|4385,4387
TotBili|4388,4395
-|4395,4396
0.7|4396,4399
<EOL>|4399,4400
_|4400,4401
_|4401,4402
_|4402,4403
04|4404,4406
:|4406,4407
02PM|4407,4411
BLOOD|4412,4417
CK|4418,4420
-|4420,4421
MB|4421,4423
-|4423,4424
3|4424,4425
cTropnT|4426,4433
-|4433,4434
<|4434,4435
0|4435,4436
.|4436,4437
01|4437,4439
proBNP|4440,4446
-|4446,4447
1284|4447,4451
*|4451,4452
<EOL>|4452,4453
_|4453,4454
_|4454,4455
_|4455,4456
04|4457,4459
:|4459,4460
02PM|4460,4464
BLOOD|4465,4470
Albumin|4471,4478
-|4478,4479
4.2|4479,4482
Calcium|4483,4490
-|4490,4491
9.7|4491,4494
Mg|4495,4497
-|4497,4498
2.2|4498,4501
<EOL>|4501,4502
_|4502,4503
_|4503,4504
_|4504,4505
04|4506,4508
:|4508,4509
34PM|4509,4513
BLOOD|4514,4519
D|4520,4521
-|4521,4522
Dimer|4522,4527
-|4527,4528
<|4528,4529
150|4529,4532
<EOL>|4532,4533
_|4533,4534
_|4534,4535
_|4535,4536
04|4537,4539
:|4539,4540
02PM|4540,4544
BLOOD|4545,4550
TSH|4551,4554
-|4554,4555
3.0|4555,4558
<EOL>|4558,4559
<EOL>|4559,4560
DISCHARGE|4560,4569
<EOL>|4569,4570
_|4570,4571
_|4571,4572
_|4572,4573
04|4574,4576
:|4576,4577
04AM|4577,4581
BLOOD|4582,4587
WBC|4588,4591
-|4591,4592
6|4592,4593
.|4593,4594
5|4594,4595
#|4595,4596
RBC|4597,4600
-|4600,4601
4|4601,4602
.|4602,4603
57|4603,4605
*|4605,4606
Hgb|4607,4610
-|4610,4611
12|4611,4613
.|4613,4614
2|4614,4615
*|4615,4616
Hct|4617,4620
-|4620,4621
36|4621,4623
.|4623,4624
8|4624,4625
*|4625,4626
<EOL>|4627,4628
MCV|4628,4631
-|4631,4632
81|4632,4634
*|4634,4635
MCH|4636,4639
-|4639,4640
26.7|4640,4644
MCHC|4645,4649
-|4649,4650
33.2|4650,4654
RDW|4655,4658
-|4658,4659
16|4659,4661
.|4661,4662
4|4662,4663
*|4663,4664
RDWSD|4665,4670
-|4670,4671
47|4671,4673
.|4673,4674
8|4674,4675
*|4675,4676
Plt|4677,4680
_|4681,4682
_|4682,4683
_|4683,4684
<EOL>|4684,4685
_|4685,4686
_|4686,4687
_|4687,4688
04|4689,4691
:|4691,4692
04AM|4692,4696
BLOOD|4697,4702
_|4703,4704
_|4704,4705
_|4705,4706
PTT|4707,4710
-|4710,4711
34.1|4711,4715
_|4716,4717
_|4717,4718
_|4718,4719
<EOL>|4719,4720
_|4720,4721
_|4721,4722
_|4722,4723
04|4724,4726
:|4726,4727
04AM|4727,4731
BLOOD|4732,4737
Glucose|4738,4745
-|4745,4746
113|4746,4749
*|4749,4750
UreaN|4751,4756
-|4756,4757
32|4757,4759
*|4759,4760
Creat|4761,4766
-|4766,4767
1|4767,4768
.|4768,4769
4|4769,4770
*|4770,4771
Na|4772,4774
-|4774,4775
133|4775,4778
<EOL>|4779,4780
K|4780,4781
-|4781,4782
3.9|4782,4785
Cl|4786,4788
-|4788,4789
94|4789,4791
*|4791,4792
HCO3|4793,4797
-|4797,4798
26|4798,4800
AnGap|4801,4806
-|4806,4807
17|4807,4809
<EOL>|4809,4810
_|4810,4811
_|4811,4812
_|4812,4813
04|4814,4816
:|4816,4817
04AM|4817,4821
BLOOD|4822,4827
ALT|4828,4831
-|4831,4832
79|4832,4834
*|4834,4835
AST|4836,4839
-|4839,4840
57|4840,4842
*|4842,4843
AlkPhos|4844,4851
-|4851,4852
83|4852,4854
TotBili|4855,4862
-|4862,4863
0.6|4863,4866
<EOL>|4866,4867
_|4867,4868
_|4868,4869
_|4869,4870
04|4871,4873
:|4873,4874
04AM|4874,4878
BLOOD|4879,4884
Calcium|4885,4892
-|4892,4893
10.0|4893,4897
Phos|4898,4902
-|4902,4903
4.4|4903,4906
Mg|4907,4909
-|4909,4910
2.0|4910,4913
<EOL>|4913,4914
<EOL>|4914,4915
ECHO|4915,4919
_|4920,4921
_|4921,4922
_|4922,4923
<EOL>|4923,4924
The|4924,4927
left|4928,4932
atrium|4933,4939
is|4940,4942
moderately|4943,4953
dilated|4954,4961
.|4961,4962
The|4963,4966
right|4967,4972
atrium|4973,4979
is|4980,4982
<EOL>|4983,4984
moderately|4984,4994
dilated|4995,5002
.|5002,5003
No|5004,5006
atrial|5007,5013
septal|5014,5020
defect|5021,5027
is|5028,5030
seen|5031,5035
by|5036,5038
2D|5039,5041
or|5042,5044
<EOL>|5045,5046
color|5046,5051
Doppler|5052,5059
.|5059,5060
Left|5061,5065
ventricular|5066,5077
wall|5078,5082
thicknesses|5083,5094
and|5095,5098
cavity|5099,5105
size|5106,5110
<EOL>|5111,5112
are|5112,5115
normal|5116,5122
.|5122,5123
There|5124,5129
is|5130,5132
mild|5133,5137
regional|5138,5146
left|5147,5151
ventricular|5152,5163
systolic|5164,5172
<EOL>|5173,5174
dysfunction|5174,5185
with|5186,5190
hypokinesis|5191,5202
of|5203,5205
the|5206,5209
mid-anterior|5210,5222
and|5223,5226
mid-distal|5227,5237
<EOL>|5238,5239
inferior|5239,5247
wall|5248,5252
.|5252,5253
The|5254,5257
estimated|5258,5267
cardiac|5268,5275
index|5276,5281
is|5282,5284
normal|5285,5291
<EOL>|5292,5293
(|5293,5294
>|5294,5295
=|5295,5296
2.5|5296,5299
L|5299,5300
/|5300,5301
min|5301,5304
/|5304,5305
m2|5305,5307
)|5307,5308
.|5308,5309
Doppler|5310,5317
parameters|5318,5328
are|5329,5332
indeterminate|5333,5346
for|5347,5350
left|5351,5355
<EOL>|5356,5357
ventricular|5357,5368
diastolic|5369,5378
function|5379,5387
.|5387,5388
The|5389,5392
right|5393,5398
ventricular|5399,5410
cavity|5411,5417
is|5418,5420
<EOL>|5421,5422
mildly|5422,5428
dilated|5429,5436
with|5437,5441
depressed|5442,5451
free|5452,5456
wall|5457,5461
contractility|5462,5475
(|5476,5477
RV|5477,5479
free|5480,5484
<EOL>|5485,5486
wall|5486,5490
is|5491,5493
not|5494,5497
well|5498,5502
seen|5503,5507
)|5507,5508
.|5508,5509
The|5510,5513
aortic|5514,5520
valve|5521,5526
leaflets|5527,5535
(|5536,5537
3|5537,5538
)|5538,5539
are|5540,5543
mildly|5544,5550
<EOL>|5551,5552
thickened|5552,5561
but|5562,5565
aortic|5566,5572
stenosis|5573,5581
is|5582,5584
not|5585,5588
present|5589,5596
.|5596,5597
The|5598,5601
mitral|5602,5608
valve|5609,5614
<EOL>|5615,5616
leaflets|5616,5624
are|5625,5628
mildly|5629,5635
thickened|5636,5645
.|5645,5646
There|5647,5652
is|5653,5655
no|5656,5658
mitral|5659,5665
valve|5666,5671
<EOL>|5672,5673
prolapse|5673,5681
.|5681,5682
Trivial|5683,5690
mitral|5691,5697
regurgitation|5698,5711
is|5712,5714
seen|5715,5719
.|5719,5720
The|5721,5724
tricuspid|5725,5734
<EOL>|5735,5736
valve|5736,5741
leaflets|5742,5750
are|5751,5754
mildly|5755,5761
thickened|5762,5771
.|5771,5772
Moderate|5773,5781
[|5782,5783
2|5783,5784
+|5784,5785
]|5785,5786
tricuspid|5787,5796
<EOL>|5797,5798
regurgitation|5798,5811
is|5812,5814
seen|5815,5819
.|5819,5820
There|5821,5826
is|5827,5829
moderate|5830,5838
pulmonary|5839,5848
artery|5849,5855
<EOL>|5856,5857
systolic|5857,5865
hypertension|5866,5878
.|5878,5879
The|5880,5883
pulmonic|5884,5892
valve|5893,5898
leaflets|5899,5907
are|5908,5911
<EOL>|5912,5913
thickened|5913,5922
.|5922,5923
There|5924,5929
is|5930,5932
no|5933,5935
pericardial|5936,5947
effusion|5948,5956
.|5956,5957
<EOL>|5958,5959
<EOL>|5959,5960
IMPRESSION|5960,5970
:|5970,5971
Mild|5972,5976
regional|5977,5985
left|5986,5990
ventricular|5991,6002
dysfunction|6003,6014
c|6015,6016
/|6016,6017
w|6017,6018
<EOL>|6019,6020
multivessel|6020,6031
CAD|6032,6035
,|6035,6036
with|6037,6041
overall|6042,6049
mildly|6050,6056
depressed|6057,6066
global|6067,6073
systolic|6074,6082
<EOL>|6083,6084
function|6084,6092
.|6092,6093
Mildly|6094,6100
dilated|6101,6108
right|6109,6114
ventricle|6115,6124
with|6125,6129
depressed|6130,6139
free|6140,6144
<EOL>|6145,6146
wall|6146,6150
systolic|6151,6159
function|6160,6168
.|6168,6169
Moderate|6170,6178
tricuspid|6179,6188
regurgitation|6189,6202
with|6203,6207
<EOL>|6208,6209
moderate|6209,6217
pulmonary|6218,6227
hypertension|6228,6240
.|6240,6241
<EOL>|6243,6244
<EOL>|6245,6246
Mr.|6269,6272
_|6273,6274
_|6274,6275
_|6275,6276
is|6277,6279
an|6280,6282
_|6283,6284
_|6284,6285
_|6285,6286
year|6287,6291
old|6292,6295
gentleman|6296,6305
with|6306,6310
history|6311,6318
of|6319,6321
CAD|6322,6325
<EOL>|6326,6327
(|6327,6328
s|6328,6329
/|6329,6330
p|6330,6331
CABG|6332,6336
and|6337,6340
PCI|6341,6344
)|6344,6345
,|6345,6346
pAF|6347,6350
,|6350,6351
PAH|6352,6355
,|6355,6356
diastolic|6357,6366
CHF|6367,6370
who|6371,6374
presents|6375,6383
with|6384,6388
<EOL>|6389,6390
weight|6390,6396
gain|6397,6401
,|6401,6402
leg|6403,6406
swelling|6407,6415
and|6416,6419
new|6420,6423
evidence|6424,6432
of|6433,6435
right|6436,6441
ventricle|6442,6451
<EOL>|6452,6453
dilation|6453,6461
concerning|6462,6472
for|6473,6476
acute|6477,6482
on|6483,6485
chronic|6486,6493
heart|6494,6499
failure|6500,6507
<EOL>|6508,6509
exacerbation|6509,6521
.|6521,6522
<EOL>|6524,6525
<EOL>|6525,6526
#|6526,6527
Acute|6527,6532
on|6533,6535
Chronic|6536,6543
Diastolic|6544,6553
Heart|6554,6559
Failure|6560,6567
Exacerbation|6568,6580
:|6580,6581
with|6582,6586
<EOL>|6587,6588
component|6588,6597
of|6598,6600
RV|6601,6603
failure|6604,6611
by|6612,6614
report|6615,6621
of|6622,6624
OSH|6625,6628
echo|6629,6633
.|6633,6634
Likely|6636,6642
primary|6643,6650
<EOL>|6651,6652
process|6652,6659
is|6660,6662
lung|6663,6667
disease|6668,6675
causing|6676,6683
elevated|6684,6692
RV|6693,6695
pressures|6696,6705
and|6706,6709
<EOL>|6710,6711
subsequent|6711,6721
poor|6722,6726
filling|6727,6734
of|6735,6737
LV|6738,6740
.|6740,6741
He|6743,6745
diuresed|6746,6754
quite|6755,6760
well|6761,6765
with|6766,6770
20|6771,6773
<EOL>|6774,6775
IV|6775,6777
Lasix|6778,6783
which|6784,6789
is|6790,6792
consistent|6793,6803
with|6804,6808
RV|6809,6811
failure|6812,6819
.|6819,6820
Started|6822,6829
on|6830,6832
<EOL>|6833,6834
torsemide|6834,6843
10|6844,6846
daily|6847,6852
but|6853,6856
this|6857,6861
is|6862,6864
likely|6865,6871
too|6872,6875
aggressive|6876,6886
.|6886,6887
We|6889,6891
<EOL>|6892,6893
obtained|6893,6901
an|6902,6904
echo|6905,6909
but|6910,6913
read|6914,6918
PND|6919,6922
at|6923,6925
time|6926,6930
of|6931,6933
discharge|6934,6943
.|6943,6944
We|6946,6948
sent|6949,6953
him|6954,6957
<EOL>|6958,6959
home|6959,6963
on|6964,6966
a|6967,6968
diuretic|6969,6977
regimen|6978,6985
on|6986,6988
torsemide|6989,6998
5|6999,7000
mg|7001,7003
daily|7004,7009
(|7010,7011
and|7011,7014
<EOL>|7015,7016
discontinued|7016,7028
home|7029,7033
triamterene|7034,7045
-|7045,7046
HCTZ|7046,7050
)|7050,7051
.|7051,7052
Close|7054,7059
follow|7060,7066
up|7067,7069
with|7070,7074
Dr|7075,7077
.|7077,7078
<EOL>|7079,7080
_|7080,7081
_|7081,7082
_|7082,7083
ensured|7084,7091
.|7091,7092
<EOL>|7092,7093
<EOL>|7093,7094
#|7094,7095
Elevated|7095,7103
Transaminases|7104,7117
:|7117,7118
Patient|7120,7127
with|7128,7132
mildly|7133,7139
elevated|7140,7148
AST|7149,7152
and|7153,7156
<EOL>|7157,7158
ALT|7158,7161
.|7161,7162
Most|7163,7167
likely|7168,7174
etiologies|7175,7185
in|7186,7188
this|7189,7193
patient|7194,7201
include|7202,7209
amiodarone|7210,7220
<EOL>|7221,7222
toxicity|7222,7230
and|7231,7234
congestive|7235,7245
hepatopathy|7246,7257
.|7257,7258
Encouraged|7260,7270
outpatient|7271,7281
<EOL>|7282,7283
trending|7283,7291
.|7291,7292
<EOL>|7293,7294
<EOL>|7294,7295
#|7295,7296
Pulmonary|7296,7305
disease|7306,7313
:|7313,7314
patient|7315,7322
with|7323,7327
extensive|7328,7337
emphysema|7338,7347
on|7348,7350
CTA|7351,7354
<EOL>|7355,7356
though|7356,7362
patient|7363,7370
has|7371,7374
no|7375,7377
history|7378,7385
of|7386,7388
smoking|7389,7396
.|7396,7397
As|7399,7401
this|7402,7406
may|7407,7410
be|7411,7413
<EOL>|7414,7415
driving|7415,7422
R|7423,7424
heart|7425,7430
failure|7431,7438
,|7438,7439
Dr.|7440,7443
_|7444,7445
_|7445,7446
_|7446,7447
requested|7448,7457
pulmonology|7458,7469
<EOL>|7470,7471
consult|7471,7478
prior|7479,7484
to|7485,7487
discharge|7488,7497
but|7498,7501
patient|7502,7509
was|7510,7513
insistent|7514,7523
on|7524,7526
leaving|7527,7534
.|7534,7535
<EOL>|7536,7537
Instead|7538,7545
scheduled|7546,7555
outpatient|7556,7566
appointment|7567,7578
.|7578,7579
<EOL>|7580,7581
<EOL>|7582,7583
#|7583,7584
Atrial|7584,7590
Fibrillation|7591,7603
:|7603,7604
Continue|7605,7613
home|7614,7618
amiodarone|7619,7629
200mg|7630,7635
daily|7636,7641
,|7641,7642
<EOL>|7643,7644
Apixaban|7644,7652
5mg|7653,7656
BID|7657,7660
<EOL>|7662,7663
<EOL>|7663,7664
#|7664,7665
CAD|7665,7668
:|7668,7669
Continue|7670,7678
ASA|7679,7682
81mg|7683,7687
,|7687,7688
rosuvastatin|7689,7701
40mg|7702,7706
qHS|7707,7710
<EOL>|7712,7713
<EOL>|7713,7714
#|7714,7715
HTN|7715,7718
:|7718,7719
continue|7720,7728
home|7729,7733
losartan|7734,7742
25mg|7743,7747
qD|7748,7750
.|7750,7751
<EOL>|7751,7752
<EOL>|7752,7753
TRANSITIONAL|7753,7765
ISSUES|7766,7772
<EOL>|7772,7773
[|7773,7774
]|7774,7775
New|7776,7779
medication|7780,7790
:|7790,7791
Torsemide|7792,7801
5|7802,7803
mg|7804,7806
daily|7807,7812
<EOL>|7812,7813
[|7813,7814
]|7814,7815
Discontinued|7816,7828
triamterene|7829,7840
/|7840,7841
HCTZ|7841,7845
in|7846,7848
favor|7849,7854
of|7855,7857
above|7858,7863
<EOL>|7863,7864
[|7864,7865
]|7865,7866
LFTs|7867,7871
mild|7872,7876
elevated|7877,7885
in|7886,7888
house|7889,7894
;|7894,7895
consider|7896,7904
possible|7905,7913
<EOL>|7914,7915
discontinuing|7915,7928
/|7928,7929
changing|7929,7937
amiodarone|7938,7948
<EOL>|7948,7949
[|7949,7950
]|7950,7951
Please|7952,7958
check|7959,7964
LFT|7965,7968
's|7968,7970
and|7971,7974
Creatinine|7975,7985
at|7986,7988
follow|7989,7995
up|7996,7998
appointment|7999,8010
as|8011,8013
<EOL>|8014,8015
these|8015,8020
were|8021,8025
elevated|8026,8034
while|8035,8040
hospitalized|8041,8053
<EOL>|8053,8054
[|8054,8055
]|8055,8056
Follow|8057,8063
up|8064,8066
appointment|8067,8078
with|8079,8083
cardiology|8084,8094
,|8094,8095
Dr.|8096,8099
_|8100,8101
_|8101,8102
_|8102,8103
<EOL>|8103,8104
[|8104,8105
]|8105,8106
Follow|8107,8113
up|8114,8116
appointment|8117,8128
with|8129,8133
pulmonology|8134,8145
<EOL>|8145,8146
[|8146,8147
]|8147,8148
Follow|8149,8155
up|8156,8158
appointment|8159,8170
with|8171,8175
PCP|8176,8179
<EOL>|8179,8180
<EOL>|8180,8181
*|8181,8182
*|8182,8183
*|8183,8184
Discharge|8184,8193
weight|8194,8200
63.1|8201,8205
kg|8206,8208
*|8208,8209
*|8209,8210
*|8210,8211
<EOL>|8213,8214
<EOL>|8215,8216
Medications|8216,8227
on|8228,8230
Admission|8231,8240
:|8240,8241
<EOL>|8241,8242
The|8242,8245
Preadmission|8246,8258
Medication|8259,8269
list|8270,8274
is|8275,8277
accurate|8278,8286
and|8287,8290
complete|8291,8299
.|8299,8300
<EOL>|8300,8301
1.|8301,8303
Amiodarone|8304,8314
200|8315,8318
mg|8319,8321
PO|8322,8324
DAILY|8325,8330
<EOL>|8331,8332
2.|8332,8334
Apixaban|8335,8343
5|8344,8345
mg|8346,8348
PO|8349,8351
BID|8352,8355
<EOL>|8356,8357
3.|8357,8359
Aspirin|8360,8367
81|8368,8370
mg|8371,8373
PO|8374,8376
DAILY|8377,8382
<EOL>|8383,8384
4.|8384,8386
Docusate|8387,8395
Sodium|8396,8402
100|8403,8406
mg|8407,8409
PO|8410,8412
BID|8413,8416
<EOL>|8417,8418
5.|8418,8420
Losartan|8421,8429
Potassium|8430,8439
25|8440,8442
mg|8443,8445
PO|8446,8448
DAILY|8449,8454
<EOL>|8455,8456
6.|8456,8458
Omeprazole|8459,8469
10|8470,8472
mg|8473,8475
PO|8476,8478
DAILY|8479,8484
<EOL>|8485,8486
7.|8486,8488
Triamterene|8489,8500
-|8500,8501
HCTZ|8501,8505
(|8506,8507
37.5|8507,8511
/|8511,8512
25|8512,8514
)|8514,8515
1|8516,8517
CAP|8518,8521
PO|8522,8524
DAILY|8525,8530
<EOL>|8531,8532
8.|8532,8534
Senna|8535,8540
17.2|8541,8545
mg|8546,8548
PO|8549,8551
HS|8552,8554
<EOL>|8555,8556
9.|8556,8558
Align|8559,8564
(|8565,8566
bifidobacterium|8566,8581
infantis|8582,8590
)|8590,8591
4|8592,8593
mg|8594,8596
oral|8597,8601
DAILY|8602,8607
<EOL>|8608,8609
10.|8609,8612
coenzyme|8613,8621
Q10|8622,8625
100|8626,8629
mg|8630,8632
oral|8633,8637
DAILY|8638,8643
<EOL>|8644,8645
11.|8645,8648
Rosuvastatin|8649,8661
Calcium|8662,8669
40|8670,8672
mg|8673,8675
PO|8676,8678
QPM|8679,8682
<EOL>|8683,8684
12.|8684,8687
Vitamin|8688,8695
D|8696,8697
1000|8698,8702
UNIT|8703,8707
PO|8708,8710
DAILY|8711,8716
<EOL>|8717,8718
13.|8718,8721
Tamsulosin|8722,8732
0.4|8733,8736
mg|8737,8739
PO|8740,8742
QHS|8743,8746
<EOL>|8747,8748
<EOL>|8748,8749
<EOL>|8750,8751
Discharge|8751,8760
Medications|8761,8772
:|8772,8773
<EOL>|8773,8774
1.|8774,8776
Amiodarone|8777,8787
200|8788,8791
mg|8792,8794
PO|8795,8797
DAILY|8798,8803
<EOL>|8804,8805
2.|8805,8807
Apixaban|8808,8816
5|8817,8818
mg|8819,8821
PO|8822,8824
BID|8825,8828
<EOL>|8829,8830
3.|8830,8832
Aspirin|8833,8840
81|8841,8843
mg|8844,8846
PO|8847,8849
DAILY|8850,8855
<EOL>|8856,8857
4.|8857,8859
Docusate|8860,8868
Sodium|8869,8875
100|8876,8879
mg|8880,8882
PO|8883,8885
BID|8886,8889
<EOL>|8890,8891
5.|8891,8893
Losartan|8894,8902
Potassium|8903,8912
25|8913,8915
mg|8916,8918
PO|8919,8921
DAILY|8922,8927
<EOL>|8928,8929
6.|8929,8931
Rosuvastatin|8932,8944
Calcium|8945,8952
40|8953,8955
mg|8956,8958
PO|8959,8961
QPM|8962,8965
<EOL>|8966,8967
7.|8967,8969
Senna|8970,8975
17.2|8976,8980
mg|8981,8983
PO|8984,8986
HS|8987,8989
<EOL>|8990,8991
RX|8991,8993
*|8994,8995
sennosides|8995,9005
[|9006,9007
senna|9007,9012
]|9012,9013
8.6|9014,9017
mg|9018,9020
1|9021,9022
capsule|9023,9030
by|9031,9033
mouth|9034,9039
once|9040,9044
a|9045,9046
day|9047,9050
Disp|9051,9055
<EOL>|9056,9057
#|9057,9058
*|9058,9059
30|9059,9061
Capsule|9062,9069
Refills|9070,9077
:|9077,9078
*|9078,9079
0|9079,9080
<EOL>|9080,9081
8.|9081,9083
Vitamin|9084,9091
D|9092,9093
1000|9094,9098
UNIT|9099,9103
PO|9104,9106
DAILY|9107,9112
<EOL>|9113,9114
9.|9114,9116
Torsemide|9117,9126
5|9127,9128
mg|9129,9131
PO|9132,9134
DAILY|9135,9140
<EOL>|9141,9142
RX|9142,9144
*|9145,9146
torsemide|9146,9155
5|9156,9157
mg|9158,9160
1|9161,9162
tablet|9163,9169
(|9169,9170
s|9170,9171
)|9171,9172
by|9173,9175
mouth|9176,9181
once|9182,9186
a|9187,9188
day|9189,9192
Disp|9193,9197
#|9198,9199
*|9199,9200
30|9200,9202
<EOL>|9203,9204
Tablet|9204,9210
Refills|9211,9218
:|9218,9219
*|9219,9220
0|9220,9221
<EOL>|9221,9222
10.|9222,9225
Align|9226,9231
(|9232,9233
bifidobacterium|9233,9248
infantis|9249,9257
)|9257,9258
4|9259,9260
mg|9261,9263
oral|9264,9268
DAILY|9269,9274
<EOL>|9275,9276
11.|9276,9279
coenzyme|9280,9288
Q10|9289,9292
100|9293,9296
mg|9297,9299
oral|9300,9304
DAILY|9305,9310
<EOL>|9311,9312
12.|9312,9315
Omeprazole|9316,9326
10|9327,9329
mg|9330,9332
PO|9333,9335
DAILY|9336,9341
<EOL>|9342,9343
13.|9343,9346
Tamsulosin|9347,9357
0.4|9358,9361
mg|9362,9364
PO|9365,9367
QHS|9368,9371
<EOL>|9372,9373
<EOL>|9373,9374
<EOL>|9375,9376
Discharge|9376,9385
Disposition|9386,9397
:|9397,9398
<EOL>|9398,9399
Home|9399,9403
<EOL>|9403,9404
<EOL>|9405,9406
Discharge|9406,9415
Diagnosis|9416,9425
:|9425,9426
<EOL>|9426,9427
Primary|9427,9434
:|9434,9435
<EOL>|9435,9436
Acute|9436,9441
on|9442,9444
chronic|9445,9452
diastolic|9453,9462
congestive|9463,9473
heart|9474,9479
failure|9480,9487
<EOL>|9487,9488
Cor|9488,9491
pulmonale|9492,9501
<EOL>|9501,9502
<EOL>|9502,9503
Secondary|9503,9512
:|9512,9513
<EOL>|9513,9514
Pulmonary|9514,9523
hypertension|9524,9536
<EOL>|9536,9537
Paroxysmal|9537,9547
atrial|9548,9554
fibrillation|9555,9567
<EOL>|9567,9568
Hyponatremia|9568,9580
<EOL>|9580,9581
<EOL>|9581,9582
<EOL>|9583,9584
Mental|9605,9611
Status|9612,9618
:|9618,9619
Clear|9620,9625
and|9626,9629
coherent|9630,9638
.|9638,9639
<EOL>|9639,9640
Level|9640,9645
of|9646,9648
Consciousness|9649,9662
:|9662,9663
Alert|9664,9669
and|9670,9673
interactive|9674,9685
.|9685,9686
<EOL>|9686,9687
Activity|9687,9695
Status|9696,9702
:|9702,9703
Ambulatory|9704,9714
-|9715,9716
Independent|9717,9728
.|9728,9729
<EOL>|9729,9730
<EOL>|9730,9731
<EOL>|9732,9733
Dear|9757,9761
Mr.|9762,9765
_|9766,9767
_|9767,9768
_|9768,9769
,|9769,9770
<EOL>|9770,9771
<EOL>|9771,9772
You|9772,9775
were|9776,9780
hospitalized|9781,9793
for|9794,9797
progressive|9798,9809
leg|9810,9813
swelling|9814,9822
over|9823,9827
the|9828,9831
past|9832,9836
<EOL>|9837,9838
week|9838,9842
and|9843,9846
a|9847,9848
half|9849,9853
.|9853,9854
We|9856,9858
started|9859,9866
you|9867,9870
on|9871,9873
a|9874,9875
new|9876,9879
medication|9880,9890
here|9891,9895
that|9896,9900
<EOL>|9901,9902
should|9902,9908
help|9909,9913
prevent|9914,9921
this|9922,9926
from|9927,9931
happening|9932,9941
.|9941,9942
Of|9944,9946
note|9947,9951
,|9951,9952
Dr.|9953,9956
_|9957,9958
_|9958,9959
_|9959,9960
was|9961,9964
<EOL>|9965,9966
concerned|9966,9975
about|9976,9981
a|9982,9983
clot|9984,9988
in|9989,9991
your|9992,9996
lungs|9997,10002
,|10002,10003
but|10004,10007
our|10008,10011
scans|10012,10017
showed|10018,10024
NO|10025,10027
<EOL>|10028,10029
clot|10029,10033
.|10033,10034
With|10036,10040
this|10041,10045
news|10046,10050
,|10050,10051
you|10052,10055
were|10056,10060
discharged|10061,10071
home|10072,10076
with|10077,10081
PCP|10082,10085
and|10086,10089
<EOL>|10090,10091
cardiology|10091,10101
follow|10102,10108
up|10109,10111
.|10111,10112
<EOL>|10112,10113
<EOL>|10113,10114
Please|10114,10120
continue|10121,10129
to|10130,10132
take|10133,10137
your|10138,10142
torsemide|10143,10152
in|10153,10155
order|10156,10161
to|10162,10164
maintain|10165,10173
your|10174,10178
<EOL>|10179,10180
weight|10180,10186
.|10186,10187
Please|10188,10194
weight|10195,10201
yourself|10202,10210
everyday|10211,10219
and|10220,10223
call|10224,10228
your|10229,10233
<EOL>|10234,10235
cardiologist|10235,10247
if|10248,10250
you|10251,10254
weight|10255,10261
changes|10262,10269
by|10270,10272
three|10273,10278
pounds|10279,10285
.|10285,10286
<EOL>|10286,10287
<EOL>|10287,10288
You|10288,10291
also|10292,10296
have|10297,10301
"|10302,10303
pulmonary|10303,10312
hypertension|10313,10325
,|10325,10326
"|10326,10327
which|10328,10333
may|10334,10337
be|10338,10340
due|10341,10344
to|10345,10347
your|10348,10352
<EOL>|10353,10354
underlying|10354,10364
lung|10365,10369
disease|10370,10377
.|10377,10378
Amiodarone|10379,10389
can|10390,10393
also|10394,10398
cause|10399,10404
lung|10405,10409
changes|10410,10417
<EOL>|10418,10419
and|10419,10422
we|10423,10425
recommend|10426,10435
following|10436,10445
up|10446,10448
with|10449,10453
the|10454,10457
lung|10458,10462
doctors|10463,10470
as|10471,10473
_|10474,10475
_|10475,10476
_|10476,10477
<EOL>|10478,10479
outpatient|10479,10489
to|10490,10492
see|10493,10496
if|10497,10499
this|10500,10504
may|10505,10508
be|10509,10511
contributing|10512,10524
.|10524,10525
<EOL>|10526,10527
<EOL>|10527,10528
It|10528,10530
was|10531,10534
a|10535,10536
pleasure|10537,10545
taking|10546,10552
care|10553,10557
of|10558,10560
you|10561,10564
!|10564,10565
<EOL>|10565,10566
Your|10566,10570
_|10571,10572
_|10572,10573
_|10573,10574
team|10575,10579
<EOL>|10579,10580
<EOL>|10581,10582
Followup|10582,10590
Instructions|10591,10603
:|10603,10604
<EOL>|10604,10605
_|10605,10606
_|10606,10607
_|10607,10608
<EOL>|10608,10609

