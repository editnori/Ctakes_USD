 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
SURGERY|155,162
<EOL>|162,163
<EOL>|164,165
Codeine|177,184
/|185,186
Augmentin|187,196
/|197,198
Topamax|199,206
<EOL>|206,207
<EOL>|208,209
Attending|209,218
:|218,219
_|220,221
_|221,222
_|222,223
<EOL>|223,224
<EOL>|225,226
_|226,227
_|227,228
_|228,229
Complaint|230,239
:|239,240
<EOL>|240,241
left|241,245
breast|246,252
swelling|253,261
and|262,265
pain|266,270
<EOL>|270,271
<EOL>|272,273
Major|273,278
Surgical|279,287
or|288,290
Invasive|291,299
Procedure|300,309
:|309,310
<EOL>|310,311
Evacuation|311,321
of|322,324
hematoma|325,333
<EOL>|334,335
<EOL>|335,336
<EOL>|337,338
_|366,367
_|367,368
_|368,369
woman|370,375
on|376,378
anticoagulation|379,394
with|395,399
L|400,401
breast|402,408
IDC|409,412
Grade|413,418
3|419,420
<EOL>|421,422
now|422,425
s|426,427
/|427,428
p|428,429
L|430,431
breast|432,438
lumpectomy|439,449
and|450,453
SLNB|454,458
with|459,463
left|464,468
breast|469,475
swelling|476,484
<EOL>|485,486
and|486,489
pain|490,494
concerning|495,505
for|506,509
a|510,511
hematoma|512,520
.|520,521
<EOL>|522,523
<EOL>|524,525
Dyslipidemia|547,559
,|559,560
varicose|561,569
veins|570,575
(|576,577
R|577,578
>|578,579
L|579,580
)|580,581
s|582,583
/|583,584
p|584,585
ligation|586,594
,|594,595
COPD|596,600
,|600,601
OSA|602,605
<EOL>|606,607
(|607,608
+|608,609
CPap|609,613
)|613,614
,|614,615
recent|616,622
URI|623,626
(|627,628
received|628,636
course|637,643
of|644,646
Zithromax|647,656
)|656,657
,|657,658
bilateral|659,668
<EOL>|669,670
PEs|670,673
(|674,675
_|675,676
_|676,677
_|677,678
)|678,679
,|679,680
antiphospholipid|681,697
antibody|698,706
syndrome|707,715
(|716,717
on|717,719
lifelong|720,728
<EOL>|729,730
anticoagulation|730,745
)|745,746
,|746,747
T2DM|748,752
(|753,754
last|754,758
A1C|759,762
6.2|763,766
on|767,769
_|770,771
_|771,772
_|772,773
,|773,774
cerebral|775,783
<EOL>|784,785
aneurysm|785,793
(|794,795
followed|795,803
by|804,806
Dr.|807,810
_|811,812
_|812,813
_|813,814
,|814,815
unchanged|816,825
)|825,826
,|826,827
GERD|828,832
,|832,833
<EOL>|834,835
diverticulosis|835,849
,|849,850
h|851,852
/|852,853
o|853,854
colon|855,860
polyps|861,867
,|867,868
depression|869,879
,|879,880
s|881,882
/|882,883
p|883,884
right|885,890
CMC|891,894
<EOL>|895,896
joint|896,901
arthroplasty|902,914
,|914,915
b|916,917
/|917,918
l|918,919
rotator|920,927
cuff|928,932
repair|933,939
,|939,940
excision|941,949
right|950,955
_|956,957
_|957,958
_|958,959
<EOL>|960,961
digit|961,966
mass|967,971
,|971,972
CCY|973,976
w|977,978
/|978,979
stone|979,984
&|985,986
pancreatic|987,997
duct|998,1002
exploration|1003,1014
(|1015,1016
_|1016,1017
_|1017,1018
_|1018,1019
)|1019,1020
,|1020,1021
<EOL>|1022,1023
hysterectomy|1023,1035
,|1035,1036
tonsillectomy|1037,1050
<EOL>|1051,1052
<EOL>|1053,1054
:|1068,1069
<EOL>|1069,1070
_|1070,1071
_|1071,1072
_|1072,1073
<EOL>|1073,1074
:|1088,1089
<EOL>|1089,1090
No|1090,1092
family|1093,1099
hx|1100,1102
of|1103,1105
DVT|1106,1109
or|1110,1112
PE|1113,1115
,|1115,1116
two|1117,1120
sisters|1121,1128
have|1129,1133
atrial|1134,1140
fibrillation|1141,1153
.|1153,1154
<EOL>|1155,1156
<EOL>|1157,1158
<EOL>|1158,1159
<EOL>|1160,1161
<EOL>|1175,1176
VS|1191,1193
:|1193,1194
_|1195,1196
_|1196,1197
_|1197,1198
0313|1199,1203
Temp|1204,1208
:|1208,1209
98.2|1210,1214
PO|1215,1217
BP|1218,1220
:|1220,1221
98|1222,1224
/|1224,1225
62|1225,1227
HR|1228,1230
:|1230,1231
79|1232,1234
RR|1235,1237
:|1237,1238
18|1239,1241
O2|1242,1244
sat|1245,1248
:|1248,1249
<EOL>|1249,1250
95|1250,1252
%|1252,1253
O2|1254,1256
delivery|1257,1265
:|1265,1266
RA|1267,1269
<EOL>|1270,1271
GEN|1271,1274
:|1274,1275
NAD|1276,1279
,|1279,1280
pleasant|1281,1289
,|1289,1290
conversant|1291,1301
<EOL>|1302,1303
HEENT|1303,1308
:|1308,1309
NCAT|1310,1314
,|1314,1315
EOMI|1316,1320
,|1320,1321
sclera|1322,1328
anicteric|1329,1338
<EOL>|1338,1339
CV|1339,1341
:|1341,1342
RRR|1343,1346
<EOL>|1346,1347
PULM|1347,1351
:|1351,1352
no|1353,1355
increased|1356,1365
work|1366,1370
of|1371,1373
breathing|1374,1383
,|1383,1384
comfortable|1385,1396
on|1397,1399
RA|1400,1402
<EOL>|1402,1403
BREAST|1403,1409
:|1409,1410
L|1411,1412
breast|1413,1419
with|1420,1424
dependent|1425,1434
ecchymosis|1435,1445
,|1445,1446
mildly|1447,1453
ttp|1454,1457
inferior|1458,1466
<EOL>|1466,1467
breast|1467,1473
,|1473,1474
incision|1475,1483
C|1484,1485
/|1485,1486
D|1486,1487
/|1487,1488
I|1488,1489
.|1489,1490
JP|1491,1493
drain|1494,1499
with|1500,1504
serosanguineous|1505,1520
output|1521,1527
.|1527,1528
<EOL>|1529,1530
ABD|1530,1533
:|1533,1534
soft|1535,1539
,|1539,1540
non-tender|1541,1551
,|1551,1552
non-distended|1553,1566
,|1566,1567
no|1568,1570
masses|1571,1577
or|1578,1580
hernia|1581,1587
<EOL>|1587,1588
EXT|1588,1591
:|1591,1592
Warm|1593,1597
,|1597,1598
well|1599,1603
-|1603,1604
perfused|1604,1612
,|1612,1613
no|1614,1616
edema|1617,1622
,|1622,1623
no|1624,1626
tenderness|1627,1637
<EOL>|1638,1639
NEURO|1639,1644
:|1644,1645
A|1646,1647
&|1647,1648
Ox3|1648,1651
,|1651,1652
no|1653,1655
focal|1656,1661
neurologic|1662,1672
deficits|1673,1681
<EOL>|1681,1682
PSYCH|1682,1687
:|1687,1688
normal|1689,1695
judgment|1696,1704
/|1704,1705
insight|1705,1712
,|1712,1713
normal|1714,1720
memory|1721,1727
,|1727,1728
normal|1729,1735
<EOL>|1736,1737
mood|1737,1741
/|1741,1742
affect|1742,1748
<EOL>|1748,1749
<EOL>|1750,1751
Pertinent|1751,1760
Results|1761,1768
:|1768,1769
<EOL>|1769,1770
_|1770,1771
_|1771,1772
_|1772,1773
07|1774,1776
:|1776,1777
33AM|1777,1781
BLOOD|1782,1787
WBC|1788,1791
-|1791,1792
4.8|1792,1795
RBC|1796,1799
-|1799,1800
2|1800,1801
.|1801,1802
86|1802,1804
*|1804,1805
Hgb|1806,1809
-|1809,1810
8|1810,1811
.|1811,1812
6|1812,1813
*|1813,1814
Hct|1815,1818
-|1818,1819
27|1819,1821
.|1821,1822
2|1822,1823
*|1823,1824
<EOL>|1825,1826
MCV|1826,1829
-|1829,1830
95|1830,1832
MCH|1833,1836
-|1836,1837
30.1|1837,1841
MCHC|1842,1846
-|1846,1847
31|1847,1849
.|1849,1850
6|1850,1851
*|1851,1852
RDW|1853,1856
-|1856,1857
14.7|1857,1861
RDWSD|1862,1867
-|1867,1868
48|1868,1870
.|1870,1871
7|1871,1872
*|1872,1873
Plt|1874,1877
_|1878,1879
_|1879,1880
_|1880,1881
<EOL>|1881,1882
_|1882,1883
_|1883,1884
_|1884,1885
07|1886,1888
:|1888,1889
33AM|1889,1893
BLOOD|1894,1899
_|1900,1901
_|1901,1902
_|1902,1903
PTT|1904,1907
-|1907,1908
26.2|1908,1912
_|1913,1914
_|1914,1915
_|1915,1916
<EOL>|1916,1917
_|1917,1918
_|1918,1919
_|1919,1920
07|1921,1923
:|1923,1924
33AM|1924,1928
BLOOD|1929,1934
Glucose|1935,1942
-|1942,1943
130|1943,1946
*|1946,1947
UreaN|1948,1953
-|1953,1954
7|1954,1955
Creat|1956,1961
-|1961,1962
0.8|1962,1965
Na|1966,1968
-|1968,1969
141|1969,1972
<EOL>|1973,1974
K|1974,1975
-|1975,1976
4.2|1976,1979
Cl|1980,1982
-|1982,1983
101|1983,1986
HCO3|1987,1991
-|1991,1992
31|1992,1994
AnGap|1995,2000
-|2000,2001
9|2001,2002
*|2002,2003
<EOL>|2003,2004
_|2004,2005
_|2005,2006
_|2006,2007
07|2008,2010
:|2010,2011
33AM|2011,2015
BLOOD|2016,2021
Calcium|2022,2029
-|2029,2030
8|2030,2031
.|2031,2032
2|2032,2033
*|2033,2034
Phos|2035,2039
-|2039,2040
3.8|2040,2043
Mg|2044,2046
-|2046,2047
2.0|2047,2050
<EOL>|2050,2051
<EOL>|2051,2052
EXAMINATION|2052,2063
:|2063,2064
CTA|2066,2069
CHEST|2070,2075
WITH|2076,2080
CONTRAST|2081,2089
<EOL>|2091,2092
COMPARISON|2092,2102
:|2102,2103
Chest|2105,2110
CT|2111,2113
dated|2114,2119
_|2120,2121
_|2121,2122
_|2122,2123
.|2123,2124
<EOL>|2125,2126
<EOL>|2128,2129
:|2137,2138
<EOL>|2140,2141
<EOL>|2143,2144
HEART|2144,2149
AND|2150,2153
VASCULATURE|2154,2165
:|2165,2166
There|2167,2172
is|2173,2175
no|2176,2178
central|2179,2186
pulmonary|2187,2196
embolism|2197,2205
.|2205,2206
<EOL>|2208,2209
The|2209,2212
thoracic|2213,2221
<EOL>|2222,2223
aorta|2223,2228
is|2229,2231
normal|2232,2238
in|2239,2241
caliber|2242,2249
without|2250,2257
evidence|2258,2266
of|2267,2269
dissection|2270,2280
or|2281,2283
<EOL>|2284,2285
intramural|2285,2295
<EOL>|2296,2297
hematoma|2297,2305
.|2305,2306
The|2308,2311
heart|2312,2317
,|2317,2318
pericardium|2319,2330
,|2330,2331
and|2332,2335
great|2336,2341
vessels|2342,2349
are|2350,2353
within|2354,2360
<EOL>|2361,2362
normal|2362,2368
limits|2369,2375
.|2375,2376
<EOL>|2377,2378
No|2378,2380
pericardial|2381,2392
effusion|2393,2401
is|2402,2404
seen|2405,2409
.|2409,2410
<EOL>|2411,2412
<EOL>|2414,2415
AXILLA|2415,2421
,|2421,2422
HILA|2423,2427
,|2427,2428
AND|2429,2432
MEDIASTINUM|2433,2444
:|2444,2445
There|2446,2451
is|2452,2454
a|2455,2456
8.8|2457,2460
x|2461,2462
5.8|2463,2466
x|2467,2468
9.8|2469,2472
cm|2473,2475
<EOL>|2476,2477
collection|2477,2487
in|2488,2490
the|2491,2494
<EOL>|2495,2496
left|2496,2500
breast|2501,2507
,|2507,2508
with|2509,2513
density|2514,2521
measuring|2522,2531
39|2532,2534
Hounsfield|2535,2545
units|2546,2551
,|2551,2552
<EOL>|2553,2554
consistent|2554,2564
with|2565,2569
<EOL>|2570,2571
hematoma|2571,2579
.|2579,2580
There|2582,2587
are|2588,2591
few|2592,2595
foci|2596,2600
of|2601,2603
air|2604,2607
within|2608,2614
the|2615,2618
collection|2619,2629
,|2629,2630
<EOL>|2631,2632
likely|2632,2638
from|2639,2643
prior|2644,2649
<EOL>|2650,2651
aspiration|2651,2661
,|2661,2662
as|2663,2665
well|2666,2670
as|2671,2673
few|2674,2677
punctate|2678,2686
hyperdensities|2687,2701
at|2702,2704
the|2705,2708
<EOL>|2709,2710
periphery|2710,2719
.|2719,2720
No|2722,2724
<EOL>|2725,2726
axillary|2726,2734
,|2734,2735
mediastinal|2736,2747
,|2747,2748
or|2749,2751
hilar|2752,2757
lymphadenopathy|2758,2773
is|2774,2776
present|2777,2784
.|2784,2785
The|2787,2790
<EOL>|2791,2792
right|2792,2797
axilla|2798,2804
<EOL>|2805,2806
is|2806,2808
not|2809,2812
included|2813,2821
on|2822,2824
the|2825,2828
study|2829,2834
.|2834,2835
No|2837,2839
mediastinal|2840,2851
mass|2852,2856
.|2856,2857
<EOL>|2858,2859
<EOL>|2861,2862
PLEURAL|2862,2869
SPACES|2870,2876
:|2876,2877
No|2878,2880
pleural|2881,2888
effusion|2889,2897
or|2898,2900
pneumothorax|2901,2913
.|2913,2914
<EOL>|2915,2916
<EOL>|2918,2919
LUNGS|2919,2924
/|2924,2925
AIRWAYS|2925,2932
:|2932,2933
Partially|2934,2943
visualized|2944,2954
lungs|2955,2960
are|2961,2964
clear|2965,2970
without|2971,2978
<EOL>|2979,2980
masses|2980,2986
or|2987,2989
areas|2990,2995
of|2996,2998
<EOL>|2999,3000
parenchymal|3000,3011
opacification|3012,3025
.|3025,3026
The|3028,3031
airways|3032,3039
are|3040,3043
patent|3044,3050
to|3051,3053
the|3054,3057
level|3058,3063
<EOL>|3064,3065
of|3065,3067
the|3068,3071
<EOL>|3072,3073
segmental|3073,3082
bronchi|3083,3090
bilaterally|3091,3102
.|3102,3103
<EOL>|3104,3105
<EOL>|3107,3108
BASE|3108,3112
OF|3113,3115
NECK|3116,3120
:|3120,3121
Visualized|3122,3132
portions|3133,3141
of|3142,3144
the|3145,3148
base|3149,3153
of|3154,3156
the|3157,3160
neck|3161,3165
show|3166,3170
<EOL>|3171,3172
no|3172,3174
abnormality|3175,3186
.|3186,3187
<EOL>|3188,3189
<EOL>|3191,3192
BONES|3192,3197
:|3197,3198
No|3199,3201
suspicious|3202,3212
osseous|3213,3220
abnormality|3221,3232
is|3233,3235
seen|3236,3240
.|3240,3241
?|3241,3242
There|3243,3248
is|3249,3251
no|3252,3254
<EOL>|3255,3256
acute|3256,3261
fracture|3262,3270
.|3270,3271
<EOL>|3272,3273
<EOL>|3275,3276
8.8|3293,3296
x|3297,3298
5.8|3299,3302
x|3303,3304
9.8|3305,3308
cm|3309,3311
left|3312,3316
breast|3317,3323
hematoma|3324,3332
,|3332,3333
with|3334,3338
no|3339,3341
evidence|3342,3350
of|3351,3353
<EOL>|3354,3355
active|3355,3361
bleed|3362,3367
.|3367,3368
<EOL>|3370,3371
Please|3371,3377
note|3378,3382
,|3382,3383
timing|3384,3390
was|3391,3394
suboptimal|3395,3405
as|3406,3408
the|3409,3412
patient|3413,3420
needed|3421,3427
to|3428,3430
be|3431,3433
<EOL>|3434,3435
re-scanned|3435,3445
due|3446,3449
<EOL>|3450,3451
to|3451,3453
incomplete|3454,3464
field|3465,3470
-|3470,3471
of|3471,3473
-|3473,3474
view|3474,3478
on|3479,3481
initial|3482,3489
images|3490,3496
,|3496,3497
however|3498,3505
,|3505,3506
the|3507,3510
<EOL>|3511,3512
density|3512,3519
of|3520,3522
the|3523,3526
<EOL>|3527,3528
collection|3528,3538
was|3539,3542
unchanged|3543,3552
on|3553,3555
all|3556,3559
series|3560,3566
.|3566,3567
<EOL>|3568,3569
<EOL>|3569,3570
<EOL>|3571,3572
Ms.|3595,3598
_|3599,3600
_|3600,3601
_|3601,3602
is|3603,3605
a|3606,3607
_|3608,3609
_|3609,3610
_|3610,3611
woman|3612,3617
who|3618,3621
was|3622,3625
admitted|3626,3634
to|3635,3637
the|3638,3641
<EOL>|3642,3643
breast|3643,3649
service|3650,3657
following|3658,3667
a|3668,3669
left|3670,3674
breast|3675,3681
lumpectomy|3682,3692
for|3693,3696
invasive|3697,3705
<EOL>|3706,3707
carcinoma|3707,3716
performed|3717,3726
on|3727,3729
_|3730,3731
_|3731,3732
_|3732,3733
.|3733,3734
She|3735,3738
presented|3739,3748
with|3749,3753
a|3754,3755
recurrent|3756,3765
<EOL>|3766,3767
left|3767,3771
breast|3772,3778
hematoma|3779,3787
after|3788,3793
it|3794,3796
was|3797,3800
evacuated|3801,3810
by|3811,3813
needle|3814,3820
aspiration|3821,3831
<EOL>|3832,3833
in|3833,3835
clinic|3836,3842
on|3843,3845
_|3846,3847
_|3847,3848
_|3848,3849
.|3849,3850
She|3851,3854
was|3855,3858
admitted|3859,3867
for|3868,3871
observation|3872,3883
and|3884,3887
<EOL>|3888,3889
surgical|3889,3897
evacuation|3898,3908
of|3909,3911
her|3912,3915
hematoma|3916,3924
.|3924,3925
<EOL>|3926,3927
<EOL>|3927,3928
On|3928,3930
_|3931,3932
_|3932,3933
_|3933,3934
she|3935,3938
was|3939,3942
brought|3943,3950
to|3951,3953
the|3954,3957
operating|3958,3967
room|3968,3972
for|3973,3976
evacuation|3977,3987
<EOL>|3988,3989
of|3989,3991
the|3992,3995
left|3996,4000
_|4001,4002
_|4002,4003
_|4003,4004
hematoma|4005,4013
and|4014,4017
placement|4018,4027
of|4028,4030
a|4031,4032
surgical|4033,4041
drain|4042,4047
.|4047,4048
<EOL>|4049,4050
Hospital|4050,4058
course|4059,4065
as|4066,4068
detailed|4069,4077
below|4078,4083
:|4083,4084
<EOL>|4084,4085
<EOL>|4085,4086
Neuro|4086,4091
:|4091,4092
pain|4093,4097
was|4098,4101
controlled|4102,4112
with|4113,4117
oral|4118,4122
pain|4123,4127
medication|4128,4138
including|4139,4148
<EOL>|4149,4150
acetaminophen|4150,4163
and|4164,4167
tramadol|4168,4176
.|4176,4177
<EOL>|4178,4179
<EOL>|4179,4180
_|4180,4181
_|4181,4182
_|4182,4183
:|4183,4184
Vital|4185,4190
signs|4191,4196
were|4197,4201
monitored|4202,4211
per|4212,4215
protocol|4216,4224
.|4224,4225
She|4226,4229
was|4230,4233
continued|4234,4243
<EOL>|4244,4245
on|4245,4247
her|4248,4251
home|4252,4256
medications|4257,4268
.|4268,4269
<EOL>|4270,4271
<EOL>|4271,4272
Resp|4272,4276
:|4276,4277
she|4278,4281
was|4282,4285
continued|4286,4295
on|4296,4298
her|4299,4302
home|4303,4307
albuterol|4308,4317
medications|4318,4329
<EOL>|4329,4330
<EOL>|4330,4331
FEN|4331,4334
/|4334,4335
GI|4335,4337
:|4337,4338
she|4339,4342
was|4343,4346
continued|4347,4356
on|4357,4359
a|4360,4361
regular|4362,4369
diet|4370,4374
throughout|4375,4385
her|4386,4389
<EOL>|4390,4391
admission|4391,4400
.|4400,4401
She|4402,4405
was|4406,4409
briefly|4410,4417
made|4418,4422
NPO|4423,4426
for|4427,4430
the|4431,4434
operating|4435,4444
room|4445,4449
and|4450,4453
<EOL>|4454,4455
hydrated|4455,4463
with|4464,4468
IV|4469,4471
fluids|4472,4478
in|4479,4481
the|4482,4485
perioperative|4486,4499
period|4500,4506
.|4506,4507
<EOL>|4508,4509
<EOL>|4509,4510
GU|4510,4512
:|4512,4513
She|4514,4517
voided|4518,4524
without|4525,4532
issue|4533,4538
throughout|4539,4549
her|4550,4553
hospital|4554,4562
course|4563,4569
<EOL>|4569,4570
<EOL>|4570,4571
Heme|4571,4575
:|4575,4576
H|4577,4578
/|4578,4579
H|4579,4580
was|4581,4584
closely|4585,4592
monitored|4593,4602
with|4603,4607
daily|4608,4613
labs|4614,4618
and|4619,4622
found|4623,4628
to|4629,4631
be|4632,4634
<EOL>|4635,4636
stable|4636,4642
.|4642,4643
Her|4644,4647
home|4648,4652
anticoagulation|4653,4668
was|4669,4672
held|4673,4677
during|4678,4684
her|4685,4688
hospital|4689,4697
<EOL>|4698,4699
course|4699,4705
.|4705,4706
She|4707,4710
was|4711,4714
resumed|4715,4722
on|4723,4725
her|4726,4729
home|4730,4734
dose|4735,4739
of|4740,4742
warfarin|4743,4751
on|4752,4754
<EOL>|4755,4756
discharge|4756,4765
without|4766,4773
a|4774,4775
lovenox|4776,4783
bridge|4784,4790
.|4790,4791
She|4792,4795
remained|4796,4804
on|4805,4807
compression|4808,4819
<EOL>|4820,4821
boots|4821,4826
during|4827,4833
her|4834,4837
hospital|4838,4846
course|4847,4853
to|4854,4856
prevent|4857,4864
DVTs|4865,4869
.|4869,4870
<EOL>|4870,4871
<EOL>|4871,4872
ID|4872,4874
:|4874,4875
She|4876,4879
was|4880,4883
given|4884,4889
ancef|4890,4895
2gm|4896,4899
IV|4900,4902
Q8hrs|4903,4908
for|4909,4912
prophylaxis|4913,4924
,|4924,4925
she|4926,4929
<EOL>|4930,4931
remained|4931,4939
afebrile|4940,4948
and|4949,4952
did|4953,4956
not|4957,4960
develop|4961,4968
a|4969,4970
leukocytosis|4971,4983
during|4984,4990
her|4991,4994
<EOL>|4995,4996
hospital|4996,5004
course|5005,5011
.|5011,5012
<EOL>|5013,5014
<EOL>|5014,5015
Endo|5015,5019
:|5019,5020
Due|5021,5024
to|5025,5027
a|5028,5029
history|5030,5037
of|5038,5040
metabolic|5041,5050
syndrome|5051,5059
and|5060,5063
pre-diabetes|5064,5076
<EOL>|5077,5078
she|5078,5081
was|5082,5085
kept|5086,5090
on|5091,5093
a|5094,5095
constant|5096,5104
carbohydrate|5105,5117
diet|5118,5122
.|5122,5123
<EOL>|5124,5125
<EOL>|5125,5126
On|5126,5128
the|5129,5132
day|5133,5136
of|5137,5139
discharge|5140,5149
she|5150,5153
was|5154,5157
tolerating|5158,5168
a|5169,5170
regular|5171,5178
diet|5179,5183
w|5184,5185
/|5185,5186
o|5186,5187
<EOL>|5188,5189
nausea|5189,5195
or|5196,5198
emesis|5199,5205
.|5205,5206
She|5207,5210
was|5211,5214
ambulating|5215,5225
independently|5226,5239
.|5239,5240
Her|5241,5244
pain|5245,5249
was|5250,5253
<EOL>|5254,5255
controlled|5255,5265
with|5266,5270
oral|5271,5275
pain|5276,5280
medications|5281,5292
.|5292,5293
She|5294,5297
was|5298,5301
afebrile|5302,5310
and|5311,5314
did|5315,5318
<EOL>|5319,5320
not|5320,5323
have|5324,5328
a|5329,5330
leukocytosis|5331,5343
,|5343,5344
all|5345,5348
antibiotics|5349,5360
were|5361,5365
discontinued|5366,5378
.|5378,5379
She|5380,5383
<EOL>|5384,5385
was|5385,5388
discharged|5389,5399
home|5400,5404
with|5405,5409
_|5410,5411
_|5411,5412
_|5412,5413
for|5414,5417
drain|5418,5423
management|5424,5434
and|5435,5438
close|5439,5444
<EOL>|5445,5446
follow|5446,5452
up|5453,5455
with|5456,5460
Dr.|5461,5464
_|5465,5466
_|5466,5467
_|5467,5468
in|5469,5471
clinic|5472,5478
for|5479,5482
drain|5483,5488
removal|5489,5496
.|5496,5497
She|5498,5501
<EOL>|5502,5503
will|5503,5507
also|5508,5512
follow|5513,5519
up|5520,5522
with|5523,5527
Dr.|5528,5531
_|5532,5533
_|5533,5534
_|5534,5535
in|5536,5538
clinic|5539,5545
in|5546,5548
early|5549,5554
_|5555,5556
_|5556,5557
_|5557,5558
<EOL>|5559,5560
for|5560,5563
routine|5564,5571
follow|5572,5578
up|5579,5581
.|5581,5582
<EOL>|5583,5584
<EOL>|5584,5585
<EOL>|5586,5587
Medications|5587,5598
on|5599,5601
Admission|5602,5611
:|5611,5612
<EOL>|5612,5613
Active|5613,5619
Medication|5620,5630
list|5631,5635
as|5636,5638
of|5639,5641
_|5642,5643
_|5643,5644
_|5644,5645
:|5645,5646
<EOL>|5646,5647
<EOL>|5648,5649
Medications|5649,5660
-|5661,5662
Prescription|5663,5675
<EOL>|5675,5676
ALBUTEROL|5676,5685
SULFATE|5686,5693
-|5694,5695
albuterol|5696,5705
sulfate|5706,5713
2.5|5714,5717
mg|5718,5720
/|5720,5721
3|5721,5722
mL|5723,5725
(|5726,5727
0.083|5727,5732
%|5733,5734
)|5734,5735
<EOL>|5735,5736
solution|5736,5744
for|5745,5748
nebulization|5749,5761
.|5761,5762
3|5763,5764
ml|5765,5767
inhalation|5768,5778
four|5779,5783
times|5784,5789
a|5790,5791
day|5792,5795
as|5796,5798
<EOL>|5798,5799
needed|5799,5805
for|5806,5809
cough|5810,5815
,|5815,5816
wheeze|5817,5823
<EOL>|5823,5824
ALBUTEROL|5824,5833
SULFATE|5834,5841
[|5842,5843
PROAIR|5843,5849
HFA|5850,5853
]|5853,5854
-|5855,5856
ProAir|5857,5863
HFA|5864,5867
90|5868,5870
mcg|5871,5874
/|5874,5875
actuation|5875,5884
<EOL>|5884,5885
aerosol|5885,5892
inhaler.|5893,5901
2|5902,5903
puffs|5904,5909
inhalation|5910,5920
q4|5921,5923
-|5923,5924
6|5924,5925
hours|5926,5931
as|5932,5934
needed|5935,5941
for|5942,5945
<EOL>|5945,5946
cough|5946,5951
/|5951,5952
wheeze|5952,5958
<EOL>|5958,5959
ATORVASTATIN|5959,5971
-|5972,5973
atorvastatin|5974,5986
40|5987,5989
mg|5990,5992
tablet.|5993,6000
1|6001,6002
(|6003,6004
One|6004,6007
)|6007,6008
tablet|6009,6015
(|6015,6016
s|6016,6017
)|6017,6018
by|6019,6021
<EOL>|6021,6022
mouth|6022,6027
at|6028,6030
bedtime|6031,6038
-|6039,6040
(|6042,6043
Prescribed|6043,6053
by|6054,6056
Other|6057,6062
Provider|6063,6071
;|6071,6072
Dose|6073,6077
<EOL>|6077,6078
adjustment|6078,6088
-|6089,6090
no|6091,6093
new|6094,6097
Rx|6098,6100
)|6100,6101
<EOL>|6101,6102
ENOXAPARIN|6102,6112
-|6113,6114
enoxaparin|6115,6125
100|6126,6129
mg|6130,6132
/|6132,6133
mL|6133,6135
subcutaneous|6136,6148
syringe|6149,6156
.|6156,6157
100|6158,6161
mg|6162,6164
<EOL>|6165,6166
SC|6166,6168
<EOL>|6168,6169
twice|6169,6174
daily|6175,6180
approximately|6181,6194
12|6195,6197
hours|6198,6203
apart|6204,6209
(|6210,6211
will|6211,6215
start|6216,6221
_|6222,6223
_|6223,6224
_|6224,6225
,|6225,6226
<EOL>|6226,6227
last|6227,6231
dose|6232,6236
_|6237,6238
_|6238,6239
_|6239,6240
AM|6241,6243
)|6243,6244
.|6244,6245
-|6246,6247
(|6249,6250
Prescribed|6250,6260
by|6261,6263
Other|6264,6269
Provider|6270,6278
;|6278,6279
Dose|6280,6284
<EOL>|6284,6285
adjustment|6285,6295
-|6296,6297
no|6298,6300
new|6301,6304
Rx|6305,6307
)|6307,6308
<EOL>|6308,6309
ERYTHROMYCIN|6309,6321
-|6322,6323
erythromycin|6324,6336
5|6337,6338
mg|6339,6341
/|6341,6342
gram|6342,6346
(|6347,6348
0.5|6348,6351
%|6352,6353
)|6353,6354
eye|6355,6358
ointment|6359,6367
.|6367,6368
<EOL>|6369,6370
Apply|6370,6375
<EOL>|6375,6376
_|6376,6377
_|6377,6378
_|6378,6379
inch|6380,6384
affected|6385,6393
eye|6394,6397
four|6398,6402
times|6403,6408
a|6409,6410
day|6411,6414
<EOL>|6414,6415
FUROSEMIDE|6415,6425
-|6426,6427
furosemide|6428,6438
20|6439,6441
mg|6442,6444
tablet|6445,6451
.|6451,6452
_|6453,6454
_|6454,6455
_|6455,6456
tablet|6457,6463
(|6463,6464
s|6464,6465
)|6465,6466
by|6467,6469
mouth|6470,6475
<EOL>|6475,6476
once|6476,6480
a|6481,6482
day|6483,6486
as|6487,6489
needed|6490,6496
for|6497,6500
leg|6501,6504
swelling|6505,6513
<EOL>|6513,6514
HYDROMORPHONE|6514,6527
-|6528,6529
hydromorphone|6530,6543
2|6544,6545
mg|6546,6548
tablet|6549,6555
.|6555,6556
_|6557,6558
_|6558,6559
_|6559,6560
tablet|6561,6567
(|6567,6568
s|6568,6569
)|6569,6570
by|6571,6573
<EOL>|6573,6574
mouth|6574,6579
every|6580,6585
four|6586,6590
(|6591,6592
4|6592,6593
)|6593,6594
hours|6595,6600
as|6601,6603
needed|6604,6610
for|6611,6614
severe|6615,6621
pain|6622,6626
do|6627,6629
not|6630,6633
<EOL>|6634,6635
drink|6635,6640
<EOL>|6640,6641
alcohol|6641,6648
or|6649,6651
drive|6652,6657
while|6658,6663
taking|6664,6670
this|6671,6675
medication|6676,6686
<EOL>|6686,6687
NEBULIZER|6687,6696
AND|6697,6700
COMPRESSOR|6701,6711
[|6712,6713
PORTABLE|6713,6721
NEBULIZER|6722,6731
SYSTEM|6732,6738
]|6738,6739
-|6740,6741
Portable|6742,6750
<EOL>|6750,6751
Nebulizer|6751,6760
System|6761,6767
.|6767,6768
Use|6769,6772
with|6773,6777
albuterol|6778,6787
nebulizer|6788,6797
soln|6798,6802
four|6803,6807
times|6808,6813
a|6814,6815
<EOL>|6815,6816
day|6816,6819
as|6820,6822
needed|6823,6829
for|6830,6833
cough|6834,6839
/|6839,6840
wheeze|6840,6846
<EOL>|6846,6847
OMEPRAZOLE|6847,6857
-|6858,6859
omeprazole|6860,6870
20|6871,6873
mg|6874,6876
capsule|6877,6884
,|6884,6885
delayed|6885,6892
release|6893,6900
.|6900,6901
TAKE|6902,6906
1|6907,6908
<EOL>|6908,6909
CAPSULE|6909,6916
TWICE|6917,6922
DAILY|6923,6928
FOR|6929,6932
GASTROESOPHAGEAL|6933,6949
REFLUXDISEASE|6950,6963
<EOL>|6963,6964
SERTRALINE|6964,6974
-|6975,6976
sertraline|6977,6987
100|6988,6991
mg|6992,6994
tablet|6995,7001
.|7001,7002
1.5|7003,7006
tablet|7007,7013
(|7013,7014
s|7014,7015
)|7015,7016
by|7017,7019
mouth|7020,7025
<EOL>|7025,7026
once|7026,7030
a|7031,7032
day|7033,7036
<EOL>|7036,7037
TRAMADOL|7037,7045
-|7046,7047
tramadol|7048,7056
50|7057,7059
mg|7060,7062
tablet.|7063,7070
one|7071,7074
tablet|7075,7081
(|7081,7082
s|7082,7083
)|7083,7084
by|7085,7087
mouth|7088,7093
three|7094,7099
<EOL>|7099,7100
times|7100,7105
a|7106,7107
day|7108,7111
<EOL>|7111,7112
TRAZODONE|7112,7121
-|7122,7123
trazodone|7124,7133
50|7134,7136
mg|7137,7139
tablet.|7140,7147
1|7148,7149
tablet|7150,7156
(|7156,7157
s|7157,7158
)|7158,7159
by|7160,7162
mouth|7163,7168
at|7169,7171
<EOL>|7171,7172
bedtime|7172,7179
as|7180,7182
needed|7183,7189
for|7190,7193
insomia|7194,7201
<EOL>|7201,7202
WARFARIN|7202,7210
-|7211,7212
warfarin|7213,7221
5|7222,7223
mg|7224,7226
tablet.|7227,7234
1|7235,7236
(|7237,7238
One|7238,7241
)|7241,7242
tablet|7243,7249
(|7249,7250
s|7250,7251
)|7251,7252
by|7253,7255
mouth|7256,7261
2|7262,7263
<EOL>|7263,7264
times|7264,7269
a|7270,7271
_|7272,7273
_|7273,7274
_|7274,7275
,|7275,7276
_|7277,7278
_|7278,7279
_|7279,7280
tabs|7281,7285
po|7286,7288
5|7289,7290
times|7291,7296
a|7297,7298
week|7299,7303
(|7304,7305
last|7305,7309
dose|7310,7314
per|7315,7318
<EOL>|7318,7319
_|7319,7320
_|7320,7321
_|7321,7322
clinic|7323,7329
_|7330,7331
_|7331,7332
_|7332,7333
-|7334,7335
(|7337,7338
Prescribed|7338,7348
by|7349,7351
Other|7352,7357
Provider|7358,7366
;|7366,7367
Dose|7368,7372
<EOL>|7372,7373
adjustment|7373,7383
-|7384,7385
no|7386,7388
new|7389,7392
Rx|7393,7395
)|7395,7396
<EOL>|7396,7397
<EOL>|7398,7399
Medications|7399,7410
-|7411,7412
OTC|7413,7416
<EOL>|7416,7417
ACETAMINOPHEN|7417,7430
-|7431,7432
acetaminophen|7433,7446
500|7447,7450
mg|7451,7453
tablet.|7454,7461
2|7462,7463
tablet|7464,7470
(|7470,7471
s|7471,7472
)|7472,7473
by|7474,7476
<EOL>|7477,7478
mouth|7478,7483
<EOL>|7483,7484
3|7484,7485
times|7486,7491
daily|7492,7497
as|7498,7500
needed|7501,7507
for|7508,7511
pain|7512,7516
-|7517,7518
_|7520,7521
_|7521,7522
_|7522,7523
DC|7524,7526
med|7527,7530
rec|7531,7534
)|7534,7535
<EOL>|7535,7536
CHOLECALCIFEROL|7536,7551
(|7552,7553
VITAMIN|7553,7560
D3|7561,7563
)|7563,7564
-|7565,7566
cholecalciferol|7567,7582
(|7583,7584
vitamin|7584,7591
D3|7592,7594
)|7594,7595
<EOL>|7596,7597
2,000|7597,7602
<EOL>|7602,7603
unit|7603,7607
tablet.|7608,7615
1|7616,7617
tablet|7618,7624
(|7624,7625
s|7625,7626
)|7626,7627
by|7628,7630
mouth|7631,7636
once|7637,7641
a|7642,7643
day|7644,7647
-|7648,7649
(|7651,7652
OTC|7652,7655
)|7655,7656
<EOL>|7656,7657
POLYETHYLENE|7657,7669
GLYCOL|7670,7676
3350|7677,7681
[|7682,7683
MIRALAX|7683,7690
]|7690,7691
-|7692,7693
Miralax|7694,7701
17|7702,7704
gram|7705,7709
/|7709,7710
dose|7710,7714
oral|7715,7719
<EOL>|7719,7720
powder.|7720,7727
1|7728,7729
powder|7730,7736
(|7736,7737
s|7737,7738
)|7738,7739
by|7740,7742
mouth|7743,7748
once|7749,7753
a|7754,7755
day|7756,7759
as|7760,7762
needed|7763,7769
for|7770,7773
<EOL>|7773,7774
constipation|7774,7786
-|7787,7788
(|7790,7791
Prescribed|7791,7801
by|7802,7804
Other|7805,7810
Provider|7811,7819
;|7819,7820
Dose|7821,7825
adjustment|7826,7836
-|7837,7838
<EOL>|7838,7839
no|7839,7841
new|7842,7845
Rx|7846,7848
)|7848,7849
<EOL>|7849,7850
SENNOSIDES|7850,7860
[|7861,7862
SENNA|7862,7867
]|7867,7868
-|7869,7870
senna|7871,7876
8.6|7877,7880
mg|7881,7883
tablet.|7884,7891
1|7892,7893
tablet|7894,7900
(|7900,7901
s|7901,7902
)|7902,7903
by|7904,7906
mouth|7907,7912
<EOL>|7912,7913
once|7913,7917
a|7918,7919
day|7920,7923
as|7924,7926
needed|7927,7933
for|7934,7937
constipation|7938,7950
-|7951,7952
(|7954,7955
OTC|7955,7958
)|7958,7959
<EOL>|7959,7960
<EOL>|7960,7961
<EOL>|7962,7963
Discharge|7963,7972
Medications|7973,7984
:|7984,7985
<EOL>|7985,7986
1.|7986,7988
TraMADol|7990,7998
50|7999,8001
mg|8002,8004
PO|8005,8007
Q4H|8008,8011
:|8011,8012
PRN|8012,8015
Pain|8016,8020
-|8021,8022
Moderate|8023,8031
<EOL>|8032,8033
Reason|8035,8041
for|8042,8045
PRN|8046,8049
duplicate|8050,8059
override|8060,8068
:|8068,8069
Alternating|8070,8081
agents|8082,8088
for|8089,8092
<EOL>|8093,8094
similar|8094,8101
severity|8102,8110
<EOL>|8110,8111
RX|8111,8113
*|8114,8115
tramadol|8115,8123
50|8124,8126
mg|8127,8129
1|8130,8131
tablet|8132,8138
(|8138,8139
s|8139,8140
)|8140,8141
by|8142,8144
mouth|8145,8150
Q4hr|8151,8155
prn|8156,8159
Disp|8160,8164
#|8165,8166
*|8166,8167
7|8167,8168
Tablet|8169,8175
<EOL>|8176,8177
Refills|8177,8184
:|8184,8185
*|8185,8186
0|8186,8187
<EOL>|8188,8189
2.|8189,8191
Atorvastatin|8193,8205
40|8206,8208
mg|8209,8211
PO|8212,8214
QPM|8215,8218
<EOL>|8220,8221
3.|8221,8223
Docusate|8225,8233
Sodium|8234,8240
100|8241,8244
mg|8245,8247
PO|8248,8250
BID|8251,8254
<EOL>|8256,8257
4.|8257,8259
Omeprazole|8261,8271
20|8272,8274
mg|8275,8277
PO|8278,8280
BID|8281,8284
<EOL>|8286,8287
5.|8287,8289
Senna|8291,8296
17.2|8297,8301
mg|8302,8304
PO|8305,8307
HS|8308,8310
<EOL>|8312,8313
6.|8313,8315
Sertraline|8317,8327
150|8328,8331
mg|8332,8334
PO|8335,8337
DAILY|8338,8343
<EOL>|8345,8346
7.|8346,8348
TraZODone|8350,8359
50|8360,8362
mg|8363,8365
PO|8366,8368
QHS|8369,8372
:|8372,8373
PRN|8373,8376
sleep|8377,8382
<EOL>|8384,8385
<EOL>|8385,8386
<EOL>|8387,8388
Discharge|8388,8397
Disposition|8398,8409
:|8409,8410
<EOL>|8410,8411
Home|8411,8415
With|8416,8420
Service|8421,8428
<EOL>|8428,8429
<EOL>|8430,8431
Facility|8431,8439
:|8439,8440
<EOL>|8440,8441
_|8441,8442
_|8442,8443
_|8443,8444
<EOL>|8444,8445
<EOL>|8446,8447
Discharge|8447,8456
Diagnosis|8457,8466
:|8466,8467
<EOL>|8467,8468
breast|8468,8474
hematoma|8475,8483
<EOL>|8484,8485
<EOL>|8485,8486
<EOL>|8487,8488
Mental|8509,8515
Status|8516,8522
:|8522,8523
Clear|8524,8529
and|8530,8533
coherent|8534,8542
.|8542,8543
<EOL>|8543,8544
Level|8544,8549
of|8550,8552
Consciousness|8553,8566
:|8566,8567
Alert|8568,8573
and|8574,8577
interactive|8578,8589
.|8589,8590
<EOL>|8590,8591
Activity|8591,8599
Status|8600,8606
:|8606,8607
Ambulatory|8608,8618
-|8619,8620
Independent|8621,8632
.|8632,8633
<EOL>|8633,8634
<EOL>|8634,8635
<EOL>|8636,8637
Personal|8661,8669
Care|8670,8674
:|8674,8675
<EOL>|8677,8678
1|8678,8679
.|8679,8680
You|8681,8684
may|8685,8688
keep|8689,8693
your|8694,8698
incisions|8699,8708
open|8709,8713
to|8714,8716
air|8717,8720
or|8721,8723
covered|8724,8731
with|8732,8736
a|8737,8738
<EOL>|8739,8740
clean|8740,8745
,|8745,8746
sterile|8747,8754
gauze|8755,8760
that|8761,8765
you|8766,8769
change|8770,8776
daily|8777,8782
.|8782,8783
<EOL>|8783,8784
2.|8784,8786
Clean|8787,8792
around|8793,8799
the|8800,8803
drain|8804,8809
site|8810,8814
(|8814,8815
s|8815,8816
)|8816,8817
,|8817,8818
where|8819,8824
the|8825,8828
tubing|8829,8835
exits|8836,8841
the|8842,8845
<EOL>|8846,8847
skin|8847,8851
,|8851,8852
with|8853,8857
soap|8858,8862
and|8863,8866
water|8867,8872
.|8872,8873
<EOL>|8875,8876
3.|8876,8878
Strip|8879,8884
drain|8885,8890
tubing|8891,8897
,|8897,8898
empty|8899,8904
bulb|8905,8909
(|8909,8910
s|8910,8911
)|8911,8912
,|8912,8913
and|8914,8917
record|8918,8924
output|8925,8931
(|8931,8932
s|8932,8933
)|8933,8934
_|8935,8936
_|8936,8937
_|8937,8938
<EOL>|8939,8940
times|8940,8945
per|8946,8949
day|8950,8953
.|8953,8954
<EOL>|8956,8957
4.|8957,8959
A|8960,8961
written|8962,8969
record|8970,8976
of|8977,8979
the|8980,8983
daily|8984,8989
output|8990,8996
from|8997,9001
each|9002,9006
drain|9007,9012
should|9013,9019
<EOL>|9020,9021
be|9021,9023
brought|9024,9031
to|9032,9034
every|9035,9040
follow|9041,9047
-|9047,9048
up|9048,9050
appointment|9051,9062
.|9062,9063
Your|9064,9068
drains|9069,9075
will|9076,9080
be|9081,9083
<EOL>|9084,9085
removed|9085,9092
as|9093,9095
soon|9096,9100
as|9101,9103
possible|9104,9112
when|9113,9117
the|9118,9121
daily|9122,9127
output|9128,9134
tapers|9135,9141
off|9142,9145
to|9146,9148
<EOL>|9149,9150
an|9150,9152
acceptable|9153,9163
amount|9164,9170
.|9170,9171
<EOL>|9173,9174
5|9174,9175
.|9175,9176
You|9177,9180
may|9181,9184
wear|9185,9189
a|9190,9191
surgical|9192,9200
bra|9201,9204
or|9205,9207
soft|9208,9212
,|9212,9213
loose|9214,9219
camisole|9220,9228
for|9229,9232
<EOL>|9233,9234
comfort|9234,9241
.|9241,9242
<EOL>|9244,9245
6.|9245,9247
Do|9248,9250
not|9251,9254
shower|9255,9261
while|9262,9267
your|9268,9272
drain|9273,9278
is|9279,9281
in|9282,9284
place|9285,9290
.|9290,9291
<EOL>|9292,9293
7.|9293,9295
The|9296,9299
Dermabond|9300,9309
skin|9310,9314
glue|9315,9319
will|9320,9324
begin|9325,9330
to|9331,9333
flake|9334,9339
off|9340,9343
in|9344,9346
about|9347,9352
_|9353,9354
_|9354,9355
_|9355,9356
<EOL>|9357,9358
days|9358,9362
.|9362,9363
<EOL>|9365,9366
<EOL>|9366,9367
Activity|9367,9375
:|9375,9376
<EOL>|9378,9379
1|9379,9380
.|9380,9381
You|9382,9385
may|9386,9389
resume|9390,9396
your|9397,9401
regular|9402,9409
diet|9410,9414
.|9414,9415
<EOL>|9417,9418
2.|9418,9420
Walk|9421,9425
several|9426,9433
times|9434,9439
a|9440,9441
day|9442,9445
.|9445,9446
<EOL>|9448,9449
3.|9449,9451
DO|9452,9454
NOT|9455,9458
lift|9459,9463
anything|9464,9472
heavier|9473,9480
than|9481,9485
5|9486,9487
pounds|9488,9494
or|9495,9497
engage|9498,9504
in|9505,9507
<EOL>|9508,9509
strenuous|9509,9518
activity|9519,9527
for|9528,9531
6|9532,9533
weeks|9534,9539
following|9540,9549
surgery|9550,9557
.|9557,9558
<EOL>|9559,9560
<EOL>|9560,9561
1.|9576,9578
Resume|9579,9585
your|9586,9590
regular|9591,9598
medications|9599,9610
unless|9611,9617
instructed|9618,9628
otherwise|9629,9638
<EOL>|9639,9640
and|9640,9643
take|9644,9648
any|9649,9652
new|9653,9656
meds|9657,9661
as|9662,9664
ordered|9665,9672
.|9673,9674
<EOL>|9676,9677
2|9677,9678
.|9678,9679
You|9680,9683
may|9684,9687
take|9688,9692
your|9693,9697
prescribed|9698,9708
pain|9709,9713
medication|9714,9724
for|9725,9728
moderate|9729,9737
to|9738,9740
<EOL>|9741,9742
severe|9742,9748
pain|9749,9753
.|9753,9754
You|9755,9758
may|9759,9762
switch|9763,9769
to|9770,9772
Tylenol|9773,9780
or|9781,9783
Extra|9784,9789
Strength|9790,9798
Tylenol|9799,9806
<EOL>|9807,9808
for|9808,9811
mild|9812,9816
pain|9817,9821
as|9822,9824
directed|9825,9833
on|9834,9836
the|9837,9840
packaging|9841,9850
.|9850,9851
Please|9852,9858
note|9859,9863
that|9864,9868
<EOL>|9869,9870
Percocet|9870,9878
and|9879,9882
Vicodin|9883,9890
have|9891,9895
Tylenol|9896,9903
as|9904,9906
an|9907,9909
active|9910,9916
ingredient|9917,9927
so|9928,9930
do|9931,9933
<EOL>|9934,9935
not|9935,9938
take|9939,9943
these|9944,9949
meds|9950,9954
with|9955,9959
additional|9960,9970
Tylenol|9971,9978
.|9978,9979
<EOL>|9981,9982
3.|9982,9984
Take|9985,9989
prescription|9990,10002
pain|10003,10007
medications|10008,10019
for|10020,10023
pain|10024,10028
not|10029,10032
relieved|10033,10041
by|10042,10044
<EOL>|10045,10046
Tylenol|10046,10053
.|10053,10054
<EOL>|10056,10057
4.|10057,10059
Take|10060,10064
Colace|10065,10071
,|10071,10072
100|10073,10076
mg|10077,10079
by|10080,10082
mouth|10083,10088
2|10089,10090
times|10091,10096
per|10097,10100
day|10101,10104
,|10104,10105
while|10106,10111
taking|10112,10118
<EOL>|10119,10120
the|10120,10123
prescription|10124,10136
pain|10137,10141
medication|10142,10152
.|10152,10153
You|10154,10157
may|10158,10161
use|10162,10165
a|10166,10167
different|10168,10177
<EOL>|10178,10179
over-the|10179,10187
-|10187,10188
counter|10188,10195
stool|10196,10201
softener|10202,10210
if|10211,10213
you|10214,10217
wish|10218,10222
.|10222,10223
<EOL>|10225,10226
5.|10226,10228
Do|10229,10231
not|10232,10235
drive|10236,10241
or|10242,10244
operate|10245,10252
heavy|10253,10258
machinery|10259,10268
while|10269,10274
taking|10275,10281
any|10282,10285
<EOL>|10286,10287
narcotic|10287,10295
pain|10296,10300
medication|10301,10311
.|10311,10312
You|10313,10316
may|10317,10320
have|10321,10325
constipation|10326,10338
when|10339,10343
taking|10344,10350
<EOL>|10351,10352
narcotic|10352,10360
pain|10361,10365
medications|10366,10377
(|10378,10379
oxycodone|10379,10388
,|10388,10389
percocet|10390,10398
,|10398,10399
vicodin|10400,10407
,|10407,10408
<EOL>|10409,10410
hydrocodone|10410,10421
,|10421,10422
dilaudid|10423,10431
,|10431,10432
etc|10433,10436
.|10436,10437
)|10437,10438
;|10438,10439
you|10440,10443
should|10444,10450
continue|10451,10459
drinking|10460,10468
<EOL>|10469,10470
fluids|10470,10476
,|10476,10477
you|10478,10481
may|10482,10485
take|10486,10490
stool|10491,10496
softeners|10497,10506
,|10506,10507
and|10508,10511
should|10512,10518
eat|10519,10522
foods|10523,10528
that|10529,10533
<EOL>|10534,10535
are|10535,10538
high|10539,10543
in|10544,10546
fiber|10547,10552
.|10552,10553
<EOL>|10555,10556
<EOL>|10556,10557
Call|10557,10561
the|10562,10565
office|10566,10572
IMMEDIATELY|10573,10584
if|10585,10587
you|10588,10591
have|10592,10596
any|10597,10600
of|10601,10603
the|10604,10607
following|10608,10617
:|10617,10618
<EOL>|10620,10621
1.|10621,10623
Signs|10624,10629
of|10630,10632
infection|10633,10642
:|10642,10643
fever|10644,10649
with|10650,10654
chills|10655,10661
,|10661,10662
increased|10663,10672
redness|10673,10680
,|10680,10681
<EOL>|10682,10683
swelling|10683,10691
,|10691,10692
warmth|10693,10699
or|10700,10702
tenderness|10703,10713
at|10714,10716
the|10717,10720
surgical|10721,10729
site|10730,10734
,|10734,10735
or|10736,10738
unusual|10739,10746
<EOL>|10747,10748
drainage|10748,10756
from|10757,10761
the|10762,10765
incision|10766,10774
(|10774,10775
s|10775,10776
)|10776,10777
.|10777,10778
<EOL>|10780,10781
2|10781,10782
.|10782,10783
A|10784,10785
large|10786,10791
amount|10792,10798
of|10799,10801
bleeding|10802,10810
from|10811,10815
the|10816,10819
incision|10820,10828
(|10828,10829
s|10829,10830
)|10830,10831
or|10832,10834
drain|10835,10840
(|10840,10841
s|10841,10842
)|10842,10843
.|10843,10844
<EOL>|10846,10847
<EOL>|10847,10848
3.|10848,10850
Fever|10851,10856
greater|10857,10864
than|10865,10869
101.5|10870,10875
oF|10876,10878
<EOL>|10880,10881
4.|10881,10883
Severe|10884,10890
pain|10891,10895
NOT|10896,10899
relieved|10900,10908
by|10909,10911
your|10912,10916
medication|10917,10927
.|10927,10928
<EOL>|10930,10931
<EOL>|10933,10934
Return|10934,10940
to|10941,10943
the|10944,10947
ER|10948,10950
if|10951,10953
:|10953,10954
<EOL>|10956,10957
*|10957,10958
If|10959,10961
you|10962,10965
are|10966,10969
vomiting|10970,10978
and|10979,10982
can|10983,10986
not|10986,10989
keep|10990,10994
in|10995,10997
fluids|10998,11004
or|11005,11007
your|11008,11012
<EOL>|11013,11014
medications|11014,11025
.|11025,11026
<EOL>|11028,11029
*|11029,11030
If|11031,11033
you|11034,11037
have|11038,11042
shaking|11043,11050
chills|11051,11057
,|11057,11058
fever|11059,11064
greater|11065,11072
than|11073,11077
101.5|11078,11083
(|11084,11085
F|11085,11086
)|11086,11087
<EOL>|11088,11089
degrees|11089,11096
or|11097,11099
38|11100,11102
(|11103,11104
C|11104,11105
)|11105,11106
degrees|11107,11114
,|11114,11115
increased|11116,11125
redness|11126,11133
,|11133,11134
swelling|11135,11143
or|11144,11146
<EOL>|11147,11148
discharge|11148,11157
from|11158,11162
incision|11163,11171
,|11171,11172
chest|11173,11178
pain|11179,11183
,|11183,11184
shortness|11185,11194
of|11195,11197
breath|11198,11204
,|11204,11205
or|11206,11208
<EOL>|11209,11210
anything|11210,11218
else|11219,11223
that|11224,11228
is|11229,11231
troubling|11232,11241
you|11242,11245
.|11245,11246
<EOL>|11248,11249
*|11249,11250
Any|11251,11254
serious|11255,11262
change|11263,11269
in|11270,11272
your|11273,11277
symptoms|11278,11286
,|11286,11287
or|11288,11290
any|11291,11294
new|11295,11298
symptoms|11299,11307
that|11308,11312
<EOL>|11313,11314
concern|11314,11321
you|11322,11325
.|11325,11326
<EOL>|11328,11329
<EOL>|11329,11330
ANTICOAGULATION|11330,11345
:|11345,11346
<EOL>|11346,11347
You|11347,11350
should|11351,11357
begin|11358,11363
taking|11364,11370
your|11371,11375
home|11376,11380
warfarin|11381,11389
dose|11390,11394
this|11395,11399
evening|11400,11407
<EOL>|11408,11409
(|11409,11410
_|11410,11411
_|11411,11412
_|11412,11413
)|11413,11414
and|11415,11418
resume|11419,11425
taking|11426,11432
warfarin|11433,11441
at|11442,11444
your|11445,11449
regular|11450,11457
scheduled|11458,11467
<EOL>|11468,11469
doses|11469,11474
.|11474,11475
You|11476,11479
will|11480,11484
not|11485,11488
need|11489,11493
a|11494,11495
bridge|11496,11502
therapy|11503,11510
to|11511,11513
begin|11514,11519
warfarin|11520,11528
.|11528,11529
<EOL>|11530,11531
<EOL>|11531,11532
DRAIN|11532,11537
DISCHARGE|11538,11547
INSTRUCTIONS|11548,11560
<EOL>|11562,11563
You|11563,11566
are|11567,11570
being|11571,11576
discharged|11577,11587
with|11588,11592
drains|11593,11599
in|11600,11602
place|11603,11608
.|11608,11609
Drain|11610,11615
care|11616,11620
is|11621,11623
a|11624,11625
<EOL>|11626,11627
clean|11627,11632
procedure|11633,11642
.|11642,11643
Wash|11644,11648
your|11649,11653
hands|11654,11659
thoroughly|11660,11670
with|11671,11675
soap|11676,11680
and|11681,11684
warm|11685,11689
<EOL>|11690,11691
water|11691,11696
before|11697,11703
performing|11704,11714
drain|11715,11720
care|11721,11725
.|11725,11726
Perform|11727,11734
drainage|11735,11743
care|11744,11748
twice|11749,11754
<EOL>|11755,11756
a|11756,11757
day|11758,11761
.|11761,11762
Try|11763,11766
to|11767,11769
empty|11770,11775
the|11776,11779
drain|11780,11785
at|11786,11788
the|11789,11792
same|11793,11797
time|11798,11802
each|11803,11807
day|11808,11811
.|11811,11812
Pull|11813,11817
<EOL>|11818,11819
the|11819,11822
stopper|11823,11830
out|11831,11834
of|11835,11837
the|11838,11841
drainage|11842,11850
bottle|11851,11857
and|11858,11861
empty|11862,11867
the|11868,11871
drainage|11872,11880
<EOL>|11881,11882
fluid|11882,11887
into|11888,11892
the|11893,11896
measuring|11897,11906
cup|11907,11910
.|11910,11911
Record|11912,11918
the|11919,11922
amount|11923,11929
of|11930,11932
drainage|11933,11941
<EOL>|11942,11943
fluid|11943,11948
on|11949,11951
the|11952,11955
record|11956,11962
sheet|11963,11968
.|11968,11969
Reestablish|11970,11981
drain|11982,11987
suction|11988,11995
.|11995,11996
<EOL>|11998,11999
Please|11999,12005
assist|12006,12012
patient|12013,12020
with|12021,12025
drain|12026,12031
care|12032,12036
.|12036,12037
A|12038,12039
daily|12040,12045
log|12046,12049
of|12050,12052
individual|12053,12063
<EOL>|12064,12065
drain|12065,12070
outputs|12071,12078
should|12079,12085
be|12086,12088
maintained|12089,12099
and|12100,12103
brought|12104,12111
with|12112,12116
patient|12117,12124
to|12125,12127
<EOL>|12128,12129
follow|12129,12135
up|12136,12138
appointment|12139,12150
with|12151,12155
your|12156,12160
surgeon|12161,12168
.|12168,12169
<EOL>|12169,12170
<EOL>|12170,12171
<EOL>|12172,12173
Followup|12173,12181
Instructions|12182,12194
:|12194,12195
<EOL>|12195,12196
_|12196,12197
_|12197,12198
_|12198,12199
<EOL>|12199,12200

