 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
NEUROSURGERY|156,168
<EOL>|168,169
<EOL>|170,171
Penicillins|183,194
/|195,196
Paxil|197,202
/|203,204
Wellbutrin|205,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
Exposed|253,260
hardware|261,269
<EOL>|269,270
<EOL>|271,272
Major|272,277
Surgical|278,286
or|287,289
Invasive|290,298
Procedure|299,308
:|308,309
<EOL>|309,310
Exposed|310,317
hardware|318,326
removal|327,334
<EOL>|335,336
<EOL>|336,337
<EOL>|338,339
The|367,370
is|371,373
a|374,375
_|376,377
_|377,378
_|378,379
year|380,384
old|385,388
female|389,395
who|396,399
had|400,403
prior|404,409
surgery|410,417
for|418,421
a|422,423
possible|424,432
<EOL>|433,434
right|434,439
parietal|440,448
<EOL>|448,449
anaplastic|449,459
astrocytoma|460,471
with|472,476
craniotomy|477,487
for|488,491
resection|492,501
on|502,504
_|505,506
_|506,507
_|507,508
<EOL>|509,510
by|510,512
Dr.|513,516
_|517,518
_|518,519
_|519,520
in|521,523
_|524,525
_|525,526
_|526,527
followed|528,536
by|537,539
involved|540,548
-|548,549
field|549,554
<EOL>|555,556
irradiation|556,567
to|568,570
6,120|571,576
cGy|577,580
_|581,582
_|582,583
_|583,584
in|585,587
_|588,589
_|589,590
_|590,591
,|591,592
3|593,594
cycles|595,601
of|602,604
<EOL>|605,606
Temodar|606,613
ended|614,619
_|620,621
_|621,622
_|622,623
and|624,627
a|628,629
second|630,636
craniotomy|637,647
for|648,651
tumor|652,657
recurrence|658,668
<EOL>|669,670
on|670,672
_|673,674
_|674,675
_|675,676
by|677,679
Dr.|680,683
_|684,685
_|685,686
_|686,687
at|688,690
_|691,692
_|692,693
_|693,694
with|695,699
PCV|700,703
(|703,704
comb|704,708
chemo|709,714
)|714,715
_|716,717
_|717,718
_|718,719
-|720,721
<EOL>|721,722
_|722,723
_|723,724
_|724,725
.|725,726
<EOL>|728,729
<EOL>|729,730
In|730,732
_|733,734
_|734,735
_|735,736
she|737,740
presented|741,750
with|751,755
exposed|756,763
hardware|764,772
to|773,775
the|776,779
office|780,786
and|787,790
<EOL>|791,792
she|792,795
needed|796,802
admission|803,812
an|813,815
complex|816,823
revision|824,832
for|833,836
a|837,838
plate|839,844
that|845,849
had|850,853
<EOL>|854,855
eroded|855,861
through|862,869
the|870,873
skin|874,878
;|878,879
Plastics|880,888
and|889,892
I|893,894
reconstructed|895,908
the|909,912
scalp|913,918
<EOL>|919,920
at|920,922
that|923,927
time|928,932
.|932,933
<EOL>|933,934
<EOL>|934,935
The|935,938
patient|939,946
presents|947,955
today|956,961
again|962,967
with|968,972
some|973,977
history|978,985
of|986,988
pruritus|989,997
<EOL>|998,999
on|999,1001
the|1002,1005
top|1006,1009
of|1010,1012
her|1013,1016
head|1017,1021
and|1022,1025
newly|1026,1031
diagnosed|1032,1041
exposed|1042,1049
hardware|1050,1058
.|1058,1059
She|1060,1063
<EOL>|1064,1065
reports|1065,1072
that|1073,1077
she|1078,1081
had|1082,1085
her|1086,1089
husband|1090,1097
look|1098,1102
at|1103,1105
the|1106,1109
top|1110,1113
of|1114,1116
her|1117,1120
head|1121,1125
"|1126,1127
a|1128,1129
<EOL>|1130,1131
few|1131,1134
ago|1135,1138
"|1138,1139
and|1140,1143
saw|1144,1147
that|1148,1152
metal|1153,1158
hardware|1159,1167
from|1168,1172
her|1173,1176
prior|1177,1182
surgery|1183,1190
was|1191,1194
<EOL>|1195,1196
present|1196,1203
.|1203,1204
<EOL>|1204,1205
<EOL>|1206,1207
right|1229,1234
parietal|1235,1243
anaplastic|1244,1254
astrocytoma|1255,1266
,|1266,1267
Craniotomy|1268,1278
_|1279,1280
_|1280,1281
_|1281,1282
by|1283,1285
<EOL>|1287,1288
Dr.|1288,1291
_|1292,1293
_|1293,1294
_|1294,1295
in|1296,1298
_|1299,1300
_|1300,1301
_|1301,1302
irradiation|1303,1314
to|1315,1317
6,120|1318,1323
<EOL>|1324,1325
<EOL>|1326,1327
cGy|1327,1330
_|1331,1332
_|1332,1333
_|1333,1334
in|1335,1337
_|1338,1339
_|1339,1340
_|1340,1341
,|1341,1342
3|1342,1343
cycles|1344,1350
of|1351,1353
Temodar|1354,1361
ended|1362,1367
_|1368,1369
_|1369,1370
_|1370,1371
<EOL>|1373,1374
craniotomy|1374,1384
on|1385,1387
_|1388,1389
_|1389,1390
_|1390,1391
by|1392,1394
Dr.|1395,1398
_|1399,1400
_|1400,1401
_|1401,1402
at|1403,1405
_|1406,1407
_|1407,1408
_|1408,1409
_|1410,1411
_|1411,1412
_|1412,1413
-|1414,1415
<EOL>|1417,1418
_|1418,1419
_|1419,1420
_|1420,1421
wound|1422,1427
revision|1428,1436
and|1437,1440
removal|1441,1448
of|1449,1451
the|1452,1455
exposed|1456,1463
craniotx|1464,1472
<EOL>|1473,1474
hardware|1474,1482
,|1482,1483
Accutane|1484,1492
for|1493,1496
2|1497,1498
weeks|1499,1504
only|1505,1509
_|1510,1511
_|1511,1512
_|1512,1513
disease|1514,1521
since|1522,1527
<EOL>|1528,1529
_|1529,1530
_|1530,1531
_|1531,1532
,|1532,1533
<EOL>|1535,1536
tubal|1536,1541
ligation|1542,1550
,|1550,1551
tonsillectomy|1551,1564
,|1564,1565
bronchitis|1566,1576
,|1576,1577
depression|1578,1588
.|1588,1589
<EOL>|1591,1592
seizures|1592,1600
<EOL>|1602,1603
<EOL>|1603,1604
<EOL>|1605,1606
:|1620,1621
<EOL>|1621,1622
_|1622,1623
_|1623,1624
_|1624,1625
<EOL>|1625,1626
:|1640,1641
<EOL>|1641,1642
NC|1642,1644
<EOL>|1644,1645
<EOL>|1646,1647
AF|1662,1664
VSS|1665,1668
<EOL>|1668,1669
obese|1669,1674
<EOL>|1674,1675
Gen|1675,1678
:|1678,1679
WD|1680,1682
/|1682,1683
WN|1683,1685
,|1685,1686
comfortable|1687,1698
,|1698,1699
NAD|1700,1703
.|1703,1704
<EOL>|1704,1705
HEENT|1705,1710
:|1710,1711
_|1712,1713
_|1713,1714
_|1714,1715
bilat|1716,1721
EOMs|1722,1726
:|1726,1727
intact|1728,1734
<EOL>|1734,1735
Neck|1735,1739
:|1739,1740
Supple|1741,1747
.|1747,1748
<EOL>|1748,1749
no|1749,1751
LNN|1752,1755
<EOL>|1755,1756
RRR|1756,1759
<EOL>|1759,1760
no|1760,1762
SOB|1763,1766
<EOL>|1766,1767
obese|1767,1772
<EOL>|1772,1773
Extrem|1773,1779
:|1779,1780
Warm|1781,1785
and|1786,1789
well|1790,1794
-|1794,1795
perfused|1795,1803
,|1803,1804
<EOL>|1805,1806
<EOL>|1806,1807
Neuro|1807,1812
:|1812,1813
<EOL>|1813,1814
Mental|1814,1820
status|1821,1827
:|1827,1828
Awake|1829,1834
and|1835,1838
alert|1839,1844
,|1844,1845
cooperative|1846,1857
with|1858,1862
exam|1863,1867
,|1867,1868
normal|1869,1875
<EOL>|1875,1876
affect|1876,1882
but|1883,1886
VERY|1887,1891
simple|1892,1898
construct|1899,1908
.|1908,1909
<EOL>|1909,1910
Orientation|1910,1921
:|1921,1922
Oriented|1923,1931
to|1932,1934
person|1935,1941
,|1941,1942
place|1943,1948
,|1948,1949
and|1950,1953
date|1954,1958
.|1958,1959
<EOL>|1959,1960
Recall|1960,1966
:|1966,1967
_|1968,1969
_|1969,1970
_|1970,1971
objects|1972,1979
at|1980,1982
5|1983,1984
minutes|1985,1992
.|1992,1993
<EOL>|1993,1994
Language|1994,2002
:|2002,2003
Speech|2004,2010
fluent|2011,2017
with|2018,2022
good|2023,2027
comprehension|2028,2041
and|2042,2045
repetition|2046,2056
.|2056,2057
<EOL>|2057,2058
Naming|2058,2064
intact|2065,2071
.|2071,2072
No|2073,2075
dysarthria|2076,2086
or|2087,2089
paraphasic|2090,2100
errors|2101,2107
.|2107,2108
<EOL>|2108,2109
<EOL>|2109,2110
Cranial|2110,2117
Nerves|2118,2124
:|2124,2125
<EOL>|2125,2126
I|2126,2127
:|2127,2128
Not|2129,2132
tested|2133,2139
<EOL>|2139,2140
II|2140,2142
:|2142,2143
Pupils|2144,2150
equally|2151,2158
round|2159,2164
and|2165,2168
reactive|2169,2177
to|2178,2180
light|2181,2186
,|2186,2187
3|2189,2190
to|2191,2193
2|2194,2195
<EOL>|2195,2196
mm|2196,2198
bilaterally|2199,2210
.|2210,2211
Visual|2212,2218
fields|2219,2225
are|2226,2229
full|2230,2234
to|2235,2237
confrontation|2238,2251
.|2251,2252
<EOL>|2252,2253
III|2253,2256
,|2256,2257
IV|2258,2260
,|2260,2261
VI|2262,2264
:|2264,2265
Extraocular|2266,2277
movements|2278,2287
intact|2288,2294
bilaterally|2295,2306
without|2307,2314
<EOL>|2314,2315
nystagmus|2315,2324
.|2324,2325
<EOL>|2325,2326
V|2326,2327
,|2327,2328
VII|2329,2332
:|2332,2333
Facial|2334,2340
strength|2341,2349
and|2350,2353
sensation|2354,2363
intact|2364,2370
and|2371,2374
symmetric|2375,2384
.|2384,2385
<EOL>|2385,2386
VIII|2386,2390
:|2390,2391
Hearing|2392,2399
intact|2400,2406
to|2407,2409
voice|2410,2415
.|2415,2416
<EOL>|2416,2417
IX|2417,2419
,|2419,2420
X|2421,2422
:|2422,2423
Palatal|2424,2431
elevation|2432,2441
symmetrical|2442,2453
.|2453,2454
<EOL>|2454,2455
XI|2455,2457
:|2457,2458
Sternocleidomastoid|2459,2478
and|2479,2482
trapezius|2483,2492
normal|2493,2499
bilaterally|2500,2511
.|2511,2512
<EOL>|2512,2513
XII|2513,2516
:|2516,2517
Tongue|2518,2524
midline|2525,2532
without|2533,2540
fasciculations|2541,2555
.|2555,2556
<EOL>|2556,2557
<EOL>|2557,2558
Motor|2558,2563
:|2563,2564
Normal|2565,2571
bulk|2572,2576
and|2577,2580
tone|2581,2585
bilaterally|2586,2597
.|2597,2598
No|2599,2601
abnormal|2602,2610
movements|2611,2620
<EOL>|2620,2621
<EOL>|2621,2622
W|2622,2623
:|2623,2624
there|2625,2630
is|2631,2633
an|2634,2636
area|2637,2641
over|2642,2646
the|2647,2650
R|2651,2652
hemiconvexity|2653,2666
that|2667,2671
shows|2672,2677
a|2678,2679
<EOL>|2680,2681
chronic|2681,2688
<EOL>|2688,2689
skin|2689,2693
defect|2694,2700
where|2701,2706
the|2707,2710
underlying|2711,2721
harware|2722,2729
has|2730,2733
eroded|2734,2740
through|2741,2748
the|2749,2752
<EOL>|2752,2753
skin|2753,2757
.|2757,2758
<EOL>|2758,2759
Different|2759,2768
from|2769,2773
previous|2774,2782
repaired|2783,2791
portion|2792,2799
and|2800,2803
represents|2804,2814
piece|2815,2820
of|2821,2823
<EOL>|2824,2825
the|2825,2828
implanted|2829,2838
miniplates|2839,2849
;|2849,2850
No|2851,2853
discharge|2854,2863
;|2863,2864
no|2865,2867
reythemal|2868,2877
no|2878,2880
<EOL>|2881,2882
swelling|2882,2890
;|2890,2891
surprisingly|2893,2905
benign|2906,2912
aspect|2913,2919
.|2919,2920
<EOL>|2920,2921
<EOL>|2921,2922
PHYSICAL|2922,2930
EXAM|2931,2935
PRIOR|2936,2941
TO|2942,2944
DISCHARGE|2945,2954
:|2954,2955
<EOL>|2956,2957
AF|2957,2959
VSS|2960,2963
<EOL>|2963,2964
obese|2964,2969
<EOL>|2969,2970
Gen|2970,2973
:|2973,2974
WD|2975,2977
/|2977,2978
WN|2978,2980
,|2980,2981
comfortable|2982,2993
,|2993,2994
NAD|2995,2998
.|2998,2999
<EOL>|2999,3000
HEENT|3000,3005
:|3005,3006
_|3007,3008
_|3008,3009
_|3009,3010
bilat|3011,3016
EOMs|3017,3021
:|3021,3022
intact|3023,3029
<EOL>|3029,3030
Neck|3030,3034
:|3034,3035
Supple|3036,3042
.|3042,3043
<EOL>|3043,3044
Incision|3044,3052
:|3052,3053
clean|3054,3059
,|3059,3060
dry|3061,3064
,|3064,3065
intact|3066,3072
.|3072,3073
No|3074,3076
redness|3077,3084
,|3084,3085
swelling|3086,3094
,|3094,3095
erythema|3096,3104
or|3105,3107
<EOL>|3108,3109
discharge|3109,3118
.|3118,3119
Sutures|3120,3127
in|3128,3130
place|3131,3136
.|3136,3137
<EOL>|3138,3139
<EOL>|3140,3141
Pertinent|3141,3150
Results|3151,3158
:|3158,3159
<EOL>|3159,3160
_|3160,3161
_|3161,3162
_|3162,3163
:|3163,3164
<EOL>|3164,3165
Hematology|3165,3175
<EOL>|3176,3177
COMPLETE|3177,3185
BLOOD|3186,3191
COUNT|3192,3197
WBC|3198,3201
RBC|3202,3205
Hgb|3206,3209
Hct|3210,3213
MCV|3214,3217
MCH|3218,3221
MCHC|3222,3226
RDW|3227,3230
Plt|3231,3234
Ct|3235,3237
<EOL>|3238,3239
_|3239,3240
_|3240,3241
_|3241,3242
06|3243,3245
:|3245,3246
25|3246,3248
4.8|3252,3255
3.49|3256,3260
*|3260,3261
11.2|3262,3266
*|3266,3267
34.4|3268,3272
*|3272,3273
98|3274,3276
31.9|3277,3281
32.5|3282,3286
16.3|3287,3291
*|3291,3292
245|3293,3296
<EOL>|3297,3298
<EOL>|3298,3299
BASIC|3299,3304
COAGULATION|3305,3316
_|3317,3318
_|3318,3319
_|3319,3320
,|3320,3321
PTT|3322,3325
,|3325,3326
PLT|3327,3330
,|3330,3331
INR|3332,3335
)|3335,3336
Plt|3337,3340
Ct|3341,3343
<EOL>|3344,3345
_|3345,3346
_|3346,3347
_|3347,3348
06|3349,3351
:|3351,3352
25|3352,3354
245|3358,3361
<EOL>|3362,3363
<EOL>|3364,3365
Chemistry|3365,3374
<EOL>|3375,3376
RENAL|3376,3381
&|3382,3383
GLUCOSE|3384,3391
Glucose|3392,3399
UreaN|3400,3405
Creat|3406,3411
Na|3412,3414
K|3415,3416
Cl|3417,3419
HCO3|3420,3424
AnGap|3425,3430
<EOL>|3431,3432
_|3432,3433
_|3433,3434
_|3434,3435
06|3436,3438
:|3438,3439
25|3439,3441
_|3445,3446
_|3446,3447
_|3447,3448
142|3449,3452
3.4|3453,3456
110|3457,3460
*|3460,3461
23|3462,3464
12|3465,3467
<EOL>|3468,3469
<EOL>|3469,3470
<EOL>|3471,3472
<EOL>|3472,3473
<EOL>|3474,3475
The|3498,3501
patient|3502,3509
presented|3510,3519
to|3520,3522
the|3523,3526
_|3527,3528
_|3528,3529
_|3529,3530
neurosurgical|3531,3544
service|3545,3552
on|3553,3555
<EOL>|3556,3557
_|3557,3558
_|3558,3559
_|3559,3560
for|3561,3564
treatment|3565,3574
of|3575,3577
exposed|3578,3585
hardware|3586,3594
from|3595,3599
a|3600,3601
previous|3602,3610
<EOL>|3611,3612
surgery|3612,3619
on|3620,3622
her|3623,3626
head|3627,3631
.|3631,3632
She|3633,3636
went|3637,3641
to|3642,3644
the|3645,3648
OR|3649,3651
on|3652,3654
_|3655,3656
_|3656,3657
_|3657,3658
,|3658,3659
where|3660,3665
a|3666,3667
<EOL>|3669,3670
was|3670,3673
performed|3674,3683
removal|3684,3691
of|3692,3694
exposed|3695,3702
hardware|3703,3711
by|3712,3714
Dr.|3715,3718
_|3719,3720
_|3720,3721
_|3721,3722
.|3722,3723
<EOL>|3724,3725
Postoperatively|3725,3740
,|3740,3741
the|3742,3745
patient|3746,3753
was|3754,3757
stable|3758,3764
.|3764,3765
Infectious|3766,3776
disease|3777,3784
<EOL>|3785,3786
consulted|3786,3795
the|3796,3799
patient|3800,3807
and|3808,3811
recommended|3812,3823
fluconazole|3824,3835
200|3836,3839
mg|3840,3842
PO|3843,3845
for|3846,3849
<EOL>|3850,3851
5|3851,3852
days|3853,3857
for|3858,3861
yeast|3862,3867
infection|3868,3877
and|3878,3881
Keflex|3882,3888
_|3889,3890
_|3890,3891
_|3891,3892
mg|3893,3895
PO|3896,3898
BID|3899,3902
for|3903,3906
7|3907,3908
days|3909,3913
.|3913,3914
<EOL>|3914,3915
<EOL>|3915,3916
For|3916,3919
DVT|3920,3923
prophylaxis|3924,3935
,|3935,3936
the|3937,3940
patient|3941,3948
received|3949,3957
subcutaneous|3958,3970
heparin|3971,3978
<EOL>|3979,3980
and|3980,3983
SCD|3984,3987
's|3987,3989
during|3990,3996
her|3997,4000
stay|4001,4005
.|4005,4006
<EOL>|4006,4007
<EOL>|4007,4008
At|4008,4010
the|4011,4014
time|4015,4019
of|4020,4022
discharge|4023,4032
,|4032,4033
the|4034,4037
patient|4038,4045
was|4046,4049
able|4050,4054
to|4055,4057
tolerate|4058,4066
PO|4067,4069
,|4069,4070
<EOL>|4071,4072
was|4072,4075
ambulatoryand|4076,4089
able|4090,4094
to|4095,4097
void|4098,4102
independently|4103,4116
.|4116,4117
She|4118,4121
was|4122,4125
able|4126,4130
to|4131,4133
<EOL>|4134,4135
verbalize|4135,4144
agreement|4145,4154
and|4155,4158
understanding|4159,4172
of|4173,4175
the|4176,4179
discharge|4180,4189
plan|4190,4194
.|4194,4195
<EOL>|4195,4196
<EOL>|4197,4198
Medications|4198,4209
on|4210,4212
Admission|4213,4222
:|4222,4223
<EOL>|4223,4224
The|4224,4227
Preadmission|4228,4240
Medication|4241,4251
list|4252,4256
may|4257,4260
be|4261,4263
inaccurate|4264,4274
and|4275,4278
requires|4279,4287
<EOL>|4288,4289
futher|4289,4295
investigation|4296,4309
.|4309,4310
<EOL>|4310,4311
1.|4311,4313
ALPRAZolam|4314,4324
0.5|4325,4328
mg|4329,4331
PO|4332,4334
TID|4335,4338
<EOL>|4339,4340
2.|4340,4342
Azathioprine|4343,4355
100|4356,4359
mg|4360,4362
PO|4363,4365
BID|4366,4369
<EOL>|4370,4371
3.|4371,4373
DiCYCLOmine|4374,4385
10|4386,4388
mg|4389,4391
PO|4392,4394
Q6H|4395,4398
:|4398,4399
PRN|4399,4402
abdominal|4403,4412
pain|4413,4417
<EOL>|4418,4419
4.|4419,4421
Fluticasone|4422,4433
-|4433,4434
Salmeterol|4434,4444
Diskus|4445,4451
(|4452,4453
500|4453,4456
/|4456,4457
50|4457,4459
)|4459,4460
1|4462,4463
INH|4464,4467
IH|4468,4470
BID|4471,4474
<EOL>|4475,4476
5.|4476,4478
Hydrocodone|4479,4490
-|4490,4491
Acetaminophen|4491,4504
(|4505,4506
5mg|4506,4509
-|4509,4510
500mg|4510,4515
)|4515,4516
1|4517,4518
TAB|4519,4522
PO|4523,4525
Q4H|4526,4529
:|4529,4530
PRN|4530,4533
pain|4534,4538
<EOL>|4539,4540
6.|4540,4542
Infliximab|4543,4553
100|4554,4557
mg|4558,4560
IV|4561,4563
Q6|4564,4566
WEEKS|4567,4572
<EOL>|4573,4574
7.|4574,4576
Levothyroxine|4577,4590
Sodium|4591,4597
50|4598,4600
mcg|4601,4604
PO|4605,4607
DAILY|4608,4613
<EOL>|4614,4615
8.|4615,4617
Mesalamine|4618,4628
500|4629,4632
mg|4633,4635
PO|4636,4638
QID|4639,4642
<EOL>|4643,4644
9.|4644,4646
Omeprazole|4647,4657
20|4658,4660
mg|4661,4663
PO|4664,4666
DAILY|4667,4672
<EOL>|4673,4674
10.|4674,4677
Promethazine|4678,4690
25|4691,4693
mg|4694,4696
PO|4697,4699
Q6H|4700,4703
:|4703,4704
PRN|4704,4707
n|4708,4709
/|4709,4710
v|4710,4711
<EOL>|4712,4713
11|4713,4715
.|4715,4716
Topiramate|4717,4727
(|4728,4729
Topamax|4729,4736
)|4736,4737
200|4738,4741
mg|4742,4744
PO|4745,4747
BID|4748,4751
<EOL>|4752,4753
12.|4753,4756
Venlafaxine|4757,4768
XR|4769,4771
150|4772,4775
mg|4776,4778
PO|4779,4781
DAILY|4782,4787
<EOL>|4788,4789
13.|4789,4792
Zolpidem|4793,4801
Tartrate|4802,4810
15|4811,4813
mg|4814,4816
PO|4817,4819
HS|4820,4822
<EOL>|4823,4824
<EOL>|4824,4825
<EOL>|4826,4827
Discharge|4827,4836
Medications|4837,4848
:|4848,4849
<EOL>|4849,4850
1.|4850,4852
ALPRAZolam|4853,4863
0.5|4864,4867
mg|4868,4870
PO|4871,4873
TID|4874,4877
<EOL>|4878,4879
2.|4879,4881
Azathioprine|4882,4894
100|4895,4898
mg|4899,4901
PO|4902,4904
BID|4905,4908
<EOL>|4909,4910
3.|4910,4912
DiCYCLOmine|4913,4924
10|4925,4927
mg|4928,4930
PO|4931,4933
Q6H|4934,4937
:|4937,4938
PRN|4938,4941
abdominal|4942,4951
pain|4952,4956
<EOL>|4957,4958
4.|4958,4960
Levothyroxine|4961,4974
Sodium|4975,4981
50|4982,4984
mcg|4985,4988
PO|4989,4991
DAILY|4992,4997
<EOL>|4998,4999
5.|4999,5001
Mesalamine|5002,5012
500|5013,5016
mg|5017,5019
PO|5020,5022
QID|5023,5026
<EOL>|5027,5028
6.|5028,5030
Omeprazole|5031,5041
20|5042,5044
mg|5045,5047
PO|5048,5050
DAILY|5051,5056
<EOL>|5057,5058
7.|5058,5060
Topiramate|5061,5071
(|5072,5073
Topamax|5073,5080
)|5080,5081
200|5082,5085
mg|5086,5088
PO|5089,5091
BID|5092,5095
<EOL>|5096,5097
8.|5097,5099
Venlafaxine|5100,5111
XR|5112,5114
150|5115,5118
mg|5119,5121
PO|5122,5124
DAILY|5125,5130
<EOL>|5131,5132
9.|5132,5134
Zolpidem|5135,5143
Tartrate|5144,5152
15|5153,5155
mg|5156,5158
PO|5159,5161
HS|5162,5164
<EOL>|5165,5166
10.|5166,5169
Hydrocodone|5170,5181
-|5181,5182
Acetaminophen|5182,5195
(|5196,5197
5mg|5197,5200
-|5200,5201
500mg|5201,5206
)|5206,5207
1|5208,5209
TAB|5210,5213
PO|5214,5216
Q4H|5217,5220
:|5220,5221
PRN|5221,5224
pain|5225,5229
<EOL>|5230,5231
11|5231,5233
.|5233,5234
Acetaminophen|5235,5248
325|5249,5252
-|5252,5253
650|5253,5256
mg|5257,5259
PO|5260,5262
Q6H|5263,5266
:|5266,5267
PRN|5267,5270
temperature|5271,5282
;|5282,5283
pain|5284,5288
<EOL>|5289,5290
12.|5290,5293
Docusate|5294,5302
Sodium|5303,5309
100|5310,5313
mg|5314,5316
PO|5317,5319
BID|5320,5323
:|5323,5324
PRN|5324,5327
constipation|5328,5340
<EOL>|5341,5342
RX|5342,5344
*|5345,5346
docusate|5346,5354
sodium|5355,5361
100|5362,5365
mg|5366,5368
100|5369,5372
capsule|5373,5380
(|5380,5381
s|5381,5382
)|5382,5383
by|5384,5386
mouth|5387,5392
twice|5393,5398
a|5399,5400
day|5401,5404
<EOL>|5405,5406
Disp|5406,5410
#|5411,5412
*|5412,5413
30|5413,5415
Capsule|5416,5423
Refills|5424,5431
:|5431,5432
*|5432,5433
0|5433,5434
<EOL>|5434,5435
13.|5435,5438
Fluconazole|5439,5450
200|5451,5454
mg|5455,5457
PO|5458,5460
Q24H|5461,5465
Duration|5466,5474
:|5474,5475
4|5476,5477
Days|5478,5482
<EOL>|5483,5484
RX|5484,5486
*|5487,5488
fluconazole|5488,5499
200|5500,5503
mg|5504,5506
1|5507,5508
tablet|5509,5515
(|5515,5516
s|5516,5517
)|5517,5518
by|5519,5521
mouth|5522,5527
daily|5528,5533
Disp|5534,5538
#|5539,5540
*|5540,5541
4|5541,5542
<EOL>|5543,5544
Tablet|5544,5550
Refills|5551,5558
:|5558,5559
*|5559,5560
0|5560,5561
<EOL>|5561,5562
14.|5562,5565
OxycoDONE|5566,5575
(|5576,5577
Immediate|5577,5586
Release|5587,5594
)|5594,5595
5|5597,5598
mg|5599,5601
PO|5602,5604
Q6H|5605,5608
:|5608,5609
PRN|5609,5612
for|5613,5616
moderate|5617,5625
<EOL>|5626,5627
pain|5627,5631
<EOL>|5632,5633
RX|5633,5635
*|5636,5637
oxycodone|5637,5646
5|5647,5648
mg|5649,5651
_|5652,5653
_|5653,5654
_|5654,5655
tablet|5656,5662
(|5662,5663
s|5663,5664
)|5664,5665
by|5666,5668
mouth|5669,5674
every|5675,5680
six|5681,5684
(|5685,5686
6|5686,5687
)|5687,5688
hours|5689,5694
<EOL>|5695,5696
Disp|5696,5700
#|5701,5702
*|5702,5703
40|5703,5705
Tablet|5706,5712
Refills|5713,5720
:|5720,5721
*|5721,5722
0|5722,5723
<EOL>|5723,5724
15.|5724,5727
Cephalexin|5728,5738
500|5739,5742
mg|5743,5745
PO|5746,5748
Q12H|5749,5753
Duration|5754,5762
:|5762,5763
7|5764,5765
Days|5766,5770
<EOL>|5771,5772
RX|5772,5774
*|5775,5776
cephalexin|5776,5786
500|5787,5790
mg|5791,5793
1|5794,5795
tablet|5796,5802
(|5802,5803
s|5803,5804
)|5804,5805
by|5806,5808
mouth|5809,5814
twice|5815,5820
a|5821,5822
day|5823,5826
Disp|5827,5831
#|5832,5833
*|5833,5834
14|5834,5836
<EOL>|5837,5838
Tablet|5838,5844
Refills|5845,5852
:|5852,5853
*|5853,5854
0|5854,5855
<EOL>|5855,5856
<EOL>|5856,5857
<EOL>|5858,5859
Discharge|5859,5868
Disposition|5869,5880
:|5880,5881
<EOL>|5881,5882
Home|5882,5886
<EOL>|5886,5887
<EOL>|5888,5889
Discharge|5889,5898
Diagnosis|5899,5908
:|5908,5909
<EOL>|5909,5910
Hardware|5910,5918
removal|5919,5926
<EOL>|5926,5927
<EOL>|5927,5928
<EOL>|5929,5930
Mental|5951,5957
Status|5958,5964
:|5964,5965
Clear|5966,5971
and|5972,5975
coherent|5976,5984
.|5984,5985
<EOL>|5985,5986
Level|5986,5991
of|5992,5994
Consciousness|5995,6008
:|6008,6009
Alert|6010,6015
and|6016,6019
interactive|6020,6031
.|6031,6032
<EOL>|6032,6033
Activity|6033,6041
Status|6042,6048
:|6048,6049
Ambulatory|6050,6060
-|6061,6062
Independent|6063,6074
.|6074,6075
<EOL>|6075,6076
<EOL>|6076,6077
<EOL>|6078,6079
|6103,6104
Please|6105,6111
take|6112,6116
Fluconazole|6117,6128
200mg|6129,6134
once|6135,6139
daily|6140,6145
for|6146,6149
4|6150,6151
days|6152,6156
.|6156,6157
Please|6158,6164
<EOL>|6165,6166
take|6166,6170
Keflex|6171,6177
for|6178,6181
7|6182,6183
days|6184,6188
for|6189,6192
wound|6193,6198
infection|6199,6208
.|6208,6209
<EOL>|6210,6211
<EOL>|6211,6212
Clearance|6212,6221
to|6222,6224
drive|6225,6230
and|6231,6234
return|6235,6241
to|6242,6244
work|6245,6249
will|6250,6254
be|6255,6257
addressed|6258,6267
at|6268,6270
your|6271,6275
<EOL>|6276,6277
post-operative|6277,6291
office|6292,6298
visit|6299,6304
.|6304,6305
<EOL>|6305,6306
CALL|6306,6310
YOUR|6311,6315
SURGEON|6316,6323
IMMEDIATELY|6324,6335
IF|6336,6338
YOU|6339,6342
EXPERIENCE|6343,6353
ANY|6354,6357
OF|6358,6360
THE|6361,6364
<EOL>|6365,6366
FOLLOWING|6366,6375
<EOL>|6375,6376
<EOL>|6376,6377
|6377,6378
New|6378,6381
onset|6382,6387
of|6388,6390
tremors|6391,6398
or|6399,6401
seizures|6402,6410
.|6410,6411
<EOL>|6411,6412
|6412,6413
Any|6413,6416
confusion|6417,6426
or|6427,6429
change|6430,6436
in|6437,6439
mental|6440,6446
status|6447,6453
.|6453,6454
<EOL>|6455,6456
|6456,6457
Any|6457,6460
numbness|6461,6469
,|6469,6470
tingling|6471,6479
,|6479,6480
weakness|6481,6489
in|6490,6492
your|6493,6497
extremities|6498,6509
.|6509,6510
<EOL>|6510,6511
|6511,6512
Pain|6512,6516
or|6517,6519
headache|6520,6528
that|6529,6533
is|6534,6536
continually|6537,6548
increasing|6549,6559
,|6559,6560
or|6561,6563
not|6564,6567
<EOL>|6568,6569
relieved|6569,6577
by|6578,6580
pain|6581,6585
medication|6586,6596
.|6596,6597
<EOL>|6597,6598
|6598,6599
Any|6599,6602
signs|6603,6608
of|6609,6611
infection|6612,6621
at|6622,6624
the|6625,6628
wound|6629,6634
site|6635,6639
:|6639,6640
increasing|6641,6651
redness|6652,6659
,|6659,6660
<EOL>|6661,6662
increased|6662,6671
swelling|6672,6680
,|6680,6681
increased|6682,6691
tenderness|6692,6702
,|6702,6703
or|6704,6706
drainage|6707,6715
.|6715,6716
<EOL>|6716,6717
|6717,6718
Fever|6718,6723
greater|6724,6731
than|6732,6736
or|6737,6739
equal|6740,6745
to|6746,6748
101|6749,6752
.|6752,6753
5|6753,6754
°|6754,6755
F|6756,6757
.|6757,6758
<EOL>|6758,6759
<EOL>|6759,6760
<EOL>|6761,6762
Followup|6762,6770
Instructions|6771,6783
:|6783,6784
<EOL>|6784,6785
_|6785,6786
_|6786,6787
_|6787,6788
<EOL>|6788,6789

