CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Sulfonamides, ophthalmologic antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamides
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamides
null|Sulfonamides, topical|Drug|false|false||Sulfonamides
null|Sulfonamides|Drug|false|false||Sulfonamides
null|Sulfonamides|Drug|false|false||Sulfonamides
null|Sulfonamides, ophthalmologic antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamides, Gynecological|Drug|false|false||Sulfonamides
null|Sulfonamides, Gynecological|Drug|false|false||Sulfonamides
null|Sulfonamides, intestinal antiinfectives|Drug|false|false||Sulfonamides
null|Sulfonamides, intestinal antiinfectives|Drug|false|false||Sulfonamidesnull|Poisoning by, adverse effect of and underdosing of sulfonamides|Disorder|false|false||Sulfonamides
null|Poisoning by sulfonamide|Disorder|false|false||Sulfonamidesnull|Adverse reaction to sulfonamides|Finding|false|false||Sulfonamidesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Bactrim|Drug|false|false||Bactrim
null|Bactrim|Drug|false|false||Bactrimnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Vomiting|Finding|false|false||vomitingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Exploratory laparotomy|Procedure|false|false||Exploratory laparotomynull|Laparotomy|Procedure|false|false||laparotomynull|Lysis of adhesions|Procedure|false|false||lysis of adhesionsnull|Lysis|Finding|false|false||lysis
null|pathologic cytolysis|Finding|false|false||lysisnull|Tissue Adhesions|Finding|false|false||adhesionsnull|Small|LabModifier|false|false||smallnull|Bowel resection|Procedure|false|false|C0021853|bowel resectionnull|Intestines|Anatomy|false|false|C0741614;C0015252;C0728940|bowelnull|removal technique|Procedure|false|false|C0021853|resection
null|Excision|Procedure|false|false|C0021853|resectionnull|Anastomosis of small intestine to small intestine|Procedure|false|false||enteroenterostomy
null|Anastomosis of intestine|Procedure|false|false||enteroenterostomynull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Uterus|Anatomy|false|false||uterinenull|Uterine Fibroids|Disorder|false|false||fibroids
null|Fibroid Tumor|Disorder|false|false||fibroidsnull|Lung excision|Procedure|false|false|C4037972;C0024109|lung resectionnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0024115;C0396565;C0740941|lung
null|Lung|Anatomy|false|false|C0024115;C0396565;C0740941|lungnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Carcinoid Tumor|Disorder|false|false||carcinoid tumornull|Carcinoid Tumor|Disorder|false|false||carcinoidnull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Surgical consultation|Procedure|false|false||surgical consultationnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Diagnosis Classification - Consultation|Finding|false|false||consultation
null|Document Type - Consultation|Finding|false|false||consultationnull|Consultation|Procedure|false|false||consultationnull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Early|Time|false|false||earlynull|Morning|Time|false|false||morningnull|Approximate|Modifier|false|false||approximatelynull|Muscle Cramp|Finding|false|false|C0000726|crampingnull|Cramping sensation quality|Modifier|false|false||crampingnull|Abdomen|Anatomy|false|false|C0026821|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Associated with|Modifier|false|false||associated withnull|Associated with|Modifier|false|false||associatednull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting bile|Finding|false|false||bilious emesisnull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Approximate|Modifier|false|false||approximatelynull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Presentation|Finding|false|false||presentationnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Intestines|Anatomy|false|false|C5975557|bowelsnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false|C0021853|timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Similarity|Modifier|false|false||similarnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Small bowel obstruction|Disorder|false|false|C4319010;C0021852;C0021853|small bowel obstructionnull|Abdomen>Small bowel|Anatomy|false|false|C0021843;C0235329;C0028778|small bowel
null|Intestines, Small|Anatomy|false|false|C0021843;C0235329;C0028778|small bowelnull|Small|LabModifier|false|false||smallnull|Intestinal Obstruction|Disorder|false|false|C4319010;C0021852;C0021853|bowel obstructionnull|Intestines|Anatomy|false|false|C0021843;C0028778;C0235329|bowelnull|Obstruction|Finding|false|false|C0021853;C4319010;C0021852|obstructionnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|Carcinoid Tumor|Disorder|false|false||carcinoid tumornull|Carcinoid Tumor|Disorder|false|false||carcinoidnull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Vitamin B 12 Deficiency|Disorder|false|false||Vitamin B12 deficiencynull|Decreased circulating vitamin B12 concentration|Finding|false|false||Vitamin B12 deficiencynull|Vitamin B12 [EPC]|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|cobalamins|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12
null|vitamin B12|Drug|false|false||Vitamin B12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||Vitamin B12null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Lung excision|Procedure|false|false|C4037972;C0024109|lung resectionnull|Lung diseases|Disorder|false|false|C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0396565;C0024115;C0740941|lung
null|Lung|Anatomy|false|false|C0396565;C0024115;C0740941|lungnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Right arm|Anatomy|false|false|C3495676;C0038895;C1457907;C1547138;C0543467;C1824218;C3715044;C1522541;C5400986;C4761640|R armnull|Anorectal Malformations|Disorder|false|false|C4048756;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078;C4048756|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078;C4048756|armnull|Protocol Treatment Arm|Procedure|false|false|C0446516;C1140618;C1269078;C4048756|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0446516;C1140618;C1269078;C4048756|arm
null|Study Arm|Procedure|false|false|C0446516;C1140618;C1269078;C4048756|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|null|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C3495676;C1522541;C5400986;C4761640|armnull|Level of Care - Surgery|Finding|false|false|C4048756|surgery
null|Surgical procedure finding|Finding|false|false|C4048756|surgery
null|Surgical aspects|Finding|false|false|C4048756|surgerynull|Operative Surgical Procedures|Procedure|false|false|C4048756|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Contribution|Event|false|false||contributorynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heartnull|Regular|Modifier|false|false||regularnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|false|false|C0004339;C1550016|lungsnull|Remote control command - Clear|Finding|false|false|C0024109|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Auscultation|Procedure|false|false|C0024109|auscultationnull|Decreased breath sounds|Finding|false|false||decreased breath soundsnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Thoracotomy Scar|Finding|false|false||thoracotomy scarnull|Thoracotomy|Procedure|false|false||thoracotomynull|Scar Tissue|Finding|false|false||scar
null|Cicatrix|Finding|false|false||scar
null|RPS4X gene|Finding|false|false||scarnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Abdomen soft|Finding|false|false|C0230168;C0000726|abdomen softnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0426663;C0153662;C0941288;C3542022|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0426663;C0153662;C0941288;C3542022|abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0230168;C0000726|softnull|Soft|Modifier|false|false||softnull|Very|Modifier|false|false||verynull|Obesity|Disorder|false|false||obesenull|Dilated|Finding|false|false||distendednull|Distended|Modifier|false|false||distendednull|Somewhat|Finding|false|false||somewhatnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|abdomennull|Protective muscle spasm|Finding|true|false||guardingnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|IPSS-R Risk Category Low|Finding|false|false|C1660780|low
null|IPSS Risk Category Low|Finding|false|false|C1660780|low
null|low confidentiality|Finding|false|false|C1660780|lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|midline cell component|Anatomy|false|false|C4510895;C3263723;C0043251;C0043250;C5203106;C4522223;C1550472;C1549529;C1547965;C1550680|midlinenull|Midline (qualifier value)|Modifier|false|false||midlinenull|Wound of abdomen|Disorder|false|false|C1660780;C0000726|abdominal woundnull|Abdomen|Anatomy|false|false|C4510895;C3263723;C0043251;C0043250|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Traumatic Wound|Disorder|false|false|C1660780;C0000726|wound
null|Wounds and Injuries|Disorder|false|false|C1660780;C0000726|wound
null|Traumatic injury|Disorder|false|false|C1660780;C0000726|woundnull|Route of Administration - Wound|Finding|false|false|C1660780|wound
null|null|Finding|false|false|C1660780|wound
null|Specimen Type - Wound|Finding|false|false|C1660780|woundnull|Body Substance Discharge|Finding|true|false||drainage
null|Body Fluid Discharge|Finding|true|false||drainagenull|Drainage procedure|Procedure|true|false||drainagenull|Erythema|Disorder|false|false||erythemanull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C4522245;C1415181;C1420113;C5960784;C1415181;C0201899;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|CT of abdomen and pelvis|Procedure|false|false|C4266535;C0030797;C0559769;C0230168;C0000726;C1508499;C0000726|CT of abdomen and pelvisnull|CT of abdomen|Procedure|false|false|C0230168;C0000726|CT of abdomennull|Abdominopelvic structure|Anatomy|false|false|C0812455;C1641132;C0941288;C0153662;C0153663|abdomen and pelvisnull|Abdomen|Anatomy|false|false|C0941288;C0153663;C0812455;C1641132;C0153662|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C1508499;C0000726;C0230168;C0000726;C4266535;C0030797;C0559769|abdomennull|Abdomen problem|Finding|false|false|C1508499;C0230168;C0000726;C0000726|abdomennull|Abdomen|Anatomy|false|false|C1641132;C0412620;C0941288;C0812455;C0153662;C0153663|abdomen
null|Abdominal Cavity|Anatomy|false|false|C1641132;C0412620;C0941288;C0812455;C0153662;C0153663|abdomennull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769;C0000726;C1508499;C0230168;C0000726|pelvisnull|Pelvis problem|Finding|false|false|C1508499;C4266535;C0030797;C0559769;C0000726;C0230168;C0000726|pelvisnull|Pelvis+|Anatomy|false|false|C1641132;C0812455;C0153663;C0153662|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C1641132;C0812455;C0153663;C0153662|pelvis
null|Pelvis|Anatomy|false|false|C1641132;C0812455;C0153663;C0153662|pelvisnull|Slightly (qualifier value)|Modifier|false|false||Slightly
null|Slight (qualifier value)|Modifier|false|false||Slightlynull|Dilated loops|Finding|false|false||dilated loopsnull|Dilated|Finding|false|false||dilatednull|null|Device|false|false||loopsnull|Abdomen>Small bowel|Anatomy|false|false|C1552853;C0456205;C1546561|small bowel
null|Intestines, Small|Anatomy|false|false|C1552853;C0456205;C1546561|small bowelnull|Small|LabModifier|false|false||smallnull|Intestines|Anatomy|false|false|C1546561;C1552853;C0456205|bowelnull|Abdomen>Small bowel|Anatomy|false|false|C1552853;C0456205;C1546561|small bowel
null|Intestines, Small|Anatomy|false|false|C1552853;C0456205;C1546561|small bowelnull|Small|LabModifier|false|false||smallnull|Bowel contents|Finding|false|false|C4319010;C0021852;C0021853;C0021853;C4319010;C0021852|bowel contentsnull|Intestines|Anatomy|false|false|C1552853;C0456205;C1546561|bowelnull|contents - HtmlLinkType|Finding|false|false|C4319010;C0021852;C0021853;C4319010;C0021852;C0021853|contents
null|Contents|Finding|false|false|C4319010;C0021852;C0021853;C4319010;C0021852;C0021853|contentsnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Collapsed|Finding|false|false||collapsed
null|Collapse (finding)|Finding|false|false||collapsednull|null|Device|false|false||loopsnull|Together|Modifier|false|false||togethernull|Early|Time|false|false||earlynull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Small|LabModifier|false|false||smallnull|Intestinal Obstruction|Disorder|false|false|C0021853|bowel obstructionnull|Intestines|Anatomy|false|false|C0021843|bowelnull|Obstruction|Finding|false|false||obstructionnull|Changing|Finding|false|false|C0035561|changesnull|Changed status|LabModifier|false|false||changesnull|Table Cell Horizontal Align - right|Finding|false|false|C0035561|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Bone structure of rib|Anatomy|false|false|C0392747;C1552823|ribsnull|Details|Modifier|false|false||detailednull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Abdoman (drug)|Drug|false|false||abdoman
null|Abdoman (drug)|Drug|false|false||abdomannull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvis|Anatomy|false|false|C0153663;C0812455|pelvisnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Small bowel obstruction|Disorder|false|false|C0021853;C4319010;C0021852|small bowel obstructionnull|Abdomen>Small bowel|Anatomy|false|false|C0021843;C0235329;C0028778|small bowel
null|Intestines, Small|Anatomy|false|false|C0021843;C0235329;C0028778|small bowelnull|Small|LabModifier|false|false||smallnull|Intestinal Obstruction|Disorder|false|false|C4319010;C0021852;C0021853|bowel obstructionnull|Intestines|Anatomy|false|false|C0028778;C0235329;C0021843|bowelnull|Obstruction|Finding|false|false|C0021853;C4319010;C0021852|obstructionnull|Transition Mutation|Disorder|false|false||Transitionnull|Transition (action)|Event|false|false||Transitionnull|Point|Modifier|false|false||pointnull|point - UnitsOfMeasure|LabModifier|false|false||pointnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Middle|Modifier|false|false||midnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Evening|Time|false|false||eveningnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Sequence Chromatogram|Finding|false|false|C4266535;C0030797;C0559769|Tracenull|Trace Dosing Unit|LabModifier|false|false||Trace
null|trace amount|LabModifier|false|false||Trace
null|unknown - trace|LabModifier|false|false||Tracenull|effusion|Finding|false|false|C4266535;C0030797;C0559769|free fluidnull|Free of (attribute)|Finding|false|false|C4266535;C0030797;C0559769|freenull|Empty (qualifier)|Modifier|false|false||freenull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false|C4266535;C0030797;C0559769|fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0332148;C0750492;C1883002;C0812455;C0332296;C0205463;C1546638;C0153663;C0013687|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0332148;C0750492;C1883002;C0812455;C0332296;C0205463;C1546638;C0153663;C0013687|pelvis
null|Pelvis|Anatomy|false|false|C0332148;C0750492;C1883002;C0812455;C0332296;C0205463;C1546638;C0153663;C0013687|pelvisnull|Probable diagnosis|Finding|false|false|C4266535;C0030797;C0559769|likely
null|Probably|Finding|false|false|C4266535;C0030797;C0559769|likelynull|Physiological|Finding|false|false|C4266535;C0030797;C0559769|physiologicnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Yellow color|Modifier|false|false||Yellownull|Cloudy|Modifier|false|false||Hazynull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|null|Lab|false|false|C0014792|URINE  RBC
null|Red blood cells urine positive|Lab|false|false|C0014792|URINE  RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792;C0221752;C2188659|RBCnull|null|Attribute|false|false|C0014792|RBCnull|bacteria aspects|Finding|false|false||BACTERIAnull|Bacteria <walking sticks>|Entity|false|false||BACTERIA
null|Bacteria|Entity|false|false||BACTERIAnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||MODnull|Yeast, Dried|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEAST
null|Candida albicans allergenic extract|Drug|false|false||YEASTnull|Saccharomyces cerevisiae|Entity|false|false||YEAST
null|Yeasts|Entity|false|false||YEASTnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|epinephrine|Drug|false|false||EPI
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||EPInull|Exocrine pancreatic insufficiency|Disorder|false|false||EPInull|Eysenck personality inventory|Finding|false|false||EPI
null|TFPI wt Allele|Finding|false|false||EPI
null|TFPI gene|Finding|false|false||EPInull|Electronic Portal Imaging|Procedure|false|false||EPI
null|Echo-Planar Imaging|Procedure|false|false||EPInull|Mucus in urine (finding)|Finding|false|false||URINE  MUCOUSnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mucus (substance)|Finding|false|false||MUCOUS
null|mucus layer|Finding|false|false||MUCOUSnull|Mucous appearance|Modifier|false|false||MUCOUSnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPT
null|SGPT - Glutamate pyruvate transaminase|Drug|false|false||SGPTnull|GPT gene|Finding|false|false||SGPTnull|Serum Alanine Transaminase Test|Procedure|false|false||SGPTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C1415181;C1420113;C5960784;C0201899;C1415181;C4522245;C0004002;C0242192;C1121182|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOT
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||SGOTnull|GOT1 gene|Finding|false|false|C1185650|SGOTnull|Aspartate aminotransferase measurement|Procedure|false|false|C1185650|SGOTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false||LDHnull|Lactate dehydrogenase measurement|Procedure|false|false||LDHnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASE
null|lipase|Drug|false|false||LIPASEnull|Lipase measurement|Procedure|false|false||LIPASEnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Nasogastric tube procedures|Procedure|false|false|C3282907|nasogastric tubenull|Nasogastric tube|Device|false|false||nasogastric tubenull|Nasogastric Route of Administration|Finding|false|false|C3282907|nasogastricnull|Nasogastric|Anatomy|false|false|C0812428;C0694637;C1427122;C1719071|nasogastricnull|Unspecified tube|Finding|false|false|C3282907|tube
null|TUBE1 gene|Finding|false|false|C3282907|tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Polyarteritis Nodosa|Disorder|false|false|C2244316|pannull|ADA2 wt Allele|Finding|false|false|C2244316|pannull|proteasome-activating nucleotidase complex|Anatomy|false|false|C0031036;C5401218|pannull|Pansexuality|Subject|false|false||pannull|Public Affairs Network of Cancer Centers|Entity|false|false||pan
null|Punjabi language|Entity|false|false||pan
null|Pan <Homininae>|Entity|false|false||pannull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|Periodicals|Finding|false|false||serialnull|Serial|Time|false|false||serialnull|physical examination (physical finding)|Finding|false|false||physical examnull|Physical Examination|Procedure|false|false||physical examnull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Nasogastric Route of Administration|Finding|false|false|C3282907|nasogastricnull|Nasogastric|Anatomy|false|false|C0694637|nasogastricnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Day hospital|Device|false|false||hospital daynull|Day hospital|Entity|false|false||hospital daynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Day 2|Finding|false|false||day 2null|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|CT of abdomen|Procedure|false|false|C0230168;C0000726;C0000726|CT of abdomennull|Abdomen|Anatomy|false|false|C0941288;C0153662;C0412620|abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726;C0000726|abdomennull|Abdomen problem|Finding|false|false|C0000726;C0230168;C0000726|abdomennull|Abdominal Cavity|Anatomy|false|false|C0153662;C0412620;C0941288|abdomen
null|Abdomen|Anatomy|false|false|C0153662;C0412620;C0941288|abdomennull|Malignant neoplasm of pelvis|Disorder|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis problem|Finding|false|false|C4266535;C0030797;C0559769|pelvisnull|Pelvis+|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvic cavity structure|Anatomy|false|false|C0153663;C0812455|pelvis
null|Pelvis|Anatomy|false|false|C0153663;C0812455|pelvisnull|Increase|Finding|false|false||increasenull|Academic degree|Finding|false|false||degreenull|Levels (qualifier value)|Modifier|false|false||degreenull|Degree Unit of Plane Angle|LabModifier|false|false||degree
null|Degree or extent|LabModifier|false|false||degreenull|Obstruction|Finding|false|false||obstructionnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|NPO - Nothing by mouth|Procedure|false|false||NPOnull|null|Entity|false|false||NPOnull|Nasogastric Route of Administration|Finding|false|false|C3282907|nasogastricnull|Nasogastric|Anatomy|false|false|C0694637|nasogastricnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Initially|Time|false|false||initiallynull|morphine|Drug|false|false|C0149576|morphine
null|morphine|Drug|false|false|C0149576|morphinenull|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|p-Chloroamphetamine|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCA
null|pyrrolidonecarboxylic acid|Drug|false|false|C0149576|PCAnull|Posterior cortical atrophy syndrome|Disorder|false|false|C0149576|PCA
null|Familial lichen amyloidosis|Disorder|false|false|C0149576|PCAnull|PCA Message Structure|Finding|false|false|C0149576|PCA
null|CHOANAL ATRESIA, POSTERIOR|Finding|false|false|C0149576|PCA
null|FLVCR1 gene|Finding|false|false|C0149576|PCAnull|Patient controlled intravenous analgesia|Procedure|false|false|C0149576|PCA
null|Passive Cutaneous Anaphylaxis|Procedure|false|false|C0149576|PCA
null|Patient-Controlled Analgesia|Procedure|false|false|C0149576|PCAnull|Structure of posterior cerebral artery|Anatomy|false|false|C0812428;C1427122;C1719071;C0220723;C1836722;C1549860;C0268398;C4275079;C0026549;C0078944;C5968782;C0030625;C0034330;C0030131|PCAnull|Principal Component Analysis|LabModifier|false|false||PCAnull|Nasogastric tube procedures|Procedure|false|false|C0149576;C3282907|nasogastric tubenull|Nasogastric tube|Device|false|false||nasogastric tubenull|Nasogastric Route of Administration|Finding|false|false|C3282907|nasogastricnull|Nasogastric|Anatomy|false|false|C1427122;C1719071;C0694637;C0812428|nasogastricnull|Unspecified tube|Finding|false|false|C3282907;C0149576|tube
null|TUBE1 gene|Finding|false|false|C3282907;C0149576|tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Clear liquid diet|Procedure|false|false||clear liquid dietnull|Clear liquid|Finding|false|false||clear liquidnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Liquid diet|Procedure|false|false||liquid dietnull|Liquid Dosage Form|Drug|false|false||liquid
null|Liquid substance|Drug|false|false||liquidnull|Liquid (finding)|Finding|false|false||liquidnull|Liquid diet|Procedure|false|false||liquidnull|Liquid (state of matter)|Modifier|false|false||liquidnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Hour|Time|false|false||hoursnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Defecation|Finding|false|false|C0021853|bowel movementsnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementsnull|Oral pain|Finding|false|false|C0226896|oral painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1549543;C0030193;C1527415;C4521986;C0221776;C3244316;C4284232|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false|C0226896|pain
null|Pain|Finding|false|false|C0226896|painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false|C0226896|medication
null|Medications|Finding|false|false|C0226896|medicationnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803;C5575035;C1554187|incisionnull|Well (answer to question)|Finding|false|false|C2338258|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Staple, Surgical|Device|false|false||staplesnull|Gender Status - Intact|Finding|false|false|C2338258|intactnull|Intact|Modifier|false|false||intactnull|Uncomplicated|Modifier|false|false||uncomplicatednull|Course|Time|false|false||coursenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MAJOR AFFECTIVE DISORDER 2|Disorder|false|false||MDInull|Myositis Damage Index|Finding|false|false||MDInull|Metered Dose Inhaler|Device|false|false||MDInull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Wheezing|Finding|false|false||wheezesnull|Flovent|Drug|false|false||Flovent
null|Flovent|Drug|false|false||Floventnull|Inhaler (unit of presentation)|Finding|false|false||inhalernull|Inhaler|Device|false|false||inhalernull|Inhaler Dosing Unit|LabModifier|false|false||inhalernull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Wheezing|Finding|false|false||wheezesnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||dailynull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|albuterol sulfate|Drug|false|false||Albuterol Sulfate
null|albuterol sulfate|Drug|false|false||Albuterol Sulfatenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|Inhalers, Aerosol|Device|false|false||Aerosol Inhalernull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Every six hours|Time|false|false||Q6Hnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Wheezing|Finding|false|false||wheezingnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Puff Dosing Unit|LabModifier|false|false||Puff
null|Picofarad|LabModifier|false|false||Puffnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false||2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Every four hours|Time|false|false||Q4Hnull|4 Hours|Time|false|false||4 hoursnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1332410;C4546282|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1332410;C4546282|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C0524463;C1325531|BIDnull|BID gene|Finding|false|false|C0524463;C1325531|BIDnull|Twice a day|Time|false|false||BIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|trazodone|Drug|false|false||Trazodone
null|trazodone|Drug|false|false||Trazodonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Wellbutrin|Drug|false|false||Wellbutrin
null|Wellbutrin|Drug|false|false||Wellbutrinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Enneking High Surgical Grade|Finding|false|false|C4319010;C0021852|High grade
null|Severe (severity modifier)|Finding|false|false|C4319010;C0021852|High gradenull|Message Waiting Priority - High|Finding|false|false||High
null|high - ActExposureLevelCode|Finding|false|false||High
null|IPSS Risk Category High|Finding|false|false||High
null|IPSS-R Risk Category High|Finding|false|false||High
null|High (finding)|Finding|false|false||Highnull|Observation Value - High|Modifier|false|false||High
null|High|Modifier|false|false||High
null|Abnormally high|Modifier|false|false||Highnull|Histopathologic Grade|Finding|false|false|C4319010;C0021852|grade
null|Grade|Finding|false|false|C4319010;C0021852|grade
null|School Grade|Finding|false|false|C4319010;C0021852|gradenull|Small bowel obstruction|Disorder|false|false|C4319010;C0021852;C0021853|small bowel obstructionnull|Abdomen>Small bowel|Anatomy|false|false|C4554016;C0205082;C0235329;C0919553;C3244287;C0441800|small bowel
null|Intestines, Small|Anatomy|false|false|C4554016;C0205082;C0235329;C0919553;C3244287;C0441800|small bowelnull|Small|LabModifier|false|false||smallnull|Intestinal Obstruction|Disorder|false|false|C0021853|bowel obstructionnull|Intestines|Anatomy|false|false|C0021843;C0235329|bowelnull|Obstruction|Finding|false|false||obstructionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Intestines|Anatomy|false|false||bowelnull|Movement|Finding|false|false||movementsnull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Nurse Practitioner - Procedure Practitioner Identifier Code Type|Finding|false|false||nurse practitioner
null|nurse practitioner Degree/license/certificate|Finding|false|false||nurse practitionernull|nurse practitioner|Subject|false|false||nurse practitionernull|Nurses|Subject|false|false||nursenull|Practitioner|Subject|false|false||practitionernull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||return tonull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Accident and Emergency department|Device|false|false||Emergency Departmentnull|interventional services emergency department|Entity|false|false||Emergency Department
null|Accident and Emergency department|Entity|false|false||Emergency Departmentnull|Level of Care - Emergency|Finding|false|false||Emergency
null|Consent Non-Disclosure Reason - Emergency|Finding|false|false||Emergency
null|Admission Type - Emergency|Finding|false|false||Emergency
null|Referral category - Emergency|Finding|false|false||Emergency
null|Emergencies [Disease/Finding]|Finding|false|false||Emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||Emergency
null|Certification patient type - Emergency|Finding|false|false||Emergency
null|Encounter Admission Source - emergency|Finding|false|false||Emergency
null|Patient Class - Emergency|Finding|false|false||Emergency
null|Visit Priority Code - Emergency|Finding|false|false||Emergencynull|emergency encounter|Procedure|false|false||Emergencynull|Emergency Situation|Phenomenon|false|false||Emergencynull|Specialty Type - Emergency|Title|false|false||Emergencynull|Bale out|Time|false|false||Emergencynull|Department - No suggested values defined|Finding|false|false||Department
null|Organization Unit Type - Department|Finding|false|false||Department
null|Department - Charge type|Finding|false|false||Departmentnull|Department|Entity|false|false||Departmentnull|Patient location type - Department|Modifier|false|false||Department
null|Department - Person location type|Modifier|false|false||Departmentnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Tightness sensation quality|Modifier|false|false||tightnessnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Wheezing|Finding|false|false||wheezenull|Vomiting|Finding|false|false||vomitingnull|Liquid substance|Drug|true|false||fluidsnull|Mouse Body Fluid or Substance|Finding|true|false||fluidsnull|Fluid Therapy|Procedure|true|false||fluidsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Dehydration|Disorder|false|false||dehydratednull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Indication of (contextual qualifier)|Finding|false|false||reasonsnull|Signs of dehydration|Finding|false|false||Signs of dehydrationnull|Aspects of signs|Finding|false|false|C0230028;C0226896|Signs
null|Physical findings|Finding|false|false|C0230028;C0226896|Signsnull|Manufactured sign|Device|false|false||Signsnull|dehydration (Na, H2O)|Disorder|false|false|C0230028;C0226896|dehydration
null|Dehydration|Disorder|false|false|C0230028;C0226896|dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|Xerostomia|Disorder|false|false|C0230028;C0226896|dry mouthnull|Oral cavity|Anatomy|false|false|C2062903;C0011175;C0220912;C0311392;C0043352|mouth
null|Oral region|Anatomy|false|false|C2062903;C0011175;C0220912;C0311392;C0043352|mouthnull|Rapid|Modifier|false|false||rapidnull|Heart beat|Finding|false|false||heartbeatnull|Pulse Rate|Attribute|false|false||heartbeatnull|feeling dizzy|Finding|false|false||feeling dizzynull|Feelings|Finding|false|false||feelingnull|Dizziness|Finding|false|false||dizzynull|Faint - appearance|Finding|false|false||faint
null|Syncope|Finding|false|false||faintnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Dark color|Modifier|false|false||darknull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Materials|Drug|false|false||materialnull|Defecation|Finding|false|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|false|false||movementnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hour|Time|false|false||hoursnull|Within 24 hours|Time|false|false||within 24 hoursnull|24 Hours|Time|false|false||24 hoursnull|Hour|Time|false|false||hoursnull|Call - dosing instruction fragment|Finding|false|false||Call
null|Call (Instruction)|Finding|false|false||Call
null|Decision|Finding|false|false||Call
null|CHL1 gene|Finding|false|false||Callnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Stat (do immediately)|Time|false|false||immediatelynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Changing|Finding|false|false|C1515974|changesnull|Changed status|LabModifier|false|false||changesnull|Transaction counts and value totals - location|Finding|false|false|C1515974|locationnull|Anatomic Site|Anatomy|false|false|C1555588;C0392747|locationnull|location participation type|Device|false|false||locationnull|location participation type|Entity|false|false||locationnull|Location|Modifier|false|false||locationnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Chills|Finding|false|false||chillsnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Degrees fahrenheit|LabModifier|false|false||Fahrenheitnull|degrees Celsius|LabModifier|false|false||degrees Celsiusnull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|degrees Celsius|LabModifier|false|false||Celsius
null|Celsius Scale|LabModifier|false|false||Celsiusnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Concern|Finding|false|false||concernnull|Regular|Modifier|false|false||regularnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Take|Procedure|false|false||takenull|New medications|Drug|false|false||new medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Several|LabModifier|false|false||severalnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Quantity|LabModifier|false|false||amountsnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Lifting|Event|false|false||liftingnull|Weights - exercise activity|Finding|false|false||weightsnull|Weight|LabModifier|false|false||weightsnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Automobile Driving|Finding|false|false||drivingnull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Incision care|Procedure|false|false|C2338258|Incision Carenull|Surgical wound|Disorder|false|false|C2338258|Incisionnull|Surgical incisions|Procedure|false|false|C2338258|Incisionnull|Cranial incision point|Anatomy|false|false|C1947933;C0580931;C2362566;C0150258;C0332803;C0184898|Incisionnull|In care (finding)|Finding|false|false|C2338258|Care
null|Continuity Assessment Record and Evaluation|Finding|false|false|C2338258|Carenull|care activity|Event|false|false|C2338258|Carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Nurse Practitioner - Procedure Practitioner Identifier Code Type|Finding|false|false||nurse practitioner
null|nurse practitioner Degree/license/certificate|Finding|false|false||nurse practitionernull|nurse practitioner|Subject|false|false||nurse practitionernull|Nurses|Subject|false|false||nursenull|Practitioner|Subject|false|false||practitionernull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false|C2338258|drainage
null|Body Fluid Discharge|Finding|false|false|C2338258|drainagenull|Drainage procedure|Procedure|false|false|C2338258|drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0012621;C2926602;C0184898;C0013103|incisionnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Surgical wound|Disorder|false|false||surgical incisionsnull|Surgical incisions|Procedure|false|false||surgical incisionsnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Surgical incisions|Procedure|false|false||incisionsnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Soap Dosage Form|Drug|false|false||soapnull|Soap|Device|false|false||soapnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Gently|Modifier|false|false||Gentlynull|Fenamole|Drug|false|false||pat
null|Fenamole|Drug|false|false||patnull|Paroxysmal atrial tachycardia|Disorder|false|false||patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||pat
null|protein acetyltransferase activity|Finding|false|false||patnull|Thermoacoustic Computed Tomography|Procedure|false|false||patnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Staple, Surgical|Device|false|false||staplesnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Steri-Strip|Device|false|false||steri-stripsnull|Silene|Entity|false|false||sterinull|strip medical device|Device|false|false||stripsnull|Own|Finding|false|false||ownnull|strip medical device|Device|false|false||stripsnull|day|Time|false|false||daysnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C1561538;C1561539|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Transaction counts and value totals - day|Finding|false|false|C1515974|day
null|Precision - day|Finding|false|false|C1515974|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Odors|Phenomenon|false|false||odornull|Yellow color|Modifier|false|false||yellownull|Bloody|Finding|false|false||bloodynull|Hemorrhagic|Modifier|false|false||bloodynull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions