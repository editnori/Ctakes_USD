 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
NEUROLOGY|156,165
<EOL>|165,166
<EOL>|167,168
amoxicillin|180,191
<EOL>|191,192
<EOL>|193,194
Attending|194,203
:|203,204
_|205,206
_|206,207
_|207,208
.|208,209
<EOL>|209,210
<EOL>|211,212
Weakness|229,237
and|238,241
lethargy|242,250
<EOL>|251,252
<EOL>|253,254
Major|254,259
Surgical|260,268
or|269,271
Invasive|272,280
Procedure|281,290
:|290,291
<EOL>|291,292
None|292,296
<EOL>|296,297
<EOL>|297,298
<EOL>|299,300
Patient|328,335
is|336,338
a|339,340
_|341,342
_|342,343
_|343,344
year|345,349
old|350,353
female|354,360
with|361,365
history|366,373
of|374,376
chronic|377,384
<EOL>|384,385
abdominal|385,394
pain|395,399
and|400,403
anemia|404,410
w|411,412
/|412,413
recent|414,420
Fe|421,423
sucrose|424,431
infusion|432,440
(|441,442
_|442,443
_|443,444
_|444,445
)|445,446
<EOL>|446,447
complicated|447,458
by|459,461
infusion|462,470
reaction|471,479
(|480,481
mottling|481,489
and|490,493
discoloration|494,507
of|508,510
<EOL>|510,511
feet|511,515
)|515,516
s|517,518
/|518,519
p|519,520
IV|521,523
steroids|524,532
who|533,536
presents|537,545
with|546,550
increasing|551,561
lethargy|562,570
and|571,574
<EOL>|574,575
headache|575,583
.|583,584
<EOL>|584,585
<EOL>|585,586
History|586,593
per|594,597
_|598,599
_|599,600
_|600,601
records|602,609
and|610,613
per|614,617
her|618,621
Aunt|622,626
as|627,629
patient|630,637
can|638,641
not|641,644
<EOL>|644,645
provide|645,652
much|653,657
history|658,665
.|665,666
Per|667,670
her|671,674
aunt|675,679
,|679,680
_|681,682
_|682,683
_|683,684
has|685,688
been|689,693
doing|694,699
well|700,704
<EOL>|704,705
recently|705,713
without|714,721
any|722,725
illness|726,733
,|733,734
behavioral|735,745
change|746,752
.|752,753
She|754,757
had|758,761
a|762,763
cold|764,768
<EOL>|768,769
she|769,772
was|773,776
getting|777,784
over|785,789
but|790,793
otherwise|794,803
doing|804,809
well|810,814
.|814,815
She|816,819
had|820,823
an|824,826
Fe|827,829
<EOL>|829,830
transfusion|830,841
on|842,844
_|845,846
_|846,847
_|847,848
around|849,855
3|856,857
:|857,858
30P|858,861
at|862,864
_|865,866
_|866,867
_|867,868
and|869,872
the|873,876
aunt|877,881
<EOL>|881,882
accompanied|882,893
her|894,897
to|898,900
the|901,904
visit|905,910
.|910,911
Towards|912,919
the|920,923
end|924,927
of|928,930
the|931,934
infusion|935,943
,|943,944
<EOL>|944,945
_|945,946
_|946,947
_|947,948
developed|949,958
mottle|959,965
purple|966,972
lower|973,978
extremities|979,990
and|991,994
was|995,998
having|999,1005
<EOL>|1005,1006
nausea|1006,1012
,|1012,1013
heart|1014,1019
racing|1020,1026
.|1026,1027
She|1028,1031
was|1032,1035
sent|1036,1040
to|1041,1043
_|1044,1045
_|1045,1046
_|1046,1047
where|1048,1053
she|1054,1057
had|1058,1061
SBP|1062,1065
<EOL>|1065,1066
up|1066,1068
to|1069,1071
144|1072,1075
.|1075,1076
Her|1077,1080
exam|1081,1085
per|1086,1089
_|1090,1091
_|1091,1092
_|1092,1093
records|1094,1101
notable|1102,1109
for|1110,1113
"|1114,1115
shivering|1115,1124
...|1124,1127
<EOL>|1127,1128
does|1128,1132
n't|1132,1135
open|1136,1140
her|1141,1144
eyes|1145,1149
...|1149,1152
mottled|1152,1159
hands|1160,1165
and|1166,1169
feet|1170,1174
"|1174,1175
.|1175,1176
There|1177,1182
was|1183,1186
no|1187,1189
<EOL>|1189,1190
concern|1190,1197
for|1198,1201
respiratory|1202,1213
distress|1214,1222
.|1222,1223
She|1224,1227
was|1228,1231
given|1232,1237
50|1238,1240
mg|1241,1243
IV|1244,1246
<EOL>|1246,1247
Benadryl|1247,1255
,|1255,1256
100|1257,1260
mg|1261,1263
IV|1264,1266
hydrocortisone|1267,1281
and|1282,1285
observed|1286,1294
for|1295,1298
5|1299,1300
hours|1301,1306
and|1307,1310
<EOL>|1310,1311
then|1311,1315
discharged|1316,1326
.|1326,1327
At|1328,1330
that|1331,1335
time|1336,1340
_|1341,1342
_|1342,1343
_|1343,1344
was|1345,1348
reportedly|1349,1359
"|1360,1361
lethargic|1361,1370
"|1370,1371
<EOL>|1371,1372
meaning|1372,1379
sleeping|1380,1388
frequently|1389,1399
but|1400,1403
able|1404,1408
to|1409,1411
sit|1412,1415
up|1416,1418
and|1419,1422
walk|1423,1427
without|1428,1435
<EOL>|1435,1436
issue|1436,1441
.|1441,1442
They|1443,1447
arrived|1448,1455
home|1456,1460
and|1461,1464
_|1465,1466
_|1466,1467
_|1467,1468
went|1469,1473
to|1474,1476
bed|1477,1480
.|1480,1481
Around|1482,1488
6|1489,1490
:|1490,1491
00|1491,1493
AM|1494,1496
<EOL>|1496,1497
on|1497,1499
_|1500,1501
_|1501,1502
_|1502,1503
,|1503,1504
_|1505,1506
_|1506,1507
_|1507,1508
aunt|1509,1513
check|1514,1519
on|1520,1522
her|1523,1526
and|1527,1530
she|1531,1534
was|1535,1538
still|1539,1544
sleeping|1545,1553
.|1553,1554
<EOL>|1554,1555
She|1555,1558
was|1559,1562
reporting|1563,1572
a|1573,1574
headache|1575,1583
(|1584,1585
which|1585,1590
the|1591,1594
transfusion|1595,1606
place|1607,1612
said|1613,1617
<EOL>|1617,1618
would|1618,1623
happen|1624,1630
)|1630,1631
but|1632,1635
did|1636,1639
not|1640,1643
mention|1644,1651
other|1652,1657
characteristic|1658,1672
.|1672,1673
<EOL>|1674,1675
_|1675,1676
_|1676,1677
_|1677,1678
<EOL>|1678,1679
aunt|1679,1683
gave|1684,1688
her|1689,1692
acetaminophen|1693,1706
and|1707,1710
water|1711,1716
and|1717,1720
_|1721,1722
_|1722,1723
_|1723,1724
went|1725,1729
back|1730,1734
to|1735,1737
<EOL>|1737,1738
sleep|1738,1743
.|1743,1744
Over|1745,1749
the|1750,1753
next|1754,1758
few|1759,1762
hours|1763,1768
,|1768,1769
she|1770,1773
heard|1774,1779
_|1780,1781
_|1781,1782
_|1782,1783
awake|1784,1789
several|1790,1797
<EOL>|1797,1798
times|1798,1803
and|1804,1807
use|1808,1811
the|1812,1815
bathroom|1816,1824
.|1824,1825
Then|1826,1830
as|1831,1833
it|1834,1836
got|1837,1840
later|1841,1846
and|1847,1850
later|1851,1856
into|1857,1861
<EOL>|1861,1862
the|1862,1865
day|1866,1869
and|1870,1873
_|1874,1875
_|1875,1876
_|1876,1877
was|1878,1881
not|1882,1885
up|1886,1888
and|1889,1892
about|1893,1898
yet|1899,1902
,|1902,1903
her|1904,1907
aunt|1908,1912
became|1913,1919
<EOL>|1919,1920
worried|1920,1927
.|1927,1928
She|1929,1932
told|1933,1937
_|1938,1939
_|1939,1940
_|1940,1941
to|1942,1944
call|1945,1949
the|1950,1953
_|1954,1955
_|1955,1956
_|1956,1957
which|1958,1963
she|1964,1967
<EOL>|1967,1968
was|1968,1971
able|1972,1976
to|1977,1979
do|1980,1982
.|1982,1983
She|1984,1987
reportedly|1988,1998
said|1999,2003
she|2004,2007
continued|2008,2017
to|2018,2020
have|2021,2025
a|2026,2027
<EOL>|2027,2028
headache|2028,2036
and|2037,2040
felt|2041,2045
sleepy|2046,2052
.|2052,2053
She|2054,2057
was|2058,2061
instructed|2062,2072
to|2073,2075
go|2076,2078
to|2079,2081
the|2082,2085
ED|2086,2088
.|2088,2089
<EOL>|2090,2091
<EOL>|2091,2092
She|2092,2095
went|2096,2100
to|2101,2103
the|2104,2107
ED|2108,2110
at|2111,2113
_|2114,2115
_|2115,2116
_|2116,2117
for|2118,2121
evaluation|2122,2132
.|2132,2133
At|2134,2136
_|2137,2138
_|2138,2139
_|2139,2140
she|2141,2144
<EOL>|2144,2145
had|2145,2148
T|2149,2150
99.5|2151,2155
,|2155,2156
P|2157,2158
58|2159,2161
,|2161,2162
RR|2163,2165
15|2166,2168
and|2169,2172
sat|2173,2176
100|2177,2180
%|2180,2181
.|2181,2182
BP|2183,2185
110|2186,2189
/|2189,2190
67|2190,2192
.|2192,2193
She|2194,2197
was|2198,2201
<EOL>|2201,2202
reportedly|2202,2212
drowsy|2213,2219
and|2220,2223
arousing|2224,2232
to|2233,2235
voice|2236,2241
,|2241,2242
"|2243,2244
alert|2244,2249
oriented|2250,2258
x3|2259,2261
"|2261,2262
,|2262,2263
<EOL>|2263,2264
consistent|2264,2274
eye|2275,2278
fluttering|2279,2289
,|2289,2290
pupils|2291,2297
reactive|2298,2306
to|2307,2309
light|2310,2315
and|2316,2319
<EOL>|2319,2320
extraocular|2320,2331
eye|2332,2335
movements|2336,2345
full|2346,2350
,|2350,2351
with|2352,2356
reportedly|2357,2367
"|2368,2369
non|2369,2372
focal|2373,2378
<EOL>|2379,2380
exam|2380,2384
"|2384,2385
.|2385,2386
<EOL>|2386,2387
Lab|2387,2390
work|2391,2395
notable|2396,2403
for|2404,2407
WBC|2408,2411
7.2|2412,2415
,|2415,2416
Hgb|2417,2420
13.2|2421,2425
,|2425,2426
Na|2427,2429
142|2430,2433
,|2433,2434
bicarb|2435,2441
26|2442,2444
,|2444,2445
Cr|2446,2448
<EOL>|2448,2449
0.9|2449,2452
,|2452,2453
Ca|2454,2456
9.4|2457,2460
,|2460,2461
normal|2462,2468
LFTs|2469,2473
,|2473,2474
Fe|2475,2477
360|2478,2481
,|2481,2482
Ferritin|2483,2491
438.|2492,2496
VBG|2497,2500
pH|2501,2503
was|2504,2507
7.43|2508,2512
,|2512,2513
<EOL>|2513,2514
PCO2|2514,2518
was|2519,2522
45.|2523,2526
She|2526,2529
had|2530,2533
a|2534,2535
normal|2536,2542
_|2543,2544
_|2544,2545
_|2545,2546
and|2547,2550
LP|2551,2553
with|2554,2558
WBC|2559,2562
2|2563,2564
,|2564,2565
100|2566,2569
%|2569,2570
<EOL>|2570,2571
monocytes|2571,2580
glucose|2581,2588
57|2589,2591
,|2591,2592
protein|2593,2600
24|2601,2603
,|2603,2604
no|2605,2607
xanthochromia|2608,2621
.|2621,2622
She|2623,2626
<EOL>|2626,2627
ultimately|2627,2637
had|2638,2641
MRA|2642,2645
and|2646,2649
MRV|2650,2653
which|2654,2659
showed|2660,2666
no|2667,2669
thrombus|2670,2678
or|2679,2681
venoous|2682,2689
<EOL>|2689,2690
thrombosis|2690,2700
.|2700,2701
She|2702,2705
was|2706,2709
transferred|2710,2721
to|2722,2724
_|2725,2726
_|2726,2727
_|2727,2728
for|2729,2732
further|2733,2740
management|2741,2751
.|2751,2752
<EOL>|2752,2753
<EOL>|2753,2754
On|2754,2756
my|2757,2759
interview|2760,2769
she|2770,2773
can|2774,2777
not|2777,2780
provide|2781,2788
much|2789,2793
history|2794,2801
other|2802,2807
than|2808,2812
to|2813,2815
<EOL>|2816,2817
say|2817,2820
<EOL>|2820,2821
she|2821,2824
is|2825,2827
here|2828,2832
because|2833,2840
"|2841,2842
I|2842,2843
'|2843,2844
m|2844,2845
tired|2846,2851
"|2851,2852
.|2852,2853
She|2854,2857
keeps|2858,2863
her|2864,2867
eyes|2868,2872
closed|2873,2879
<EOL>|2880,2881
during|2881,2887
<EOL>|2887,2888
questioning|2888,2899
.|2899,2900
She|2901,2904
reports|2905,2912
headache|2913,2921
but|2922,2925
can|2926,2929
not|2929,2932
describe|2933,2941
where|2942,2947
it|2948,2950
<EOL>|2951,2952
is|2952,2954
<EOL>|2954,2955
or|2955,2957
features|2958,2966
other|2967,2972
than|2973,2977
+|2978,2979
photophobia|2979,2990
.|2990,2991
She|2992,2995
is|2996,2998
unable|2999,3005
to|3006,3008
<EOL>|3009,3010
participate|3010,3021
<EOL>|3021,3022
in|3022,3024
other|3025,3030
questioning|3031,3042
,|3042,3043
often|3044,3049
getting|3050,3057
tearful|3058,3065
and|3066,3069
saying|3070,3076
"|3077,3078
the|3078,3081
<EOL>|3081,3082
questions|3082,3091
are|3092,3095
hard|3096,3100
"|3100,3101
.|3101,3102
<EOL>|3103,3104
<EOL>|3104,3105
Per|3105,3108
her|3109,3112
father|3113,3119
and|3120,3123
aunt|3124,3128
,|3128,3129
she|3130,3133
has|3134,3137
no|3138,3140
history|3141,3148
of|3149,3151
seizures|3152,3160
,|3160,3161
or|3162,3164
CNS|3165,3168
<EOL>|3168,3169
infection|3169,3178
.|3178,3179
She|3180,3183
did|3184,3187
have|3188,3192
a|3193,3194
concussion|3195,3205
at|3206,3208
_|3209,3210
_|3210,3211
_|3211,3212
years|3213,3218
old|3219,3222
.|3222,3223
<EOL>|3224,3225
<EOL>|3226,3227
Anemia|3249,3255
<EOL>|3256,3257
<EOL>|3258,3259
:|3273,3274
<EOL>|3274,3275
_|3275,3276
_|3276,3277
_|3277,3278
<EOL>|3278,3279
:|3293,3294
<EOL>|3294,3295
Mother|3295,3301
with|3302,3306
a|3307,3308
celiac|3309,3315
disease|3316,3323
and|3324,3327
autoimmune|3328,3338
hypothyroidism|3339,3353
.|3353,3354
Dad|3355,3358
<EOL>|3358,3359
is|3359,3361
healthy|3362,3369
.|3369,3370
She|3371,3374
has|3375,3378
a|3379,3380
cousin|3381,3387
with|3388,3392
seizures|3393,3401
.|3401,3402
<EOL>|3402,3403
<EOL>|3404,3405
Admission|3420,3429
exam|3430,3434
:|3434,3435
<EOL>|3435,3436
98.1|3436,3440
76|3441,3443
130|3444,3447
/|3447,3448
78|3448,3450
14|3451,3453
96|3454,3456
%|3456,3457
RA|3458,3460
<EOL>|3461,3462
General|3462,3469
:|3469,3470
appears|3471,3478
to|3479,3481
be|3482,3484
sleeping|3485,3493
,|3493,3494
occasional|3495,3505
eye|3506,3509
lid|3510,3513
fluttering|3514,3524
,|3524,3525
<EOL>|3525,3526
lip|3526,3529
movements|3530,3539
,|3539,3540
occasional|3541,3551
slow|3552,3556
movements|3557,3566
of|3567,3569
head|3570,3574
from|3575,3579
side|3580,3584
to|3585,3587
<EOL>|3587,3588
side|3588,3592
<EOL>|3592,3593
HEENT|3593,3598
:|3598,3599
no|3600,3602
trauma|3603,3609
,|3609,3610
no|3611,3613
jaundice|3614,3622
,|3622,3623
no|3624,3626
lesions|3627,3634
of|3635,3637
oropharynx|3638,3648
<EOL>|3649,3650
CV|3650,3652
:|3652,3653
RRR|3654,3657
,|3657,3658
wwp|3659,3662
<EOL>|3662,3663
Pulm|3663,3667
:|3667,3668
breathing|3669,3678
comfortably|3679,3690
on|3691,3693
RA|3694,3696
<EOL>|3697,3698
Ext|3698,3701
:|3701,3702
clammy|3703,3709
,|3709,3710
warm|3711,3715
and|3716,3719
no|3720,3722
rash|3723,3727
<EOL>|3727,3728
<EOL>|3728,3729
Neurologic|3729,3739
:|3739,3740
<EOL>|3740,3741
<EOL>|3741,3742
-|3742,3743
Mental|3743,3749
Status|3750,3756
:|3756,3757
She|3758,3761
frequently|3762,3772
gets|3773,3777
upset|3778,3783
during|3784,3790
exam|3791,3795
and|3796,3799
is|3800,3802
<EOL>|3802,3803
tearful|3803,3810
at|3811,3813
times|3814,3819
,|3819,3820
then|3821,3825
abulic|3826,3832
at|3833,3835
other|3836,3841
times|3842,3847
.|3847,3848
Eyes|3849,3853
open|3854,3858
only|3859,3863
<EOL>|3863,3864
briefly|3864,3871
to|3872,3874
voice|3875,3880
.|3880,3881
She|3882,3885
is|3886,3888
oriented|3889,3897
to|3898,3900
_|3901,3902
_|3902,3903
_|3903,3904
but|3905,3908
not|3909,3912
full|3913,3917
<EOL>|3917,3918
date|3918,3922
.|3922,3923
Knows|3924,3929
she|3930,3933
is|3934,3936
in|3937,3939
a|3940,3941
"|3942,3943
hospital|3943,3951
"|3951,3952
but|3953,3956
not|3957,3960
the|3961,3964
name|3965,3969
.|3969,3970
She|3971,3974
says|3975,3979
<EOL>|3980,3981
she|3981,3984
<EOL>|3984,3985
is|3985,3987
in|3988,3990
the|3991,3994
hospital|3995,4003
because|4004,4011
,|4011,4012
"|4013,4014
I|4014,4015
'|4015,4016
m|4016,4017
tired|4018,4023
"|4023,4024
.|4024,4025
She|4026,4029
is|4030,4032
unable|4033,4039
to|4040,4042
<EOL>|4043,4044
provide|4044,4051
<EOL>|4051,4052
history|4052,4059
.|4059,4060
Speech|4061,4067
is|4068,4070
not|4071,4074
dysarthric|4075,4085
,|4085,4086
says|4087,4091
_|4092,4093
_|4093,4094
_|4094,4095
words|4096,4101
when|4102,4106
asked|4107,4112
<EOL>|4112,4113
questions|4113,4122
,|4122,4123
no|4124,4126
spontaneous|4127,4138
speech|4139,4145
output|4146,4152
.|4152,4153
Follows|4154,4161
simple|4162,4168
commands|4169,4177
<EOL>|4177,4178
like|4178,4182
open|4183,4187
eyes|4188,4192
,|4192,4193
lift|4194,4198
legs|4199,4203
.|4203,4204
She|4205,4208
is|4209,4211
able|4212,4216
to|4217,4219
name|4220,4224
"|4225,4226
key|4226,4229
"|4229,4230
and|4231,4234
<EOL>|4234,4235
"|4235,4236
feather|4236,4243
"|4243,4244
on|4245,4247
stroke|4248,4254
card|4255,4259
but|4260,4263
then|4264,4268
stops|4269,4274
naming|4275,4281
and|4282,4285
closes|4286,4292
her|4293,4296
<EOL>|4296,4297
eyes|4297,4301
.|4301,4302
She|4303,4306
reads|4307,4312
the|4313,4316
first|4317,4322
sentence|4323,4331
on|4332,4334
stroke|4335,4341
card|4342,4346
but|4347,4350
then|4351,4355
no|4356,4358
<EOL>|4358,4359
more|4359,4363
and|4364,4367
closes|4368,4374
her|4375,4378
eyes|4379,4383
.|4383,4384
When|4385,4389
asked|4390,4395
to|4396,4398
describe|4399,4407
stroke|4408,4414
card|4415,4419
<EOL>|4419,4420
picture|4420,4427
she|4428,4431
says|4432,4436
,|4436,4437
"|4438,4439
dishes|4439,4445
"|4445,4446
.|4446,4447
She|4448,4451
does|4452,4456
not|4457,4460
participate|4461,4472
in|4473,4475
further|4476,4483
<EOL>|4483,4484
exam|4484,4488
.|4488,4489
<EOL>|4489,4490
<EOL>|4490,4491
-|4491,4492
Cranial|4492,4499
Nerves|4500,4506
:|4506,4507
<EOL>|4507,4508
II|4509,4511
,|4511,4512
III|4513,4516
,|4516,4517
IV|4518,4520
,|4520,4521
VI|4522,4524
:|4524,4525
Pupils|4527,4533
8|4534,4535
mm|4536,4538
-|4538,4539
>|4539,4540
6|4540,4541
mm|4542,4544
.|4544,4545
EOMI|4546,4550
without|4551,4558
nystagmus|4559,4568
.|4568,4569
<EOL>|4570,4571
VFF|4571,4574
<EOL>|4574,4575
to|4575,4577
confrontation|4578,4591
.|4591,4592
Fundoscopic|4594,4605
exam|4606,4610
revealed|4611,4619
no|4620,4622
papilledema|4623,4634
,|4634,4635
<EOL>|4635,4636
exudates|4636,4644
,|4644,4645
or|4646,4648
hemorrhages|4649,4660
.|4660,4661
<EOL>|4661,4662
VII|4663,4666
:|4666,4667
No|4668,4670
facial|4671,4677
droop|4678,4683
,|4683,4684
facial|4685,4691
musculature|4692,4703
symmetric|4704,4713
with|4714,4718
<EOL>|4719,4720
grimace|4720,4727
.|4727,4728
<EOL>|4728,4729
VIII|4730,4734
:|4734,4735
Hearing|4736,4743
intact|4744,4750
to|4751,4753
exam|4754,4758
<EOL>|4758,4759
IX|4760,4762
,|4762,4763
X|4764,4765
:|4765,4766
Palate|4767,4773
elevates|4774,4782
symmetrically|4783,4796
.|4796,4797
<EOL>|4797,4798
XII|4799,4802
:|4802,4803
Tongue|4804,4810
protrudes|4811,4820
in|4821,4823
midline|4824,4831
.|4831,4832
<EOL>|4832,4833
<EOL>|4833,4834
-|4834,4835
Motor|4835,4840
:|4840,4841
Normal|4842,4848
bulk|4849,4853
,|4853,4854
tone|4855,4859
throughout|4860,4870
.|4870,4871
She|4872,4875
says|4876,4880
she|4881,4884
can|4885,4888
not|4888,4891
move|4892,4896
<EOL>|4896,4897
her|4897,4900
arms|4901,4905
.|4905,4906
When|4907,4911
arms|4912,4916
placed|4917,4923
over|4924,4928
her|4929,4932
head|4933,4937
,|4937,4938
her|4939,4942
arms|4943,4947
slowly|4948,4954
miss|4955,4959
<EOL>|4959,4960
her|4960,4963
face|4964,4968
and|4969,4972
slowly|4973,4979
drops|4980,4985
to|4986,4988
the|4989,4992
bed|4993,4996
in|4997,4999
a|5000,5001
controlled|5002,5012
fashion|5013,5020
.|5020,5021
<EOL>|5022,5023
She|5023,5026
<EOL>|5026,5027
does|5027,5031
lift|5032,5036
her|5037,5040
arms|5041,5045
to|5046,5048
hold|5049,5053
the|5054,5057
side|5058,5062
rails|5063,5068
of|5069,5071
the|5072,5075
bed|5076,5079
<EOL>|5079,5080
spontaneously|5080,5093
.|5093,5094
She|5095,5098
lifts|5099,5104
her|5105,5108
legs|5109,5113
antigravity|5114,5125
and|5126,5129
holds|5130,5135
them|5136,5140
<EOL>|5140,5141
without|5141,5148
drift|5149,5154
.|5154,5155
<EOL>|5155,5156
<EOL>|5156,5157
-|5157,5158
Sensory|5158,5165
:|5165,5166
slightly|5167,5175
withdrawals|5176,5187
in|5188,5190
upper|5191,5196
extremities|5197,5208
and|5209,5212
says|5213,5217
<EOL>|5217,5218
"|5218,5219
ouch|5219,5223
"|5223,5224
,|5224,5225
briskly|5226,5233
withdrawals|5234,5245
in|5246,5248
lower|5249,5254
extremities|5255,5266
to|5267,5269
noxious|5270,5277
<EOL>|5277,5278
stimuli|5278,5285
and|5286,5289
says|5290,5294
"|5295,5296
ouch|5296,5300
"|5300,5301
<EOL>|5301,5302
<EOL>|5302,5303
-|5303,5304
DTRs|5304,5308
:|5308,5309
<EOL>|5309,5310
_|5313,5314
_|5314,5315
_|5315,5316
Tri|5317,5320
_|5321,5322
_|5322,5323
_|5323,5324
Pat|5325,5328
Ach|5329,5332
<EOL>|5332,5333
L|5334,5335
2|5337,5338
2|5340,5341
0|5345,5346
3|5350,5351
2|5354,5355
<EOL>|5355,5356
R|5357,5358
2|5360,5361
2|5363,5364
0|5368,5369
3|5373,5374
2|5377,5378
<EOL>|5378,5379
Plantar|5380,5387
response|5388,5396
was|5397,5400
flexor|5401,5407
bilaterally|5408,5419
.|5419,5420
<EOL>|5420,5421
<EOL>|5421,5422
-|5422,5423
Coordination|5423,5435
:|5435,5436
patient|5437,5444
could|5445,5450
not|5451,5454
participate|5455,5466
<EOL>|5466,5467
<EOL>|5467,5468
-|5468,5469
Gait|5469,5473
:|5473,5474
could|5475,5480
not|5481,5484
assess|5485,5491
as|5492,5494
patient|5495,5502
would|5503,5508
not|5509,5512
get|5513,5516
out|5517,5520
of|5521,5523
bed|5524,5527
<EOL>|5527,5528
<EOL>|5528,5529
Discharge|5529,5538
Exam|5539,5543
:|5543,5544
<EOL>|5544,5545
General|5545,5552
:|5552,5553
sitting|5554,5561
up|5562,5564
in|5565,5567
her|5568,5571
chair|5572,5577
with|5578,5582
eyes|5583,5587
closed|5588,5594
<EOL>|5594,5595
HEENT|5595,5600
:|5600,5601
no|5602,5604
trauma|5605,5611
,|5611,5612
no|5613,5615
jaundice|5616,5624
,|5624,5625
no|5626,5628
lesions|5629,5636
of|5637,5639
oropharynx|5640,5650
<EOL>|5651,5652
CV|5652,5654
:|5654,5655
sinus|5656,5661
bradycardia|5662,5673
,|5673,5674
no|5675,5677
m|5678,5679
/|5679,5680
r|5680,5681
/|5681,5682
g|5682,5683
<EOL>|5683,5684
Pulm|5684,5688
:|5688,5689
Breathing|5690,5699
comfortably|5700,5711
on|5712,5714
RA|5715,5717
<EOL>|5718,5719
Ext|5719,5722
:|5722,5723
Warm|5724,5728
and|5729,5732
well|5733,5737
perfused|5738,5746
,|5746,5747
no|5748,5750
rash|5751,5755
or|5756,5758
mottling|5759,5767
<EOL>|5767,5768
<EOL>|5768,5769
Neurologic|5769,5779
:|5779,5780
<EOL>|5780,5781
<EOL>|5781,5782
-|5782,5783
Mental|5783,5789
Status|5790,5796
:|5796,5797
Answering|5798,5807
questions|5808,5817
with|5818,5822
slow|5823,5827
short|5828,5833
sentence|5834,5842
.|5842,5843
<EOL>|5843,5844
More|5844,5848
humor|5849,5854
and|5855,5858
complex|5859,5866
sentences|5867,5876
observed|5877,5885
today|5886,5891
.|5891,5892
<EOL>|5892,5893
Eyes|5893,5897
intermittently|5898,5912
close|5913,5918
while|5919,5924
she|5925,5928
is|5929,5931
talking|5932,5939
.|5939,5940
Speech|5941,5947
<EOL>|5947,5948
is|5948,5950
not|5951,5954
dysarthric|5955,5965
,|5965,5966
no|5967,5969
spontaneous|5970,5981
speech|5982,5988
output|5989,5995
.|5995,5996
Follows|5997,6004
<EOL>|6004,6005
simple|6005,6011
commands|6012,6020
.|6020,6021
<EOL>|6021,6022
<EOL>|6022,6023
-|6023,6024
Cranial|6024,6031
Nerves|6032,6038
:|6038,6039
<EOL>|6039,6040
II|6040,6042
,|6042,6043
III|6044,6047
,|6047,6048
IV|6049,6051
,|6051,6052
VI|6053,6055
:|6055,6056
Pupils|6057,6063
8|6064,6065
mm|6066,6068
-|6068,6069
>|6069,6070
4|6070,6071
mm|6072,6074
.|6074,6075
EOMI|6076,6080
without|6081,6088
nystagmus|6089,6098
.|6098,6099
<EOL>|6100,6101
V|6101,6102
:|6102,6103
facial|6104,6110
sensation|6111,6120
intact|6121,6127
throughout|6128,6138
<EOL>|6138,6139
VII|6139,6142
:|6142,6143
No|6144,6146
facial|6147,6153
droop|6154,6159
,|6159,6160
facial|6161,6167
musculature|6168,6179
symmetric|6180,6189
with|6190,6194
grimace|6195,6202
<EOL>|6202,6203
but|6203,6206
limited|6207,6214
facial|6215,6221
movements|6222,6231
.|6231,6232
<EOL>|6232,6233
IX|6233,6235
,|6235,6236
X|6237,6238
,|6238,6239
XII|6240,6243
:|6243,6244
palate|6245,6251
elevates|6252,6260
symmetrically|6261,6274
,|6274,6275
tongue|6276,6282
midline|6283,6290
<EOL>|6290,6291
<EOL>|6291,6292
-|6292,6293
Motor|6293,6298
:|6298,6299
Normal|6300,6306
bulk|6307,6311
,|6311,6312
tone|6313,6317
throughout|6318,6328
.|6328,6329
Lifting|6330,6337
arms|6338,6342
and|6343,6346
legs|6347,6351
<EOL>|6351,6352
against|6352,6359
gravity|6360,6367
but|6368,6371
not|6372,6375
against|6376,6383
resistance|6384,6394
(|6395,6396
_|6396,6397
_|6397,6398
_|6398,6399
)|6399,6400
<EOL>|6400,6401
<EOL>|6401,6402
-|6402,6403
Sensory|6403,6410
:|6410,6411
Sensation|6412,6421
intact|6422,6428
to|6429,6431
touch|6432,6437
and|6438,6441
temperature|6442,6453
throughout|6454,6464
<EOL>|6464,6465
<EOL>|6465,6466
-|6466,6467
DTRs|6467,6471
:|6471,6472
1|6473,6474
+|6474,6475
patellar|6476,6484
,|6484,6485
biceps|6486,6492
,|6492,6493
brachioradialis|6494,6509
throughout|6510,6520
<EOL>|6520,6521
<EOL>|6521,6522
-|6522,6523
Coordination|6523,6535
:|6535,6536
No|6537,6539
dysmetria|6540,6549
or|6550,6552
tremor|6553,6559
.|6559,6560
<EOL>|6561,6562
<EOL>|6562,6563
-|6563,6564
Gait|6564,6568
:|6568,6569
Ambulated|6570,6579
well|6580,6584
with|6585,6589
a|6590,6591
_|6592,6593
_|6593,6594
_|6594,6595
.|6595,6596
<EOL>|6596,6597
<EOL>|6598,6599
Pertinent|6599,6608
Results|6609,6616
:|6616,6617
<EOL>|6617,6618
Admission|6618,6627
labs|6628,6632
:|6632,6633
<EOL>|6633,6634
=|6634,6635
=|6635,6636
=|6636,6637
=|6637,6638
=|6638,6639
=|6639,6640
=|6640,6641
=|6641,6642
=|6642,6643
=|6643,6644
=|6644,6645
=|6645,6646
=|6646,6647
=|6647,6648
=|6648,6649
<EOL>|6649,6650
_|6650,6651
_|6651,6652
_|6652,6653
12|6654,6656
:|6656,6657
59PM|6657,6661
GLUCOSE|6664,6671
-|6671,6672
77|6672,6674
UREA|6675,6679
N|6680,6681
-|6681,6682
8|6682,6683
CREAT|6684,6689
-|6689,6690
0.7|6690,6693
SODIUM|6694,6700
-|6700,6701
142|6701,6704
<EOL>|6705,6706
POTASSIUM|6706,6715
-|6715,6716
3.8|6716,6719
CHLORIDE|6720,6728
-|6728,6729
104|6729,6732
TOTAL|6733,6738
CO2|6739,6742
-|6742,6743
24|6743,6745
ANION|6746,6751
GAP|6752,6755
-|6755,6756
14|6756,6758
<EOL>|6758,6759
_|6759,6760
_|6760,6761
_|6761,6762
12|6763,6765
:|6765,6766
59PM|6766,6770
ALT|6773,6776
(|6776,6777
SGPT|6777,6781
)|6781,6782
-|6782,6783
9|6783,6784
AST|6785,6788
(|6788,6789
SGOT|6789,6793
)|6793,6794
-|6794,6795
13|6795,6797
ALK|6798,6801
PHOS|6802,6806
-|6806,6807
39|6807,6809
TOT|6810,6813
<EOL>|6814,6815
BILI|6815,6819
-|6819,6820
0.3|6820,6823
<EOL>|6823,6824
_|6824,6825
_|6825,6826
_|6826,6827
12|6828,6830
:|6830,6831
59PM|6831,6835
CALCIUM|6838,6845
-|6845,6846
8.7|6846,6849
PHOSPHATE|6850,6859
-|6859,6860
4.0|6860,6863
MAGNESIUM|6864,6873
-|6873,6874
1.7|6874,6877
<EOL>|6877,6878
_|6878,6879
_|6879,6880
_|6880,6881
12|6882,6884
:|6884,6885
59PM|6885,6889
tTG|6892,6895
-|6895,6896
IgA|6896,6899
-|6899,6900
7|6900,6901
<EOL>|6901,6902
_|6902,6903
_|6903,6904
_|6904,6905
12|6906,6908
:|6908,6909
59PM|6909,6913
WBC|6916,6919
-|6919,6920
5.0|6920,6923
RBC|6924,6927
-|6927,6928
3|6928,6929
.|6929,6930
89|6930,6932
*|6932,6933
HGB|6934,6937
-|6937,6938
11.5|6938,6942
HCT|6943,6946
-|6946,6947
34.4|6947,6951
MCV|6952,6955
-|6955,6956
88|6956,6958
<EOL>|6959,6960
MCH|6960,6963
-|6963,6964
29.6|6964,6968
MCHC|6969,6973
-|6973,6974
33.4|6974,6978
RDW|6979,6982
-|6982,6983
12.4|6983,6987
RDWSD|6988,6993
-|6993,6994
39.8|6994,6998
<EOL>|6998,6999
_|6999,7000
_|7000,7001
_|7001,7002
12|7003,7005
:|7005,7006
59PM|7006,7010
PLT|7013,7016
COUNT|7017,7022
-|7022,7023
235|7023,7026
<EOL>|7026,7027
_|7027,7028
_|7028,7029
_|7029,7030
05|7031,7033
:|7033,7034
11AM|7034,7038
URINE|7039,7044
HOURS|7046,7051
-|7051,7052
RANDOM|7052,7058
<EOL>|7058,7059
_|7059,7060
_|7060,7061
_|7061,7062
05|7063,7065
:|7065,7066
11AM|7066,7070
URINE|7071,7076
UCG|7078,7081
-|7081,7082
NEGATIVE|7082,7090
<EOL>|7090,7091
_|7091,7092
_|7092,7093
_|7093,7094
05|7095,7097
:|7097,7098
11AM|7098,7102
URINE|7103,7108
bnzodzpn|7110,7118
-|7118,7119
NEG|7119,7122
barbitrt|7123,7131
-|7131,7132
NEG|7132,7135
opiates|7136,7143
-|7143,7144
NEG|7144,7147
<EOL>|7148,7149
cocaine|7149,7156
-|7156,7157
NEG|7157,7160
amphetmn|7161,7169
-|7169,7170
NEG|7170,7173
oxycodn|7174,7181
-|7181,7182
NEG|7182,7185
mthdone|7186,7193
-|7193,7194
NEG|7194,7197
<EOL>|7197,7198
_|7198,7199
_|7199,7200
_|7200,7201
05|7202,7204
:|7204,7205
11AM|7205,7209
URINE|7210,7215
COLOR|7217,7222
-|7222,7223
Straw|7223,7228
APPEAR|7229,7235
-|7235,7236
Clear|7236,7241
SP|7242,7244
_|7245,7246
_|7246,7247
_|7247,7248
<EOL>|7248,7249
_|7249,7250
_|7250,7251
_|7251,7252
05|7253,7255
:|7255,7256
11AM|7256,7260
URINE|7261,7266
BLOOD|7268,7273
-|7273,7274
LG|7274,7276
*|7276,7277
NITRITE|7278,7285
-|7285,7286
NEG|7286,7289
PROTEIN|7290,7297
-|7297,7298
NEG|7298,7301
<EOL>|7302,7303
GLUCOSE|7303,7310
-|7310,7311
NEG|7311,7314
KETONE|7315,7321
-|7321,7322
TR|7322,7324
*|7324,7325
BILIRUBIN|7326,7335
-|7335,7336
NEG|7336,7339
UROBILNGN|7340,7349
-|7349,7350
NEG|7350,7353
PH|7354,7356
-|7356,7357
7.0|7357,7360
<EOL>|7361,7362
LEUK|7362,7366
-|7366,7367
NEG|7367,7370
<EOL>|7370,7371
_|7371,7372
_|7372,7373
_|7373,7374
05|7375,7377
:|7377,7378
11AM|7378,7382
URINE|7383,7388
RBC|7390,7393
-|7393,7394
5|7394,7395
*|7395,7396
WBC|7397,7400
-|7400,7401
1|7401,7402
BACTERIA|7403,7411
-|7411,7412
FEW|7412,7415
*|7415,7416
YEAST|7417,7422
-|7422,7423
NONE|7423,7427
<EOL>|7428,7429
EPI|7429,7432
-|7432,7433
0|7433,7434
<EOL>|7434,7435
_|7435,7436
_|7436,7437
_|7437,7438
05|7439,7441
:|7441,7442
11AM|7442,7446
URINE|7447,7452
MUCOUS|7454,7460
-|7460,7461
RARE|7461,7465
*|7465,7466
<EOL>|7466,7467
_|7467,7468
_|7468,7469
_|7469,7470
04|7471,7473
:|7473,7474
34AM|7474,7478
_|7481,7482
_|7482,7483
_|7483,7484
PTT|7485,7488
-|7488,7489
27.2|7489,7493
_|7494,7495
_|7495,7496
_|7496,7497
<EOL>|7497,7498
_|7498,7499
_|7499,7500
_|7500,7501
04|7502,7504
:|7504,7505
28AM|7505,7509
WBC|7512,7515
-|7515,7516
6.4|7516,7519
RBC|7520,7523
-|7523,7524
4|7524,7525
.|7525,7526
17|7526,7528
HGB|7529,7532
-|7532,7533
12.6|7533,7537
HCT|7538,7541
-|7541,7542
37.4|7542,7546
MCV|7547,7550
-|7550,7551
90|7551,7553
<EOL>|7554,7555
MCH|7555,7558
-|7558,7559
30.2|7559,7563
MCHC|7564,7568
-|7568,7569
33.7|7569,7573
RDW|7574,7577
-|7577,7578
12.4|7578,7582
RDWSD|7583,7588
-|7588,7589
40.8|7589,7593
<EOL>|7593,7594
_|7594,7595
_|7595,7596
_|7596,7597
04|7598,7600
:|7600,7601
28AM|7601,7605
NEUTS|7608,7613
-|7613,7614
58.2|7614,7618
_|7619,7620
_|7620,7621
_|7621,7622
MONOS|7623,7628
-|7628,7629
7.1|7629,7632
EOS|7633,7636
-|7636,7637
0|7637,7638
.|7638,7639
2|7639,7640
*|7640,7641
<EOL>|7642,7643
BASOS|7643,7648
-|7648,7649
0.6|7649,7652
IM|7653,7655
_|7656,7657
_|7657,7658
_|7658,7659
AbsNeut|7660,7667
-|7667,7668
3|7668,7669
.|7669,7670
70|7670,7672
AbsLymp|7673,7680
-|7680,7681
2.14|7681,7685
AbsMono|7686,7693
-|7693,7694
0|7694,7695
.|7695,7696
45|7696,7698
<EOL>|7699,7700
AbsEos|7700,7706
-|7706,7707
0|7707,7708
.|7708,7709
01|7709,7711
*|7711,7712
AbsBaso|7713,7720
-|7720,7721
0.04|7721,7725
<EOL>|7725,7726
_|7726,7727
_|7727,7728
_|7728,7729
04|7730,7732
:|7732,7733
28AM|7733,7737
PLT|7740,7743
COUNT|7744,7749
-|7749,7750
246|7750,7753
<EOL>|7753,7754
_|7754,7755
_|7755,7756
_|7756,7757
04|7758,7760
:|7760,7761
11AM|7761,7765
_|7768,7769
_|7769,7770
_|7770,7771
PO2|7772,7775
-|7775,7776
50|7776,7778
*|7778,7779
PCO2|7780,7784
-|7784,7785
34|7785,7787
*|7787,7788
PH|7789,7791
-|7791,7792
7.44|7792,7796
TOTAL|7797,7802
<EOL>|7803,7804
CO2|7804,7807
-|7807,7808
24|7808,7810
BASE|7811,7815
XS|7816,7818
-|7818,7819
0|7819,7820
COMMENTS|7821,7829
-|7829,7830
GREEN|7830,7835
TOP|7836,7839
<EOL>|7839,7840
_|7840,7841
_|7841,7842
_|7842,7843
04|7844,7846
:|7846,7847
10AM|7847,7851
GLUCOSE|7854,7861
-|7861,7862
84|7862,7864
UREA|7865,7869
N|7870,7871
-|7871,7872
7|7872,7873
CREAT|7874,7879
-|7879,7880
0.8|7880,7883
SODIUM|7884,7890
-|7890,7891
143|7891,7894
<EOL>|7895,7896
POTASSIUM|7896,7905
-|7905,7906
3.6|7906,7909
CHLORIDE|7910,7918
-|7918,7919
106|7919,7922
TOTAL|7923,7928
CO2|7929,7932
-|7932,7933
23|7933,7935
ANION|7936,7941
GAP|7942,7945
-|7945,7946
14|7946,7948
<EOL>|7948,7949
_|7949,7950
_|7950,7951
_|7951,7952
04|7953,7955
:|7955,7956
10AM|7956,7960
estGFR|7963,7969
-|7969,7970
Using|7970,7975
this|7976,7980
<EOL>|7980,7981
_|7981,7982
_|7982,7983
_|7983,7984
04|7985,7987
:|7987,7988
10AM|7988,7992
ALT|7995,7998
(|7998,7999
SGPT|7999,8003
)|8003,8004
-|8004,8005
9|8005,8006
AST|8007,8010
(|8010,8011
SGOT|8011,8015
)|8015,8016
-|8016,8017
14|8017,8019
CK|8020,8022
(|8022,8023
CPK|8023,8026
)|8026,8027
-|8027,8028
67|8028,8030
ALK|8031,8034
<EOL>|8035,8036
PHOS|8036,8040
-|8040,8041
41|8041,8043
TOT|8044,8047
BILI|8048,8052
-|8052,8053
0.3|8053,8056
<EOL>|8056,8057
_|8057,8058
_|8058,8059
_|8059,8060
04|8061,8063
:|8063,8064
10AM|8064,8068
CK|8071,8073
-|8073,8074
MB|8074,8076
-|8076,8077
<|8077,8078
1|8078,8079
<EOL>|8079,8080
_|8080,8081
_|8081,8082
_|8082,8083
04|8084,8086
:|8086,8087
10AM|8087,8091
ALBUMIN|8094,8101
-|8101,8102
3.9|8102,8105
CALCIUM|8106,8113
-|8113,8114
8.8|8114,8117
PHOSPHATE|8118,8127
-|8127,8128
2.9|8128,8131
<EOL>|8132,8133
MAGNESIUM|8133,8142
-|8142,8143
1.8|8143,8146
<EOL>|8146,8147
_|8147,8148
_|8148,8149
_|8149,8150
04|8151,8153
:|8153,8154
10AM|8154,8158
VIT|8161,8164
B12|8165,8168
-|8168,8169
227|8169,8172
*|8172,8173
<EOL>|8173,8174
_|8174,8175
_|8175,8176
_|8176,8177
04|8178,8180
:|8180,8181
10AM|8181,8185
TSH|8188,8191
-|8191,8192
2.7|8192,8195
<EOL>|8195,8196
_|8196,8197
_|8197,8198
_|8198,8199
04|8200,8202
:|8202,8203
10AM|8203,8207
TSH|8210,8213
-|8213,8214
2.6|8214,8217
<EOL>|8217,8218
_|8218,8219
_|8219,8220
_|8220,8221
04|8222,8224
:|8224,8225
10AM|8225,8229
_|8232,8233
_|8233,8234
_|8234,8235
TITER|8236,8241
-|8241,8242
1|8242,8243
:|8243,8244
1280|8244,8248
*|8248,8249
CRP|8250,8253
-|8253,8254
3.4|8254,8257
<EOL>|8258,8259
dsDNA|8259,8264
-|8264,8265
NEGATIVE|8265,8273
<EOL>|8273,8274
_|8274,8275
_|8275,8276
_|8276,8277
04|8278,8280
:|8280,8281
10AM|8281,8285
C3|8288,8290
-|8290,8291
121|8291,8294
C4|8295,8297
-|8297,8298
27|8298,8300
<EOL>|8300,8301
_|8301,8302
_|8302,8303
_|8303,8304
04|8305,8307
:|8307,8308
10AM|8308,8312
ASA|8315,8318
-|8318,8319
NEG|8319,8322
ETHANOL|8323,8330
-|8330,8331
NEG|8331,8334
ACETMNPHN|8335,8344
-|8344,8345
NEG|8345,8348
<EOL>|8349,8350
tricyclic|8350,8359
-|8359,8360
NEG|8360,8363
<EOL>|8363,8364
<EOL>|8364,8365
EEG|8365,8368
_|8369,8370
_|8370,8371
_|8371,8372
:|8372,8373
<EOL>|8373,8374
=|8374,8375
=|8375,8376
=|8376,8377
=|8377,8378
=|8378,8379
=|8379,8380
=|8380,8381
=|8381,8382
=|8382,8383
=|8383,8384
=|8384,8385
=|8385,8386
=|8386,8387
=|8387,8388
<EOL>|8388,8389
IMPRESSION|8389,8399
:|8399,8400
This|8401,8405
telemetry|8406,8415
captured|8416,8424
no|8425,8427
pushbutton|8428,8438
activations|8439,8450
.|8450,8451
<EOL>|8452,8453
The|8453,8456
background|8457,8467
showed|8468,8474
normal|8475,8481
waking|8482,8488
and|8489,8492
sleep|8493,8498
patterns|8499,8507
.|8507,8508
There|8509,8514
<EOL>|8515,8516
were|8516,8520
no|8521,8523
focal|8524,8529
abnormalities|8530,8543
,|8543,8544
epileptiform|8545,8557
features|8558,8566
,|8566,8567
or|8568,8570
<EOL>|8571,8572
electrographic|8572,8586
seizures|8587,8595
.|8595,8596
A|8597,8598
bradycardia|8599,8610
was|8611,8614
noted|8615,8620
.|8620,8621
<EOL>|8622,8623
<EOL>|8623,8624
IMAGING|8624,8631
:|8631,8632
<EOL>|8632,8633
=|8633,8634
=|8634,8635
=|8635,8636
=|8636,8637
=|8637,8638
=|8638,8639
=|8639,8640
=|8640,8641
<EOL>|8641,8642
MRI|8642,8645
BRAIN|8646,8651
WITH|8652,8656
/|8656,8657
WITHOUT|8657,8664
CONTRAST|8665,8673
_|8674,8675
_|8675,8676
_|8676,8677
<EOL>|8677,8678
<EOL>|8678,8679
:|8687,8688
<EOL>|8690,8691
<EOL>|8693,8694
A|8694,8695
5|8696,8697
mm|8698,8700
FLAIR|8701,8706
hypointense|8707,8718
and|8719,8722
T1|8723,8725
isointense|8726,8736
lesion|8737,8743
at|8744,8746
midline|8747,8754
<EOL>|8755,8756
between|8756,8763
the|8764,8767
<EOL>|8768,8769
anterior|8769,8777
and|8778,8781
posterior|8782,8791
pituitary|8792,8801
is|8802,8804
noted|8805,8810
.|8810,8811
There|8812,8817
is|8818,8820
no|8821,8823
evidence|8824,8832
<EOL>|8833,8834
of|8834,8836
<EOL>|8837,8838
hemorrhage|8838,8848
,|8848,8849
edema|8850,8855
,|8855,8856
mass|8857,8861
effect|8862,8868
,|8868,8869
midline|8870,8877
shift|8878,8883
or|8884,8886
infarction|8887,8897
.|8897,8898
The|8899,8902
<EOL>|8903,8904
ventricles|8904,8914
and|8915,8918
sulci|8919,8924
are|8925,8928
normal|8929,8935
in|8936,8938
caliber|8939,8946
and|8947,8950
configuration|8951,8964
.|8964,8965
<EOL>|8966,8967
There|8967,8972
is|8973,8975
no|8976,8978
abnormal|8979,8987
enhancement|8988,8999
after|9000,9005
contrast|9006,9014
administration|9015,9029
.|9029,9030
<EOL>|9031,9032
<EOL>|9034,9035
A|9052,9053
5|9054,9055
mm|9056,9058
FLAIR|9059,9064
hypointense|9065,9076
and|9077,9080
T1|9081,9083
isointense|9084,9094
lesion|9095,9101
at|9102,9104
midline|9105,9112
<EOL>|9113,9114
between|9114,9121
the|9122,9125
<EOL>|9126,9127
anterior|9127,9135
and|9136,9139
posterior|9140,9149
pituitary|9150,9159
likely|9160,9166
represents|9167,9177
a|9178,9179
Rathke|9180,9186
's|9186,9188
<EOL>|9189,9190
cleft|9190,9195
cyst|9196,9200
.|9200,9201
<EOL>|9203,9204
Further|9204,9211
evaluation|9212,9222
is|9223,9225
needed|9226,9232
,|9232,9233
dedicated|9234,9243
pituitary|9244,9253
MR|9254,9256
may|9257,9260
be|9261,9263
<EOL>|9264,9265
obtained|9265,9273
.|9273,9274
<EOL>|9275,9276
<EOL>|9278,9279
<EOL>|9279,9280
<EOL>|9281,9282
See|9305,9308
worksheet|9309,9318
<EOL>|9318,9319
<EOL>|9320,9321
Medications|9321,9332
on|9333,9335
Admission|9336,9345
:|9345,9346
<EOL>|9346,9347
famotidine|9347,9357
40|9358,9360
mg|9361,9363
daily|9364,9369
<EOL>|9369,9370
birth|9370,9375
control|9376,9383
per|9384,9387
her|9388,9391
aunt|9392,9396
<EOL>|9396,9397
<EOL>|9398,9399
_|9399,9400
_|9400,9401
_|9401,9402
:|9402,9403
<EOL>|9403,9404
1.|9404,9406
_|9408,9409
_|9409,9410
_|9410,9411
250|9412,9415
mcg|9416,9419
PO|9420,9422
DAILY|9423,9428
<EOL>|9430,9431
2.|9431,9433
Famotidine|9435,9445
40|9446,9448
mg|9449,9451
PO|9452,9454
DAILY|9455,9460
<EOL>|9462,9463
3.|9463,9465
Metoprolol|9467,9477
Tartrate|9478,9486
12.5|9487,9491
mg|9492,9494
PO|9495,9497
DAILY|9498,9503
<EOL>|9505,9506
4.|9506,9508
Multivitamins|9510,9523
W|9524,9525
/|9525,9526
minerals|9526,9534
1|9535,9536
TAB|9537,9540
PO|9541,9543
DAILY|9544,9549
<EOL>|9551,9552
5.|9552,9554
Nortriptyline|9556,9569
10|9570,9572
mg|9573,9575
PO|9576,9578
QHS|9579,9582
<EOL>|9584,9585
6.|9585,9587
_|9589,9590
_|9590,9591
_|9591,9592
1|9593,9594
item|9595,9599
miscellaneous|9600,9613
ONCE|9614,9618
<EOL>|9619,9620
Prognosis|9620,9629
:|9629,9630
Good|9631,9635
<EOL>|9635,9636
_|9636,9637
_|9637,9638
_|9638,9639
:|9639,9640
13|9641,9643
months|9644,9650
<EOL>|9651,9652
RX|9652,9654
_|9655,9656
_|9656,9657
_|9657,9658
Once|9661,9665
Disp|9666,9670
#|9671,9672
*|9672,9673
1|9673,9674
Each|9675,9679
Refills|9680,9687
:|9687,9688
*|9688,9689
0|9689,9690
<EOL>|9691,9692
<EOL>|9692,9693
<EOL>|9694,9695
Discharge|9695,9704
Disposition|9705,9716
:|9716,9717
<EOL>|9717,9718
Extended|9718,9726
Care|9727,9731
<EOL>|9731,9732
<EOL>|9733,9734
Facility|9734,9742
:|9742,9743
<EOL>|9743,9744
_|9744,9745
_|9745,9746
_|9746,9747
<EOL>|9747,9748
<EOL>|9749,9750
Discharge|9750,9759
Diagnosis|9760,9769
:|9769,9770
<EOL>|9770,9771
Functional|9771,9781
neurological|9782,9794
syndrome|9795,9803
<EOL>|9804,9805
<EOL>|9805,9806
<EOL>|9807,9808
Mental|9829,9835
Status|9836,9842
:|9842,9843
Clear|9844,9849
and|9850,9853
coherent|9854,9862
.|9862,9863
<EOL>|9863,9864
Level|9864,9869
of|9870,9872
Consciousness|9873,9886
:|9886,9887
Lethargic|9888,9897
but|9898,9901
arousable|9902,9911
.|9911,9912
<EOL>|9912,9913
Activity|9913,9921
Status|9922,9928
:|9928,9929
Ambulatory|9930,9940
-|9941,9942
Independent|9943,9954
.|9954,9955
<EOL>|9955,9956
<EOL>|9956,9957
<EOL>|9958,9959
Dear|9983,9987
Ms.|9988,9991
_|9992,9993
_|9993,9994
_|9994,9995
,|9995,9996
<EOL>|9996,9997
<EOL>|9997,9998
It|9998,10000
was|10001,10004
a|10005,10006
pleasure|10007,10015
taking|10016,10022
care|10023,10027
of|10028,10030
you|10031,10034
at|10035,10037
_|10038,10039
_|10039,10040
_|10040,10041
<EOL>|10042,10043
_|10043,10044
_|10044,10045
_|10045,10046
.|10046,10047
<EOL>|10047,10048
<EOL>|10048,10049
You|10049,10052
were|10053,10057
in|10058,10060
the|10061,10064
hospital|10065,10073
because|10074,10081
of|10082,10084
headache|10085,10093
,|10093,10094
lethargy|10095,10103
,|10103,10104
and|10105,10108
<EOL>|10109,10110
weakness|10110,10118
after|10119,10124
an|10125,10127
iron|10128,10132
infusion|10133,10141
.|10141,10142
<EOL>|10142,10143
<EOL>|10143,10144
You|10144,10147
had|10148,10151
a|10152,10153
number|10154,10160
of|10161,10163
tests|10164,10169
performed|10170,10179
in|10180,10182
the|10183,10186
hospital|10187,10195
,|10195,10196
all|10197,10200
of|10201,10203
<EOL>|10204,10205
which|10205,10210
were|10211,10215
reassuring|10216,10226
.|10226,10227
An|10228,10230
MRI|10231,10234
of|10235,10237
your|10238,10242
brain|10243,10248
showed|10249,10255
no|10256,10258
evidence|10259,10267
<EOL>|10268,10269
of|10269,10271
stroke|10272,10278
or|10279,10281
inflammation|10282,10294
.|10294,10295
An|10296,10298
EEG|10299,10302
to|10303,10305
monitor|10306,10313
your|10314,10318
brain|10319,10324
waves|10325,10330
<EOL>|10331,10332
showed|10332,10338
no|10339,10341
evidence|10342,10350
of|10351,10353
seizure|10354,10361
.|10361,10362
Your|10363,10367
weakness|10368,10376
gradually|10377,10386
improved|10387,10395
<EOL>|10396,10397
over|10397,10401
the|10402,10405
course|10406,10412
of|10413,10415
your|10416,10420
hospitalization|10421,10436
and|10437,10440
will|10441,10445
continue|10446,10454
to|10455,10457
<EOL>|10458,10459
improve|10459,10466
after|10467,10472
you|10473,10476
leave|10477,10482
the|10483,10486
hospital|10487,10495
.|10495,10496
<EOL>|10497,10498
<EOL>|10498,10499
After|10499,10504
leaving|10505,10512
the|10513,10516
hospital|10517,10525
,|10525,10526
you|10527,10530
should|10531,10537
continue|10538,10546
to|10547,10549
work|10550,10554
on|10555,10557
<EOL>|10558,10559
improving|10559,10568
your|10569,10573
strength|10574,10582
.|10582,10583
It|10584,10586
will|10587,10591
improve|10592,10599
as|10600,10602
long|10603,10607
as|10608,10610
you|10611,10614
work|10615,10619
<EOL>|10620,10621
hard|10621,10625
!|10625,10626
<EOL>|10626,10627
<EOL>|10627,10628
We|10628,10630
wish|10631,10635
you|10636,10639
the|10640,10643
best|10644,10648
,|10648,10649
<EOL>|10649,10650
Your|10650,10654
_|10655,10656
_|10656,10657
_|10657,10658
Care|10659,10663
Team|10664,10668
<EOL>|10668,10669
<EOL>|10670,10671
Followup|10671,10679
Instructions|10680,10692
:|10692,10693
<EOL>|10693,10694
_|10694,10695
_|10695,10696
_|10696,10697
<EOL>|10697,10698

