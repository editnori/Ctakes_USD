 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
amoxicillin|179,190
/|191,192
iron|193,197
<EOL>|197,198
<EOL>|199,200
Attending|200,209
:|209,210
_|211,212
_|212,213
_|213,214
.|214,215
<EOL>|215,216
<EOL>|217,218
Major|218,223
Surgical|224,232
or|233,235
Invasive|236,244
Procedure|245,254
:|254,255
<EOL>|255,256
None|256,260
<EOL>|260,261
<EOL>|261,262
attach|262,268
<EOL>|268,269
<EOL>|270,271
Pertinent|271,280
Results|281,288
:|288,289
<EOL>|289,290
ADMISSION|290,299
LABS|300,304
:|304,305
<EOL>|305,306
=|306,307
=|307,308
=|308,309
=|309,310
=|310,311
=|311,312
=|312,313
=|313,314
=|314,315
=|315,316
=|316,317
=|317,318
=|318,319
=|319,320
=|320,321
<EOL>|321,322
_|322,323
_|323,324
_|324,325
10|326,328
:|328,329
45PM|329,333
PLT|336,339
COUNT|340,345
-|345,346
244|346,349
<EOL>|349,350
_|350,351
_|351,352
_|352,353
10|354,356
:|356,357
45PM|357,361
NEUTS|364,369
-|369,370
55.7|370,374
_|375,376
_|376,377
_|377,378
MONOS|379,384
-|384,385
10.8|385,389
EOS|390,393
-|393,394
0|394,395
.|395,396
7|396,397
*|397,398
<EOL>|399,400
BASOS|400,405
-|405,406
0.9|406,409
IM|410,412
_|413,414
_|414,415
_|415,416
AbsNeut|417,424
-|424,425
2|425,426
.|426,427
99|427,429
AbsLymp|430,437
-|437,438
1|438,439
.|439,440
70|440,442
AbsMono|443,450
-|450,451
0|451,452
.|452,453
58|453,455
<EOL>|456,457
AbsEos|457,463
-|463,464
0|464,465
.|465,466
04|466,468
AbsBaso|469,476
-|476,477
0|477,478
.|478,479
05|479,481
<EOL>|481,482
_|482,483
_|483,484
_|484,485
10|486,488
:|488,489
45PM|489,493
WBC|496,499
-|499,500
5.4|500,503
RBC|504,507
-|507,508
4|508,509
.|509,510
19|510,512
HGB|513,516
-|516,517
13.4|517,521
HCT|522,525
-|525,526
41.2|526,530
MCV|531,534
-|534,535
98|535,537
<EOL>|538,539
MCH|539,542
-|542,543
32.0|543,547
MCHC|548,552
-|552,553
32.5|553,557
RDW|558,561
-|561,562
12.4|562,566
RDWSD|567,572
-|572,573
44.2|573,577
<EOL>|577,578
_|578,579
_|579,580
_|580,581
10|582,584
:|584,585
45PM|585,589
ASA|592,595
-|595,596
NEG|596,599
ETHANOL|600,607
-|607,608
NEG|608,611
ACETMNPHN|612,621
-|621,622
NEG|622,625
<EOL>|626,627
tricyclic|627,636
-|636,637
NEG|637,640
<EOL>|640,641
_|641,642
_|642,643
_|643,644
10|645,647
:|647,648
45PM|648,652
ALBUMIN|655,662
-|662,663
4.8|663,666
CALCIUM|667,674
-|674,675
9.6|675,678
PHOSPHATE|679,688
-|688,689
3.0|689,692
<EOL>|693,694
MAGNESIUM|694,703
-|703,704
2.1|704,707
<EOL>|707,708
_|708,709
_|709,710
_|710,711
10|712,714
:|714,715
45PM|715,719
LIPASE|722,728
-|728,729
31|729,731
<EOL>|731,732
_|732,733
_|733,734
_|734,735
10|736,738
:|738,739
45PM|739,743
ALT|746,749
(|749,750
SGPT|750,754
)|754,755
-|755,756
20|756,758
AST|759,762
(|762,763
SGOT|763,767
)|767,768
-|768,769
26|769,771
ALK|772,775
PHOS|776,780
-|780,781
48|781,783
TOT|784,787
<EOL>|788,789
BILI|789,793
-|793,794
0.4|794,797
<EOL>|797,798
_|798,799
_|799,800
_|800,801
10|802,804
:|804,805
45PM|805,809
GLUCOSE|812,819
-|819,820
128|820,823
*|823,824
UREA|825,829
N|830,831
-|831,832
15|832,834
CREAT|835,840
-|840,841
1.1|841,844
SODIUM|845,851
-|851,852
137|852,855
<EOL>|856,857
POTASSIUM|857,866
-|866,867
3.7|867,870
CHLORIDE|871,879
-|879,880
100|880,883
TOTAL|884,889
CO2|890,893
-|893,894
23|894,896
ANION|897,902
GAP|903,906
-|906,907
14|907,909
<EOL>|909,910
_|910,911
_|911,912
_|912,913
03|914,916
:|916,917
17AM|917,921
URINE|922,927
BLOOD|929,934
-|934,935
NEG|935,938
NITRITE|939,946
-|946,947
NEG|947,950
PROTEIN|951,958
-|958,959
NEG|959,962
<EOL>|963,964
GLUCOSE|964,971
-|971,972
NEG|972,975
KETONE|976,982
-|982,983
10|983,985
*|985,986
BILIRUBIN|987,996
-|996,997
NEG|997,1000
UROBILNGN|1001,1010
-|1010,1011
NORMAL|1011,1017
PH|1018,1020
-|1020,1021
6.5|1021,1024
<EOL>|1025,1026
LEUK|1026,1030
-|1030,1031
NEG|1031,1034
<EOL>|1034,1035
_|1035,1036
_|1036,1037
_|1037,1038
03|1039,1041
:|1041,1042
17AM|1042,1046
URINE|1047,1052
COLOR|1054,1059
-|1059,1060
Straw|1060,1065
APPEAR|1066,1072
-|1072,1073
CLEAR|1073,1078
SP|1079,1081
_|1082,1083
_|1083,1084
_|1084,1085
<EOL>|1085,1086
_|1086,1087
_|1087,1088
_|1088,1089
03|1090,1092
:|1092,1093
17AM|1093,1097
URINE|1098,1103
bnzodzpn|1105,1113
-|1113,1114
NEG|1114,1117
barbitrt|1118,1126
-|1126,1127
NEG|1127,1130
opiates|1131,1138
-|1138,1139
NEG|1139,1142
<EOL>|1143,1144
cocaine|1144,1151
-|1151,1152
NEG|1152,1155
amphetmn|1156,1164
-|1164,1165
NEG|1165,1168
oxycodn|1169,1176
-|1176,1177
NEG|1177,1180
mthdone|1181,1188
-|1188,1189
NEG|1189,1192
<EOL>|1192,1193
_|1193,1194
_|1194,1195
_|1195,1196
03|1197,1199
:|1199,1200
17AM|1200,1204
URINE|1205,1210
UCG|1212,1215
-|1215,1216
NEGATIVE|1216,1224
<EOL>|1224,1225
_|1225,1226
_|1226,1227
_|1227,1228
03|1229,1231
:|1231,1232
17AM|1232,1236
URINE|1237,1242
HOURS|1244,1249
-|1249,1250
RANDOM|1250,1256
<EOL>|1256,1257
<EOL>|1257,1258
PERTINENT|1258,1267
LABS|1268,1272
:|1272,1273
<EOL>|1273,1274
=|1274,1275
=|1275,1276
=|1276,1277
=|1277,1278
=|1278,1279
=|1279,1280
=|1280,1281
=|1281,1282
=|1282,1283
=|1283,1284
=|1284,1285
=|1285,1286
=|1286,1287
=|1287,1288
=|1288,1289
<EOL>|1289,1290
_|1290,1291
_|1291,1292
_|1292,1293
05|1294,1296
:|1296,1297
45AM|1297,1301
BLOOD|1302,1307
VitB12|1308,1314
-|1314,1315
956|1315,1318
*|1318,1319
<EOL>|1319,1320
_|1320,1321
_|1321,1322
_|1322,1323
05|1324,1326
:|1326,1327
45AM|1327,1331
BLOOD|1332,1337
TSH|1338,1341
-|1341,1342
0.99|1342,1346
<EOL>|1346,1347
_|1347,1348
_|1348,1349
_|1349,1350
05|1351,1353
:|1353,1354
45AM|1354,1358
BLOOD|1359,1364
Free|1365,1369
T4|1370,1372
-|1372,1373
1.3|1373,1376
<EOL>|1376,1377
_|1377,1378
_|1378,1379
_|1379,1380
05|1381,1383
:|1383,1384
45AM|1384,1388
BLOOD|1389,1394
VITAMIN|1395,1402
B1|1403,1405
-|1405,1406
WHOLE|1406,1411
BLOOD|1412,1417
-|1417,1418
PND|1418,1421
<EOL>|1421,1422
<EOL>|1422,1423
MICRO|1423,1428
:|1428,1429
<EOL>|1429,1430
=|1430,1431
=|1431,1432
=|1432,1433
=|1433,1434
=|1434,1435
=|1435,1436
<EOL>|1436,1437
_|1437,1438
_|1438,1439
_|1439,1440
3|1441,1442
:|1442,1443
17|1443,1445
am|1446,1448
URINE|1449,1454
<EOL>|1454,1455
<EOL>|1455,1456
*|1484,1485
*|1485,1486
FINAL|1486,1491
REPORT|1492,1498
_|1499,1500
_|1500,1501
_|1501,1502
<EOL>|1502,1503
<EOL>|1503,1504
URINE|1507,1512
CULTURE|1513,1520
(|1521,1522
Final|1522,1527
_|1528,1529
_|1529,1530
_|1530,1531
:|1531,1532
<EOL>|1533,1534
MIXED|1540,1545
BACTERIAL|1546,1555
FLORA|1556,1561
(|1562,1563
>|1564,1565
=|1565,1566
3|1567,1568
COLONY|1569,1575
TYPES|1576,1581
)|1581,1582
,|1582,1583
CONSISTENT|1584,1594
<EOL>|1595,1596
WITH|1596,1600
SKIN|1601,1605
<EOL>|1605,1606
AND|1612,1615
/|1615,1616
OR|1616,1618
GENITAL|1619,1626
CONTAMINATION|1627,1640
.|1640,1641
<EOL>|1642,1643
<EOL>|1643,1644
IMAGING|1644,1651
:|1651,1652
<EOL>|1652,1653
=|1653,1654
=|1654,1655
=|1655,1656
=|1656,1657
=|1657,1658
=|1658,1659
=|1659,1660
=|1660,1661
<EOL>|1661,1662
none|1662,1666
<EOL>|1666,1667
<EOL>|1667,1668
DISCHARGE|1668,1677
LABS|1678,1682
:|1682,1683
<EOL>|1683,1684
=|1684,1685
=|1685,1686
=|1686,1687
=|1687,1688
=|1688,1689
=|1689,1690
=|1690,1691
=|1691,1692
=|1692,1693
=|1693,1694
=|1694,1695
=|1695,1696
=|1696,1697
=|1697,1698
=|1698,1699
<EOL>|1699,1700
no|1700,1702
labs|1703,1707
on|1708,1710
day|1711,1714
of|1715,1717
discharge|1718,1727
<EOL>|1727,1728
<EOL>|1728,1729
DISCHARGE|1729,1738
PHYSICAL|1739,1747
EXAM|1748,1752
:|1752,1753
<EOL>|1753,1754
=|1754,1755
=|1755,1756
=|1756,1757
=|1757,1758
=|1758,1759
=|1759,1760
=|1760,1761
=|1761,1762
=|1762,1763
=|1763,1764
=|1764,1765
=|1765,1766
=|1766,1767
=|1767,1768
=|1768,1769
=|1769,1770
=|1770,1771
=|1771,1772
=|1772,1773
=|1773,1774
=|1774,1775
=|1775,1776
=|1776,1777
=|1777,1778
<EOL>|1778,1779
VITALS|1779,1785
:|1785,1786
_|1787,1788
_|1788,1789
_|1789,1790
1136|1791,1795
Temp|1796,1800
:|1800,1801
98.1|1802,1806
PO|1807,1809
BP|1810,1812
:|1812,1813
107|1814,1817
/|1817,1818
68|1818,1820
R|1821,1822
lying|1823,1828
HR|1829,1831
:|1831,1832
68|1833,1835
<EOL>|1836,1837
RR|1837,1839
:|1839,1840
18|1841,1843
O2|1844,1846
<EOL>|1846,1847
sat|1847,1850
:|1850,1851
100|1852,1855
%|1855,1856
O2|1857,1859
delivery|1860,1868
:|1868,1869
RA|1870,1872
<EOL>|1874,1875
GENERAL|1875,1882
:|1882,1883
NAD|1885,1888
,|1888,1889
sitting|1890,1897
up|1898,1900
in|1901,1903
chair|1904,1909
,|1909,1910
smiling|1911,1918
,|1918,1919
moving|1920,1926
head|1927,1931
around|1932,1938
<EOL>|1938,1939
EYES|1939,1943
:|1943,1944
Sclera|1945,1951
anicteric|1952,1961
and|1962,1965
without|1966,1973
injection|1974,1983
.|1983,1984
<EOL>|1985,1986
CARDIAC|1986,1993
:|1993,1994
RRR|1995,1998
.|1998,1999
Audible|2000,2007
S1|2008,2010
and|2011,2014
S2|2015,2017
.|2017,2018
No|2019,2021
murmurs|2022,2029
/|2029,2030
rubs|2030,2034
/|2034,2035
gallops|2035,2042
.|2042,2043
<EOL>|2043,2044
RESP|2044,2048
:|2048,2049
Clear|2050,2055
to|2056,2058
auscultation|2059,2071
bilaterally|2072,2083
.|2083,2084
No|2085,2087
wheezes|2088,2095
,|2095,2096
rhonchi|2097,2104
or|2105,2107
<EOL>|2107,2108
rales|2108,2113
.|2113,2114
No|2115,2117
increased|2118,2127
work|2128,2132
of|2133,2135
breathing|2136,2145
.|2145,2146
<EOL>|2146,2147
ABDOMEN|2147,2154
:|2154,2155
Normal|2156,2162
bowels|2163,2169
sounds|2170,2176
,|2176,2177
non|2178,2181
distended|2182,2191
,|2191,2192
non-tender|2193,2203
.|2203,2204
<EOL>|2204,2205
EXTREMITIES|2205,2216
:|2216,2217
Pulses|2218,2224
DP|2225,2227
/|2227,2228
Radial|2228,2234
2|2235,2236
+|2236,2237
bilaterally|2238,2249
.|2249,2250
<EOL>|2250,2251
SKIN|2251,2255
:|2255,2256
Warm|2257,2261
.|2261,2262
Cap|2263,2266
refill|2267,2273
<|2274,2275
2s|2275,2277
.|2277,2278
No|2279,2281
rash|2282,2286
.|2286,2287
<EOL>|2287,2288
NEUROLOGIC|2288,2298
:|2298,2299
Speech|2300,2306
slow|2307,2311
but|2312,2315
markedly|2316,2324
improved|2325,2333
today|2334,2339
and|2340,2343
speaks|2344,2350
<EOL>|2351,2352
in|2352,2354
simple|2355,2361
<EOL>|2361,2362
sentences|2362,2371
.|2371,2372
Sitting|2373,2380
in|2381,2383
a|2384,2385
chair|2386,2391
and|2392,2395
able|2396,2400
to|2401,2403
move|2404,2408
all|2409,2412
extremities|2413,2424
,|2424,2425
<EOL>|2426,2427
follow|2427,2433
commands|2434,2442
such|2443,2447
as|2448,2450
moving|2451,2457
fingers|2458,2465
/|2465,2466
toes|2466,2470
on|2471,2473
command|2474,2481
and|2482,2485
<EOL>|2486,2487
sticking|2487,2495
thumb|2496,2501
up|2502,2504
.|2504,2505
<EOL>|2505,2506
PSYCH|2506,2511
:|2511,2512
Alert|2513,2518
and|2519,2522
awake|2523,2528
,|2528,2529
pleasant|2530,2538
,|2538,2539
smiling|2540,2547
<EOL>|2548,2549
<EOL>|2549,2550
<EOL>|2551,2552
Brief|2552,2557
Hospital|2558,2566
Course|2567,2573
:|2573,2574
<EOL>|2574,2575
BRIEF|2575,2580
HOSPITAL|2581,2589
SUMMARY|2590,2597
:|2597,2598
<EOL>|2598,2599
=|2599,2600
=|2600,2601
=|2601,2602
=|2602,2603
=|2603,2604
=|2604,2605
=|2605,2606
=|2606,2607
=|2607,2608
=|2608,2609
=|2609,2610
=|2610,2611
=|2611,2612
=|2612,2613
=|2613,2614
=|2614,2615
=|2615,2616
=|2616,2617
=|2617,2618
=|2618,2619
=|2619,2620
=|2620,2621
=|2621,2622
<EOL>|2622,2623
_|2623,2624
_|2624,2625
_|2625,2626
female|2627,2633
with|2634,2638
history|2639,2646
of|2647,2649
disordered|2650,2660
eating|2661,2667
,|2667,2668
PTSD|2669,2673
,|2673,2674
GAD|2675,2678
<EOL>|2679,2680
with|2680,2684
panic|2685,2690
disorder|2691,2699
,|2699,2700
depression|2701,2711
and|2712,2715
functional|2716,2726
neurological|2727,2739
<EOL>|2740,2741
disorder|2741,2749
presenting|2750,2760
from|2761,2765
a|2766,2767
therapy|2768,2775
session|2776,2783
with|2784,2788
weakness|2789,2797
,|2797,2798
<EOL>|2799,2800
abnormal|2800,2808
movement|2809,2817
,|2817,2818
and|2819,2822
aphasia|2823,2830
concerning|2831,2841
for|2842,2845
an|2846,2848
acute|2849,2854
<EOL>|2855,2856
functional|2856,2866
neurological|2867,2879
episode|2880,2887
.|2887,2888
She|2889,2892
was|2893,2896
evaluated|2897,2906
by|2907,2909
neurology|2910,2919
<EOL>|2920,2921
and|2921,2924
psychology|2925,2935
who|2936,2939
felt|2940,2944
this|2945,2949
was|2950,2953
consistent|2954,2964
with|2965,2969
functional|2970,2980
<EOL>|2981,2982
neurological|2982,2994
disorder|2995,3003
,|3003,3004
similar|3005,3012
to|3013,3015
her|3016,3019
prior|3020,3025
presentation|3026,3038
.|3038,3039
She|3040,3043
<EOL>|3044,3045
began|3045,3050
working|3051,3058
with|3059,3063
_|3064,3065
_|3065,3066
_|3066,3067
and|3068,3071
OT|3072,3074
and|3075,3078
had|3079,3082
made|3083,3087
great|3088,3093
improvement|3094,3105
at|3106,3108
<EOL>|3109,3110
time|3110,3114
of|3115,3117
discharge|3118,3127
to|3128,3130
acute|3131,3136
rehab|3137,3142
.|3142,3143
<EOL>|3144,3145
<EOL>|3145,3146
TRANSITIONAL|3146,3158
ISSUES|3159,3165
:|3165,3166
<EOL>|3166,3167
=|3167,3168
=|3168,3169
=|3169,3170
=|3170,3171
=|3171,3172
=|3172,3173
=|3173,3174
=|3174,3175
=|3175,3176
=|3176,3177
=|3177,3178
=|3178,3179
=|3179,3180
=|3180,3181
=|3181,3182
=|3182,3183
=|3183,3184
=|3184,3185
=|3185,3186
=|3186,3187
<EOL>|3187,3188
For|3188,3191
rehab|3192,3197
:|3197,3198
<EOL>|3198,3199
[|3199,3200
]|3200,3201
Please|3202,3208
continue|3209,3217
aggressive|3218,3228
_|3229,3230
_|3230,3231
_|3231,3232
and|3233,3236
OT|3237,3239
for|3240,3243
further|3244,3251
improvement|3252,3263
<EOL>|3264,3265
in|3265,3267
functional|3268,3278
status|3279,3285
.|3285,3286
<EOL>|3287,3288
[|3288,3289
]|3289,3290
On|3291,3293
discharge|3294,3303
,|3303,3304
please|3305,3311
ensure|3312,3318
patient|3319,3326
has|3327,3330
follow|3331,3337
up|3338,3340
with|3341,3345
her|3346,3349
<EOL>|3350,3351
PCP|3351,3354
and|3355,3358
her|3359,3362
therapist|3363,3372
.|3372,3373
<EOL>|3374,3375
[|3375,3376
]|3376,3377
Patient|3378,3385
was|3386,3389
having|3390,3396
some|3397,3401
intermittent|3402,3414
nausea|3415,3421
as|3422,3424
appetite|3425,3433
<EOL>|3434,3435
improved|3435,3443
.|3443,3444
Please|3445,3451
continue|3452,3460
Zofran|3461,3467
TID|3468,3471
prn|3472,3475
.|3475,3476
QTc|3477,3480
was|3481,3484
441|3485,3488
on|3489,3491
EKG|3492,3495
on|3496,3498
<EOL>|3499,3500
_|3500,3501
_|3501,3502
_|3502,3503
.|3503,3504
If|3505,3507
continuing|3508,3518
Zofran|3519,3525
use|3526,3529
for|3530,3533
>|3534,3535
1|3535,3536
week|3537,3541
,|3541,3542
please|3543,3549
recheck|3550,3557
QTc|3558,3561
<EOL>|3562,3563
on|3563,3565
_|3566,3567
_|3567,3568
_|3568,3569
and|3570,3573
d|3574,3575
/|3575,3576
c|3576,3577
medication|3578,3588
if|3589,3591
prolonged|3592,3601
.|3601,3602
<EOL>|3602,3603
[|3603,3604
]|3604,3605
Patient|3606,3613
has|3614,3617
a|3618,3619
history|3620,3627
of|3628,3630
disordered|3631,3641
and|3642,3645
restrictive|3646,3657
eating|3658,3664
.|3664,3665
<EOL>|3666,3667
She|3667,3670
does|3671,3675
well|3676,3680
eating|3681,3687
with|3688,3692
encouragement|3693,3706
and|3707,3710
did|3711,3714
not|3715,3718
show|3719,3723
any|3724,3727
<EOL>|3728,3729
evidence|3729,3737
of|3738,3740
eating|3741,3747
disorder|3748,3756
while|3757,3762
inpatient|3763,3772
.|3772,3773
Please|3774,3780
continue|3781,3789
<EOL>|3790,3791
ensure|3791,3797
supplements|3798,3809
TID|3810,3813
with|3814,3818
meals|3819,3824
.|3824,3825
<EOL>|3826,3827
<EOL>|3827,3828
For|3828,3831
PCP|3832,3835
/|3835,3836
therapist|3836,3845
:|3845,3846
<EOL>|3846,3847
[|3847,3848
]|3848,3849
Please|3850,3856
refer|3857,3862
patient|3863,3870
to|3871,3873
psychiatrist|3874,3886
for|3887,3890
further|3891,3898
titration|3899,3908
of|3909,3911
<EOL>|3912,3913
psychiatric|3913,3924
medications|3925,3936
,|3936,3937
given|3938,3943
report|3944,3950
of|3951,3953
previous|3954,3962
sensitivity|3963,3974
to|3975,3977
<EOL>|3978,3979
medications|3979,3990
and|3991,3994
concern|3995,4002
for|4003,4006
possible|4007,4015
bipolar|4016,4023
disorder|4024,4032
diagnosis|4033,4042
.|4042,4043
<EOL>|4044,4045
<EOL>|4045,4046
[|4046,4047
]|4047,4048
Please|4049,4055
follow|4056,4062
up|4063,4065
pending|4066,4073
thiamine|4074,4082
level|4083,4088
.|4088,4089
<EOL>|4090,4091
<EOL>|4091,4092
ACUTE|4092,4097
ISSUES|4098,4104
:|4104,4105
<EOL>|4105,4106
=|4106,4107
=|4107,4108
=|4108,4109
=|4109,4110
=|4110,4111
=|4111,4112
=|4112,4113
=|4113,4114
=|4114,4115
=|4115,4116
=|4116,4117
=|4117,4118
=|4118,4119
<EOL>|4119,4120
#|4120,4121
GAD|4122,4125
/|4125,4126
Panic|4126,4131
disorder|4132,4140
<EOL>|4140,4141
#|4141,4142
Depression|4143,4153
<EOL>|4153,4154
#|4154,4155
PTSD|4156,4160
<EOL>|4160,4161
#|4161,4162
Functional|4163,4173
neurological|4174,4186
disorder|4187,4195
<EOL>|4195,4196
Patient|4196,4203
presented|4204,4213
from|4214,4218
a|4219,4220
therapy|4221,4228
session|4229,4236
where|4237,4242
she|4243,4246
had|4247,4250
acute|4251,4256
<EOL>|4257,4258
onset|4258,4263
of|4264,4266
weakness|4267,4275
,|4275,4276
abnormal|4277,4285
movement|4286,4294
and|4295,4298
aphasia|4299,4306
in|4307,4309
the|4310,4313
setting|4314,4321
<EOL>|4322,4323
of|4323,4325
potential|4326,4335
trigger|4336,4343
of|4344,4346
seeing|4347,4353
shadows|4354,4361
outside|4362,4369
the|4370,4373
door|4374,4378
.|4378,4379
Per|4380,4383
her|4384,4387
<EOL>|4388,4389
therapist|4389,4398
,|4398,4399
over|4400,4404
the|4405,4408
past|4409,4413
several|4414,4421
weeks|4422,4427
she|4428,4431
has|4432,4435
been|4436,4440
increasingly|4441,4453
<EOL>|4454,4455
more|4455,4459
hypervigilant|4460,4473
and|4474,4477
stressed|4478,4486
about|4487,4492
going|4493,4498
home|4499,4503
for|4504,4507
the|4508,4511
<EOL>|4512,4513
holidays|4513,4521
to|4522,4524
see|4525,4528
her|4529,4532
mom|4533,4536
,|4536,4537
which|4538,4543
is|4544,4546
a|4547,4548
major|4549,4554
trigger|4555,4562
for|4563,4566
her|4567,4570
PTSD|4571,4575
.|4575,4576
<EOL>|4577,4578
Her|4578,4581
therapist|4582,4591
also|4592,4596
reports|4597,4604
a|4605,4606
history|4607,4614
of|4615,4617
sexual|4618,4624
/|4624,4625
physical|4625,4633
/|4633,4634
verbal|4634,4640
<EOL>|4641,4642
abuse|4642,4647
but|4648,4651
patient|4652,4659
is|4660,4662
very|4663,4667
guarded|4668,4675
about|4676,4681
it|4682,4684
and|4685,4688
will|4689,4693
not|4694,4697
discuss|4698,4705
<EOL>|4706,4707
it|4707,4709
.|4709,4710
On|4711,4713
presentation|4714,4726
to|4727,4729
the|4730,4733
_|4734,4735
_|4735,4736
_|4736,4737
had|4738,4741
significant|4742,4753
and|4754,4757
acute|4758,4763
<EOL>|4764,4765
functional|4765,4775
neurological|4776,4788
symptoms|4789,4797
,|4797,4798
including|4799,4808
weakness|4809,4817
,|4817,4818
abnormal|4819,4827
<EOL>|4828,4829
movement|4829,4837
,|4837,4838
and|4839,4842
aphasia|4843,4850
,|4850,4851
resulting|4852,4861
in|4862,4864
impaired|4865,4873
functioning|4874,4885
.|4885,4886
There|4887,4892
<EOL>|4893,4894
was|4894,4897
concern|4898,4905
for|4906,4909
catatonia|4910,4919
and|4920,4923
she|4924,4927
improved|4928,4936
after|4937,4942
1|4943,4944
mg|4945,4947
IV|4948,4950
ativan|4951,4957
<EOL>|4958,4959
in|4959,4961
the|4962,4965
ER|4966,4968
.|4968,4969
She|4970,4973
endorsed|4974,4982
significant|4983,4994
anxiety|4995,5002
,|5002,5003
but|5004,5007
denied|5008,5014
SI|5015,5017
and|5018,5021
,|5021,5022
<EOL>|5023,5024
per|5024,5027
Psychiatry|5028,5038
,|5038,5039
she|5040,5043
did|5044,5047
not|5048,5051
meet|5052,5056
_|5057,5058
_|5058,5059
_|5059,5060
criteria|5061,5069
.|5069,5070
She|5071,5074
had|5075,5078
a|5079,5080
<EOL>|5081,5082
similar|5082,5089
episode|5090,5097
in|5098,5100
_|5101,5102
_|5102,5103
_|5103,5104
after|5105,5110
IV|5111,5113
iron|5114,5118
infusion|5119,5127
and|5128,5131
was|5132,5135
<EOL>|5136,5137
admitted|5137,5145
to|5146,5148
the|5149,5152
neurology|5153,5162
service|5163,5170
,|5170,5171
where|5172,5177
she|5178,5181
was|5182,5185
diagnosed|5186,5195
with|5196,5200
<EOL>|5201,5202
functional|5202,5212
neurological|5213,5225
disorder|5226,5234
and|5235,5238
she|5239,5242
improved|5243,5251
with|5252,5256
_|5257,5258
_|5258,5259
_|5259,5260
and|5261,5264
<EOL>|5265,5266
rehab|5266,5271
.|5271,5272
She|5273,5276
was|5277,5280
also|5281,5285
started|5286,5293
on|5294,5296
nortriptyline|5297,5310
10|5311,5313
mg|5314,5316
QHS|5317,5320
at|5321,5323
that|5324,5328
<EOL>|5329,5330
time|5330,5334
.|5334,5335
Per|5336,5339
her|5340,5343
therapist|5344,5353
,|5353,5354
she|5355,5358
is|5359,5361
sensitive|5362,5371
to|5372,5374
medications|5375,5386
and|5387,5390
<EOL>|5391,5392
when|5392,5396
she|5397,5400
was|5401,5404
on|5405,5407
SSRIs|5408,5413
she|5414,5417
became|5418,5424
manic|5425,5430
,|5430,5431
although|5432,5440
she|5441,5444
has|5445,5448
not|5449,5452
<EOL>|5453,5454
formally|5454,5462
been|5463,5467
diagnosed|5468,5477
with|5478,5482
bipolar|5483,5490
disorder|5491,5499
.|5499,5500
Once|5501,5505
admitted|5506,5514
,|5514,5515
<EOL>|5516,5517
she|5517,5520
was|5521,5524
re-evaluated|5525,5537
by|5538,5540
neuro|5541,5546
and|5547,5550
psychiatry|5551,5561
who|5562,5565
determined|5566,5576
this|5577,5581
<EOL>|5582,5583
was|5583,5586
not|5587,5590
consistent|5591,5601
with|5602,5606
catatonia|5607,5616
and|5617,5620
instead|5621,5628
was|5629,5632
likely|5633,5639
<EOL>|5640,5641
functional|5641,5651
neurological|5652,5664
disorder|5665,5673
.|5673,5674
She|5675,5678
was|5679,5682
recommended|5683,5694
for|5695,5698
acute|5699,5704
<EOL>|5705,5706
rehab|5706,5711
to|5712,5714
continue|5715,5723
aggressive|5724,5734
_|5735,5736
_|5736,5737
_|5737,5738
.|5738,5739
She|5740,5743
was|5744,5747
continued|5748,5757
on|5758,5760
home|5761,5765
<EOL>|5766,5767
nortriptyline|5767,5780
10mg|5781,5785
qhs|5786,5789
.|5789,5790
<EOL>|5790,5791
<EOL>|5791,5792
#|5792,5793
Disordered|5793,5803
eating|5804,5810
<EOL>|5810,5811
#|5811,5812
Restrictive|5812,5823
eating|5824,5830
<EOL>|5830,5831
#|5831,5832
Over-exercising|5832,5847
<EOL>|5848,5849
She|5849,5852
has|5853,5856
a|5857,5858
history|5859,5866
of|5867,5869
restrictive|5870,5881
eating|5882,5888
and|5889,5892
over-exercising|5893,5908
and|5909,5912
<EOL>|5913,5914
in|5914,5916
the|5917,5920
past|5921,5925
she|5926,5929
has|5930,5933
had|5934,5937
bradycardia|5938,5949
and|5950,5953
electrolyte|5954,5965
<EOL>|5966,5967
abnormalities|5967,5980
.|5980,5981
Per|5982,5985
her|5986,5989
therapist|5990,5999
,|5999,6000
her|6001,6004
disordered|6005,6015
eating|6016,6022
has|6023,6026
<EOL>|6027,6028
become|6028,6034
much|6035,6039
worse|6040,6045
over|6046,6050
the|6051,6054
past|6055,6059
few|6060,6063
months|6064,6070
in|6071,6073
the|6074,6077
setting|6078,6085
of|6086,6088
<EOL>|6089,6090
traveling|6090,6099
a|6100,6101
lot|6102,6105
for|6106,6109
work|6110,6114
.|6114,6115
She|6116,6119
started|6120,6127
an|6128,6130
intensive|6131,6140
outpatient|6141,6151
<EOL>|6152,6153
program|6153,6160
at|6161,6163
_|6164,6165
_|6165,6166
_|6166,6167
Eating|6168,6174
_|6175,6176
_|6176,6177
_|6177,6178
on|6179,6181
_|6182,6183
_|6183,6184
_|6184,6185
.|6185,6186
Per|6187,6190
her|6191,6194
<EOL>|6195,6196
therapist|6196,6205
,|6205,6206
she|6207,6210
restricts|6211,6220
her|6221,6224
calories|6225,6233
to|6234,6236
about|6237,6242
1,000|6243,6248
or|6249,6251
less|6252,6256
a|6257,6258
<EOL>|6259,6260
day|6260,6263
and|6264,6267
over-exercises|6268,6282
and|6283,6286
is|6287,6289
good|6290,6294
at|6295,6297
hiding|6298,6304
it|6305,6307
from|6308,6312
people|6313,6319
.|6319,6320
<EOL>|6321,6322
From|6322,6326
review|6327,6333
of|6334,6336
OMR|6337,6340
,|6340,6341
her|6342,6345
BMI|6346,6349
seems|6350,6355
to|6356,6358
be|6359,6361
normal|6362,6368
(|6369,6370
between|6370,6377
_|6378,6379
_|6379,6380
_|6380,6381
<EOL>|6382,6383
and|6383,6386
she|6387,6390
currently|6391,6400
does|6401,6405
not|6406,6409
have|6410,6414
any|6415,6418
electrolyte|6419,6430
abnormalities|6431,6444
<EOL>|6445,6446
but|6446,6449
she|6450,6453
has|6454,6457
been|6458,6462
intermittently|6463,6477
bradycardic|6478,6489
with|6490,6494
HR|6495,6497
in|6498,6500
the|6501,6504
_|6505,6506
_|6506,6507
_|6507,6508
.|6508,6509
<EOL>|6510,6511
Her|6511,6514
appetite|6515,6523
improved|6524,6532
as|6533,6535
her|6536,6539
neurological|6540,6552
symptoms|6553,6561
began|6562,6567
<EOL>|6568,6569
resolving|6569,6578
.|6578,6579
Per|6580,6583
nutrition|6584,6593
evaluation|6594,6604
,|6604,6605
no|6606,6608
need|6609,6613
for|6614,6617
eating|6618,6624
disorder|6625,6633
<EOL>|6634,6635
protocol|6635,6643
while|6644,6649
inpatient|6650,6659
.|6659,6660
She|6661,6664
received|6665,6673
Ensure|6674,6680
supplements|6681,6692
.|6692,6693
Heart|6694,6699
<EOL>|6700,6701
rates|6701,6706
were|6707,6711
stable|6712,6718
,|6718,6719
bradycardic|6720,6731
in|6732,6734
_|6735,6736
_|6736,6737
_|6737,6738
.|6738,6739
Electrolytes|6740,6752
were|6753,6757
<EOL>|6758,6759
monitored|6759,6768
.|6768,6769
TSH|6770,6773
,|6773,6774
T4|6775,6777
and|6778,6781
B12|6782,6785
levels|6786,6792
were|6793,6797
all|6798,6801
normal|6802,6808
.|6808,6809
She|6810,6813
received|6814,6822
<EOL>|6823,6824
thiamine|6824,6832
supplementation|6833,6848
.|6848,6849
She|6850,6853
received|6854,6862
Zofran|6863,6869
PRN|6870,6873
for|6874,6877
nausea|6878,6884
<EOL>|6885,6886
(|6886,6887
QTc|6887,6890
441|6891,6894
)|6894,6895
.|6895,6896
<EOL>|6896,6897
<EOL>|6897,6898
CORE|6898,6902
MEASURES|6903,6911
<EOL>|6911,6912
=|6912,6913
=|6913,6914
=|6914,6915
=|6915,6916
=|6916,6917
=|6917,6918
=|6918,6919
=|6919,6920
=|6920,6921
=|6921,6922
=|6922,6923
=|6923,6924
=|6924,6925
<EOL>|6925,6926
#|6926,6927
CODE|6927,6931
:|6931,6932
full|6933,6937
code|6938,6942
<EOL>|6943,6944
#|6944,6945
CONTACT|6945,6952
:|6952,6953
Per|6954,6957
patient|6958,6965
's|6965,6967
request|6968,6975
,|6975,6976
do|6977,6979
not|6980,6983
contact|6984,6991
her|6992,6995
mother|6996,7002
<EOL>|7002,7003
(|7003,7004
_|7004,7005
_|7005,7006
_|7006,7007
)|7007,7008
<EOL>|7008,7009
-|7010,7011
Emergency|7011,7020
Contacts|7021,7029
:|7029,7030
_|7031,7032
_|7032,7033
_|7033,7034
(|7035,7036
_|7036,7037
_|7037,7038
_|7038,7039
)|7039,7040
_|7041,7042
_|7042,7043
_|7043,7044
and|7045,7048
_|7049,7050
_|7050,7051
_|7051,7052
(|7053,7054
Uncle|7054,7059
)|7059,7060
_|7061,7062
_|7062,7063
_|7063,7064
<EOL>|7065,7066
-|7067,7068
Therapist|7068,7077
:|7077,7078
_|7079,7080
_|7080,7081
_|7081,7082
,|7082,7083
_|7084,7085
_|7085,7086
_|7086,7087
_|7088,7089
_|7089,7090
_|7090,7091
and|7092,7095
coordinates|7096,7107
<EOL>|7107,7108
all|7108,7111
of|7112,7114
her|7115,7118
care|7119,7123
and|7124,7127
available|7128,7137
for|7138,7141
questions|7142,7151
/|7151,7152
calls|7152,7157
at|7158,7160
anytime|7161,7168
<EOL>|7168,7169
<EOL>|7169,7170
<EOL>|7171,7172
Medications|7172,7183
on|7184,7186
Admission|7187,7196
:|7196,7197
<EOL>|7197,7198
The|7198,7201
Preadmission|7202,7214
Medication|7215,7225
list|7226,7230
is|7231,7233
accurate|7234,7242
and|7243,7246
complete|7247,7255
.|7255,7256
<EOL>|7256,7257
1.|7257,7259
Nortriptyline|7260,7273
10|7274,7276
mg|7277,7279
PO|7280,7282
QHS|7283,7286
<EOL>|7287,7288
<EOL>|7288,7289
<EOL>|7290,7291
Discharge|7291,7300
Medications|7301,7312
:|7312,7313
<EOL>|7313,7314
1.|7314,7316
Multivitamins|7318,7331
W|7332,7333
/|7333,7334
minerals|7334,7342
1|7343,7344
TAB|7345,7348
PO|7349,7351
DAILY|7352,7357
<EOL>|7359,7360
2.|7360,7362
Ondansetron|7364,7375
ODT|7376,7379
4|7380,7381
mg|7382,7384
PO|7385,7387
Q8H|7388,7391
:|7391,7392
PRN|7392,7395
Nausea|7396,7402
/|7402,7403
Vomiting|7403,7411
-|7412,7413
First|7414,7419
Line|7420,7424
<EOL>|7425,7426
<EOL>|7427,7428
3.|7428,7430
Thiamine|7432,7440
100|7441,7444
mg|7445,7447
PO|7448,7450
DAILY|7451,7456
<EOL>|7458,7459
4.|7459,7461
Nortriptyline|7463,7476
10|7477,7479
mg|7480,7482
PO|7483,7485
QHS|7486,7489
<EOL>|7491,7492
<EOL>|7492,7493
<EOL>|7494,7495
Discharge|7495,7504
Disposition|7505,7516
:|7516,7517
<EOL>|7517,7518
Extended|7518,7526
Care|7527,7531
<EOL>|7531,7532
<EOL>|7533,7534
Facility|7534,7542
:|7542,7543
<EOL>|7543,7544
_|7544,7545
_|7545,7546
_|7546,7547
<EOL>|7547,7548
<EOL>|7549,7550
Discharge|7550,7559
Diagnosis|7560,7569
:|7569,7570
<EOL>|7570,7571
#|7571,7572
Functional|7572,7582
neurological|7583,7595
disorder|7596,7604
<EOL>|7604,7605
#|7605,7606
GAD|7606,7609
/|7609,7610
depression|7610,7620
<EOL>|7620,7621
#|7621,7622
PTSD|7622,7626
<EOL>|7626,7627
#|7627,7628
H|7628,7629
/|7629,7630
o|7630,7631
disordered|7632,7642
eating|7643,7649
<EOL>|7650,7651
<EOL>|7651,7652
<EOL>|7653,7654
Discharge|7654,7663
Condition|7664,7673
:|7673,7674
<EOL>|7674,7675
Mental|7675,7681
Status|7682,7688
:|7688,7689
Clear|7690,7695
and|7696,7699
coherent|7700,7708
.|7708,7709
<EOL>|7709,7710
Level|7710,7715
of|7716,7718
Consciousness|7719,7732
:|7732,7733
Alert|7734,7739
and|7740,7743
interactive|7744,7755
.|7755,7756
<EOL>|7756,7757
Activity|7757,7765
Status|7766,7772
:|7772,7773
Out|7774,7777
of|7778,7780
Bed|7781,7784
with|7785,7789
assistance|7790,7800
to|7801,7803
chair|7804,7809
or|7810,7812
<EOL>|7813,7814
wheelchair|7814,7824
.|7824,7825
<EOL>|7825,7826
<EOL>|7826,7827
<EOL>|7828,7829
Discharge|7829,7838
Instructions|7839,7851
:|7851,7852
<EOL>|7852,7853
Dear|7853,7857
Ms.|7858,7861
_|7862,7863
_|7863,7864
_|7864,7865
,|7865,7866
<EOL>|7866,7867
<EOL>|7867,7868
It|7868,7870
was|7871,7874
a|7875,7876
privilege|7877,7886
taking|7887,7893
care|7894,7898
of|7899,7901
you|7902,7905
at|7906,7908
_|7909,7910
_|7910,7911
_|7911,7912
<EOL>|7913,7914
_|7914,7915
_|7915,7916
_|7916,7917
.|7917,7918
<EOL>|7920,7921
<EOL>|7921,7922
WHY|7922,7925
WAS|7926,7929
I|7930,7931
ADMITTED|7932,7940
TO|7941,7943
THE|7944,7947
HOSPITAL|7948,7956
?|7956,7957
<EOL>|7957,7958
=|7958,7959
=|7959,7960
=|7960,7961
=|7961,7962
=|7962,7963
=|7963,7964
=|7964,7965
=|7965,7966
=|7966,7967
=|7967,7968
=|7968,7969
=|7969,7970
=|7970,7971
=|7971,7972
=|7972,7973
=|7973,7974
=|7974,7975
=|7975,7976
=|7976,7977
=|7977,7978
=|7978,7979
=|7979,7980
=|7980,7981
=|7981,7982
=|7982,7983
=|7983,7984
=|7984,7985
=|7985,7986
=|7986,7987
=|7987,7988
=|7988,7989
=|7989,7990
=|7990,7991
=|7991,7992
=|7992,7993
<EOL>|7993,7994
-|7994,7995
You|7995,7998
came|7999,8003
to|8004,8006
the|8007,8010
hospital|8011,8019
because|8020,8027
you|8028,8031
acutely|8032,8039
had|8040,8043
trouble|8044,8051
moving|8052,8058
<EOL>|8059,8060
and|8060,8063
speaking|8064,8072
.|8072,8073
<EOL>|8074,8075
<EOL>|8075,8076
WHAT|8076,8080
HAPPENED|8081,8089
WHILE|8090,8095
I|8096,8097
WAS|8098,8101
IN|8102,8104
THE|8105,8108
HOSPITAL|8109,8117
?|8117,8118
<EOL>|8118,8119
=|8119,8120
=|8120,8121
=|8121,8122
=|8122,8123
=|8123,8124
=|8124,8125
=|8125,8126
=|8126,8127
=|8127,8128
=|8128,8129
=|8129,8130
=|8130,8131
=|8131,8132
=|8132,8133
=|8133,8134
=|8134,8135
=|8135,8136
=|8136,8137
=|8137,8138
=|8138,8139
=|8139,8140
=|8140,8141
=|8141,8142
=|8142,8143
=|8143,8144
=|8144,8145
=|8145,8146
=|8146,8147
=|8147,8148
=|8148,8149
=|8149,8150
=|8150,8151
=|8151,8152
=|8152,8153
=|8153,8154
=|8154,8155
=|8155,8156
=|8156,8157
=|8157,8158
=|8158,8159
=|8159,8160
=|8160,8161
<EOL>|8161,8162
-|8162,8163
You|8163,8166
were|8167,8171
seen|8172,8176
by|8177,8179
the|8180,8183
neurologists|8184,8196
who|8197,8200
diagnosed|8201,8210
you|8211,8214
with|8215,8219
<EOL>|8220,8221
functional|8221,8231
neurological|8232,8244
disorder|8245,8253
.|8253,8254
<EOL>|8255,8256
-|8256,8257
You|8257,8260
worked|8261,8267
with|8268,8272
physical|8273,8281
and|8282,8285
occupational|8286,8298
therapists|8299,8309
.|8309,8310
<EOL>|8310,8311
-|8311,8312
Your|8312,8316
symptoms|8317,8325
began|8326,8331
to|8332,8334
improve|8335,8342
.|8342,8343
<EOL>|8343,8344
<EOL>|8344,8345
WHAT|8345,8349
SHOULD|8350,8356
I|8357,8358
DO|8359,8361
AFTER|8362,8367
I|8368,8369
LEAVE|8370,8375
THE|8376,8379
HOSPITAL|8380,8388
?|8388,8389
<EOL>|8389,8390
=|8390,8391
=|8391,8392
=|8392,8393
=|8393,8394
=|8394,8395
=|8395,8396
=|8396,8397
=|8397,8398
=|8398,8399
=|8399,8400
=|8400,8401
=|8401,8402
=|8402,8403
=|8403,8404
=|8404,8405
=|8405,8406
=|8406,8407
=|8407,8408
=|8408,8409
=|8409,8410
=|8410,8411
=|8411,8412
=|8412,8413
=|8413,8414
=|8414,8415
=|8415,8416
=|8416,8417
=|8417,8418
=|8418,8419
=|8419,8420
=|8420,8421
=|8421,8422
=|8422,8423
=|8423,8424
=|8424,8425
=|8425,8426
=|8426,8427
=|8427,8428
=|8428,8429
=|8429,8430
=|8430,8431
=|8431,8432
=|8432,8433
=|8433,8434
<EOL>|8436,8437
-|8437,8438
Please|8439,8445
continue|8446,8454
to|8455,8457
take|8458,8462
all|8463,8466
your|8467,8471
medications|8472,8483
and|8484,8487
follow|8488,8494
up|8495,8497
<EOL>|8498,8499
with|8499,8503
your|8504,8508
doctors|8509,8516
at|8517,8519
your|8520,8524
_|8525,8526
_|8526,8527
_|8527,8528
appointments|8529,8541
.|8541,8542
<EOL>|8544,8545
-|8545,8546
Please|8547,8553
continue|8554,8562
to|8563,8565
work|8566,8570
with|8571,8575
your|8576,8580
physical|8581,8589
and|8590,8593
occupational|8594,8606
<EOL>|8607,8608
therapists|8608,8618
.|8618,8619
<EOL>|8619,8620
<EOL>|8620,8621
We|8621,8623
wish|8624,8628
you|8629,8632
all|8633,8636
the|8637,8640
best|8641,8645
!|8645,8646
<EOL>|8646,8647
<EOL>|8647,8648
Sincerely|8648,8657
,|8657,8658
<EOL>|8659,8660
<EOL>|8661,8662
Your|8662,8666
_|8667,8668
_|8668,8669
_|8669,8670
Care|8671,8675
Team|8676,8680
<EOL>|8682,8683
<EOL>|8684,8685
Followup|8685,8693
Instructions|8694,8706
:|8706,8707
<EOL>|8707,8708
_|8708,8709
_|8709,8710
_|8710,8711
<EOL>|8711,8712

