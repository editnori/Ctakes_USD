CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Pharmaceutical Preparations|Drug|false|false||Drugsnull|Drugs - dental services|Procedure|false|false||Drugsnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Poorly controlled|Finding|false|false||poorly controllednull|Bad|Modifier|false|false||poorlynull|Type 2|Finding|false|false||type 2null|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Diabetes Mellitus, Insulin-Dependent|Disorder|false|false||IDDMnull|Hypertensive disease|Disorder|false|false||HTNnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|Past Week|Time|false|false||past weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Jan.|Time|false|false||jannull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|Fatigue|Finding|false|false||fatiguednull|Hospital admission|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|Admitsnull|Radiation Ionizing Radiotherapy|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|radiation
null|Radiotherapy Research|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|radiation
null|Radiation therapy (procedure)|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|radiationnull|Electromagnetic Radiation|Phenomenon|false|false|C4048756;C0446516;C1140618;C1269078|radiation
null|Radiation|Phenomenon|false|false|C4048756;C0446516;C1140618;C1269078|radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Right arm|Anatomy|false|false|C1522449;C1524020;C1524021;C3495676;C1522541;C5400986;C4761640;C1824218;C3715044;C0034519;C0851346;C0184666|R armnull|Anorectal Malformations|Disorder|false|false|C4048756;C0446516;C1140618;C1269078|armnull|AKR1A1 wt Allele|Finding|false|false|C0446516;C1140618;C1269078;C4048756|arm
null|ARMC9 gene|Finding|false|false|C0446516;C1140618;C1269078;C4048756|armnull|Protocol Treatment Arm|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C4048756;C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C3495676;C1522449;C1524020;C1524021;C1824218;C3715044;C1522541;C5400986;C4761640;C0034519;C0851346;C0184666|arm
null|null|Anatomy|false|false|C3495676;C1522449;C1524020;C1524021;C1824218;C3715044;C1522541;C5400986;C4761640;C0034519;C0851346;C0184666|arm
null|Upper Extremity|Anatomy|false|false|C3495676;C1522449;C1524020;C1524021;C1824218;C3715044;C1522541;C5400986;C4761640;C0034519;C0851346;C0184666|armnull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Felt faint|Finding|false|false||felt faintnull|Faint - appearance|Finding|false|false||faint
null|Syncope|Finding|false|false||faintnull|Chest tightness|Finding|false|false|C1527391;C0817096|chest tightnessnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0232292|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0232292|chestnull|Tightness sensation quality|Modifier|false|false||tightnessnull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Associated with|Modifier|false|false||associatednull|Dyspnea|Finding|true|false||SOBnull|Increased sweating|Finding|true|false||Diaphoresisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Dyspnea|Finding|false|false||SOBnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Chest Pain|Finding|true|false|C1527391;C0817096|chest painnull|null|Attribute|true|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Dyspnea|Finding|true|false||SOBnull|Current (present time)|Time|false|false||currentlynull|All other|Finding|false|false||All othernull|Reactive Oxygen Species|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|Reactive Oxygen Species|Drug|false|false|C0262327|ROSnull|ROS1 wt Allele|Finding|false|false|C0262327|ROS
null|ROS1 gene|Finding|false|false|C0262327|ROSnull|Review of systems (procedure)|Procedure|false|false|C0262327|ROSnull|rostral sulcus|Anatomy|false|false|C0812281;C1709820;C0289313;C0162772;C0489633|ROSnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Asthma|Disorder|false|false||asthmanull|Pulmonary Emphysema|Disorder|false|false||emphysemanull|Pathological accumulation of air in tissues|Finding|false|false||emphysemanull|Bronchitis, Chronic|Disorder|false|false||chronic bronchitisnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Acute bronchitis|Disorder|false|false||bronchitis
null|Bronchitis|Disorder|false|false||bronchitisnull|Hypertensive disease|Disorder|false|false||HTNnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|null|Device|false|false||stentsnull|Migraine Disorders|Disorder|false|false||migrainesnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Pills|Drug|false|false||pillsnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Neuropathy|Disorder|false|false||neuropathynull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|parent|Subject|false|false||parentsnull|Daughter|Subject|false|false||daughternull|Hypertensive disease|Disorder|false|false||htnnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Male Gender|Finding|false|false||malenull|Male, Self-Reported|Subject|false|false||male
null|Males|Subject|false|false||malenull|Male Phenotype|Modifier|false|false||malenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0036412;C2228481;C0205180|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false|C0229274;C0009758|Conjunctiva
null|Conjunctival Diseases|Disorder|false|false|C0229274;C0009758|Conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false|C0229274;C0009758|Conjunctiva
null|null|Finding|false|false|C0229274;C0009758|Conjunctivanull|examination of conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctiva
null|Procedure on conjunctiva|Procedure|false|false|C0229274;C0009758|Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false|C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759|Conjunctiva
null|conjunctiva|Anatomy|false|false|C1550624;C1546576;C0872390;C2228431;C0153628;C0154025;C0009759|Conjunctivanull|Pink color|Modifier|false|false||pinknull|Pallor of skin|Finding|true|false|C0026724;C0026639|pallornull|Cyanosis|Finding|true|false|C0026724;C0026639|cyanosisnull|Oral mucous membrane structure|Anatomy|false|false|C1272919;C0010520;C1561514;C1527415;C4521986;C0241137|oral mucosanull|Oral Dosage Form|Drug|false|false|C0026639;C0026724;C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896;C0026639;C0026724|oral
null|Oral (intended site)|Finding|false|false|C0226896;C0026639;C0026724|oralnull|Oral cavity|Anatomy|false|false|C1561514;C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|null|Finding|false|false|C0226896;C0026639;C0026724|mucosanull|Mucous Membrane|Anatomy|false|false|C0010520;C1272919;C0241137;C1527415;C4521986;C1561514|mucosanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Jugular venous engorgement|Finding|true|false||JVDnull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C0741025|Chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|Chestnull|cetrimonium bromide|Drug|false|false||CTABnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C4037978;C0003483;C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055;C0869784|Abd
null|Abdomen|Anatomy|false|false|C3811055;C0869784|Abdnull|Procedure on aorta|Procedure|false|false|C4037978;C0003483;C0449202;C0000726|aortanull|Chest+Abdomen>Aorta|Anatomy|false|false|C3811055;C0869784|aorta
null|Aorta|Anatomy|false|false|C3811055;C0869784|aortanull|Palpation|Procedure|false|false||palpationnull|Bruit|Finding|true|false||bruitsnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Femur|Anatomy|false|false|C0006318|femoralnull|Bruit|Finding|true|false|C0015811|bruitsnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0178298;C0496955|Skinnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|false|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||Pulsesnull|Physiologic pulse|Finding|false|false||Pulsesnull|Pulse taking|Procedure|false|false||Pulsesnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Stress bismuth subsalicylate|Drug|false|false||Stress
null|Stress bismuth subsalicylate|Drug|false|false||Stressnull|Stress|Finding|false|false||Stressnull|W stress|Attribute|false|false||Stressnull|Interpretation Process|Finding|false|false||INTERPRETATIONnull|null|Attribute|false|false||INTERPRETATIONnull|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus, Insulin-Dependent|Disorder|false|false||IDDMnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|null|Device|false|false||stentnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C2926613;C1549543;C0030193;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C2926613;C1549543;C0030193;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|mg/kg/min|LabModifier|false|false||mg/kg/minnull|ug/g|LabModifier|false|false||mg/kgnull|kg/min|Finding|false|false||kg/minnull|Per Minute|Time|false|false||/minnull|Minangkabau Language|Entity|false|false||minnull|Minute of time|Time|false|false||minnull|Minimum|Modifier|false|false||minnull|Minute Unit of Plane Angle|LabModifier|false|false||min
null|minim|LabModifier|false|false||minnull|Persantine|Drug|false|false||persantine
null|Persantine|Drug|false|false||persantinenull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Inspiration (function)|Finding|false|false||inspirationnull|Symptoms|Finding|false|false||symptomnull|null|Attribute|false|false||symptomnull|null|Finding|false|false||aminophylline was givennull|aminophylline|Drug|false|false||aminophylline
null|aminophylline|Drug|false|false||aminophyllinenull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|ST segment|Finding|false|false||ST segmentnull|Anatomical segmentation|Modifier|false|false||segmentnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C1305231;C0030471|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0723346;C0016169|sinus
null|Nasal sinus|Anatomy|false|false|C0723346;C0016169|sinusnull|Hemodynamics|Finding|false|false||Hemodynamicnull|hemodynamics (procedure)|Procedure|false|false||Hemodynamicnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Appropriate|Modifier|false|false||appropriatenull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Possible|Finding|false|false||Possiblenull|Possible diagnosis|Modifier|false|false||Possible
null|Possibly Related to Intervention|Modifier|false|false||Possiblenull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Ischemic|Finding|false|false||ischemicnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Nuclear (incident type)|Modifier|false|false||Nuclear
null|Nuclear (nucleus)|Modifier|false|false||Nuclearnull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Myocardial perfusion|Subject|false|false||myocardial perfusionnull|Myocardium|Anatomy|false|false|C4281794;C4723760;C4721534;C0031001|myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Perfusion (biological)|Finding|false|false|C0027061|perfusion
null|Perfusion route|Finding|false|false|C0027061|perfusionnull|Chemotherapeutic Perfusion|Procedure|false|false|C0027061|perfusion
null|Perfusion (procedure)|Procedure|false|false|C0027061|perfusionnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Hypertensive disease|Disorder|false|false||HTNnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|Atypical chest pain|Finding|false|false|C1527391;C0817096|atypical chest painnull|atypia morphology|Finding|false|false||atypicalnull|Atypical|Modifier|false|false||atypicalnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0262384;C2926613;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0262384;C2926613;C0741025|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Poorly controlled|Finding|false|false||poorly controllednull|Bad|Modifier|false|false||poorlynull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Twi language|Entity|false|false||TWInull|Atypical Vascular Proliferation|Finding|false|false||AVLnull|Augmented Vector Left|Modifier|false|false||AVLnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|Numerous|LabModifier|false|false||multiplenull|Episode of|Time|false|false||episodesnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Exertion|Finding|false|false||exertionnull|Lacking|Modifier|false|false||lacknull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Rh Negative Blood Group|Finding|false|false|C0018787|negative
null|Negative|Finding|false|false|C0018787|negative
null|Negative Finding|Finding|false|false|C0018787|negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Cardiac enzymes|Drug|false|false|C0018787|cardiac enzymes
null|Cardiac enzymes|Drug|false|false|C0018787|cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false|C0018787|cardiac enzymesnull|null|Attribute|false|false|C0018787|cardiac enzymesnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C0443763;C0014445;C1314974;C2699077;C0205160;C1513916;C0201934;C2926589|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false|C0018787|enzymesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Nuclear (incident type)|Modifier|false|false||nuclear
null|Nuclear (nucleus)|Modifier|false|false||nuclearnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Patient Class - Inpatient|Finding|false|false||inpatient
null|Referral category - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Perfusion (biological)|Finding|false|false||perfusion
null|Perfusion route|Finding|false|false||perfusionnull|Chemotherapeutic Perfusion|Procedure|false|false||perfusion
null|Perfusion (procedure)|Procedure|false|false||perfusionnull|defects aspect|Finding|false|false||defectsnull|Continuous|Finding|false|false||Continuenull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|ACE protein, human|Drug|false|false||ACE
null|ACE protein, human|Drug|false|false||ACEnull|ACE gene|Finding|false|false||ACE
null|Adverse Childhood Experience questionnaire|Finding|false|false||ACEnull|cisplatin, cytarabine, and etoposide chemotherapy protocol|Procedure|false|false||ACE
null|cyclophosphamide/doxorubicin protocol|Procedure|false|false||ACE
null|CDE protocol|Procedure|false|false||ACE
null|CDE Regimen|Procedure|false|false||ACEnull|Achinese language|Entity|false|false||ACEnull|Continuous|Finding|false|false||Continuenull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||Statinnull|EEF1A2 gene|Finding|false|false||Statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||Statinnull|matrix metalloproteinase 7 activity|Finding|false|false||Pumpnull|null|Device|false|false||Pumpnull|Pump Dosing Unit|LabModifier|false|false||Pumpnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Rhythm|Finding|false|false||Rhythm
null|rhythmic process (biological)|Finding|false|false||Rhythmnull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|Hypertensive disease|Disorder|false|false||HTNnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Concern|Finding|false|false||Concernnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Compliance behavior|Finding|false|false||compliantnull|Compliant (qualifier value)|Modifier|false|false||compliantnull|Medication Regimen|Procedure|false|false||medication regimennull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Imdur|Drug|false|false||Imdur
null|Imdur|Drug|false|false||Imdurnull|Structure of subparietal sulcus|Anatomy|false|false||SBPsnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Titration Method|Procedure|false|false||titrationnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|Glycosylated hemoglobin A|Drug|false|false||HbA1c
null|Glycosylated hemoglobin A|Drug|false|false||HbA1cnull|Glucohemoglobin measurement|Procedure|false|false||HbA1cnull|Poorly controlled|Finding|false|false||Poorly controllednull|Bad|Modifier|false|false||Poorlynull|Current (present time)|Time|false|false||Currentlynull|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemirnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|metformin|Drug|false|false||Metformin
null|metformin|Drug|false|false||Metforminnull|three times a day at institution-specified times|Time|false|false||tid
null|Three times daily|Time|false|false||tidnull|Compliance behavior|Finding|true|false||compliantnull|Compliant (qualifier value)|Modifier|false|false||compliantnull|Continuous|Finding|false|false||Continuenull|metformin|Drug|false|false||metformin
null|metformin|Drug|false|false||metforminnull|Continuous|Finding|false|false||Continuenull|Lantus|Drug|false|false||Lantus
null|Lantus|Drug|false|false||Lantusnull|Every morning|Time|false|false||qAMnull|Once a day, at bedtime|Time|false|false||qHSnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Continuous|Finding|false|false||Continuenull|Lipitor|Drug|false|false||Lipitor
null|Lipitor|Drug|false|false||Lipitornull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Advair|Drug|false|false||Advair
null|Advair|Drug|false|false||Advairnull|Daily|Time|false|false||dailynull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|CIAO3 gene|Finding|false|false||prnnull|As required|Time|false|false||prn
null|Pro Re Nata|Time|false|false||prnnull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Daily|Time|false|false||dailynull|atenolol|Drug|false|false||Atenolol
null|atenolol|Drug|false|false||Atenololnull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||dailynull|metformin|Drug|false|false||Metformin
null|metformin|Drug|false|false||Metforminnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||dailynull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Daily|Time|false|false||dailynull|potassium chloride|Drug|false|false||Potassium chloride
null|potassium chloride|Drug|false|false||Potassium chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||chloride
null|Chlorides|Drug|false|false||chloridenull|Chloride metabolic function|Finding|false|false||chloridenull|Chloride measurement|Procedure|false|false||chloridenull|mEq|LabModifier|false|false||mEqnull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|fluticasone / salmeterol|Drug|false|false||Fluticasone-Salmeterolnull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|salmeterol|Drug|false|false||Salmeterol
null|salmeterol|Drug|false|false||Salmeterolnull|microgram|LabModifier|false|false||mcgnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C0034789;C0993608;C1550509|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329;C1556138|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Disk Drug Form|Drug|false|false|C1556138|Disknull|Disc - Body Part|Anatomy|false|false|C0993608;C1550509;C1561538;C1561539;C4546282;C0004048;C0205535;C1332410;C4035627|Disknull|Disk Device|Device|false|false||Disk
null|Disk - package|Device|false|false||Disknull|Disk Shape|Modifier|false|false||Disknull|Disk Dosing Unit|LabModifier|false|false||Disknull|Participation Type - device|Finding|false|false|C1556138|Devicenull|Medical Devices|Device|false|false||Device
null|Devices|Device|false|false||Devicenull|Kind of quantity - Device|LabModifier|false|false||Devicenull|Inhalation Route of Administration|Finding|false|false|C1556138|Inhalation
null|Inspiration (function)|Finding|false|false|C1556138|Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false|C1556138|BIDnull|BID gene|Finding|false|false|C1556138|BIDnull|Twice a day|Time|false|false||BIDnull|2 times|Finding|false|false|C1556138|2 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false|C1556138|day
null|Precision - day|Finding|false|false|C1556138|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|mcg/actuation|LabModifier|false|false||mcg/Actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||Actuationnull|Aerosol Dose Form|Drug|false|false||Aerosolnull|Aerosols|Device|false|false||Aerosolnull|Puff Dosing Unit|LabModifier|false|false||Puffsnull|Inhalation Route of Administration|Finding|false|false||Inhalation
null|Inspiration (function)|Finding|false|false||Inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||Inhalationnull|Every six hours|Time|false|false||Q6Hnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C1283071;C0391871;C0030685;C0680255;C1963578;C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C1283071;C0391871;C0030685;C0680255;C1963578;C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C1283071;C0391871;C0030685;C0680255;C1963578|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|acetaminophen / oxycodone|Drug|false|false||Oxycodone-Acetaminophennull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|Every six hours|Time|false|false||Q6Hnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemir
null|Levemir|Drug|false|false||Levemirnull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Solution Dosage Form|Drug|false|false||Solution
null|Solutions|Drug|false|false||Solution
null|Pharmaceutical Solutions|Drug|false|false||Solutionnull|Resolution|Finding|false|false||Solutionnull|Subcutaneous Route of Administration|Finding|false|false||Subcutaneousnull|subcutaneous|Modifier|false|false||Subcutaneousnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Every morning|Time|false|false||qAMnull|QPM|Time|false|false||qPM
null|Once a day, in the evening|Time|false|false||qPMnull|metformin|Drug|false|false||Metformin
null|metformin|Drug|false|false||Metforminnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false|C0524463;C1325531|Chloridenull|mEq|LabModifier|false|false||mEqnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935;C0201952;C0443318|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935;C0201952;C0443318|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Sustained Release Dosage Form|Drug|false|false||Sustained Releasenull|Sustained|Finding|false|false|C0524463;C1325531|Sustainednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C1561538;C1561539;C1720092;C0030685;C0680255;C1963578;C0006935;C1283071;C0391871|Capsule
null|Structure of organ capsule|Anatomy|false|false|C1561538;C1561539;C1720092;C0030685;C0680255;C1963578;C0006935;C1283071;C0391871|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Release - action (qualifier value)|Finding|false|false|C0524463;C1325531|Release
null|Released (action)|Finding|false|false|C0524463;C1325531|Releasenull|Discharge (release)|Procedure|false|false|C0524463;C1325531|Release
null|Release (procedure)|Procedure|false|false|C0524463;C1325531|Release
null|Patient Discharge|Procedure|false|false|C0524463;C1325531|Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false|C0524463;C1325531|oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false|C0524463;C1325531|day
null|Precision - day|Finding|false|false|C0524463;C1325531|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|Sublingual Tablet|Drug|false|false||Tablet, Sublingualnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Sig
null|Receptors, Antigen, B-Cell|Drug|false|false|C0262329|Signull|Receptors, Antigen, B-Cell|Finding|false|false|C0262329|Signull|Short insular gyrus|Anatomy|false|false|C0034789;C0034789|Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Sublingual Route of Administration|Finding|false|false||Sublingual
null|Sublingual (intended site)|Finding|false|false||Sublingualnull|Sublingual location|Modifier|false|false||Sublingualnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0741025;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Does sit|Finding|false|false||Sit
null|Sitting position|Finding|false|false||Sit
null|HHAT gene|Finding|false|false||Sit
null|SIT1 gene|Finding|false|false||Sitnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Tablet Dosage Form|Drug|false|false||tabnull|Tablet Dosing Unit|LabModifier|false|false||tabnull|5 minutes Office visit|Procedure|false|false||5 minutesnull|5 minutes|Time|false|false||5 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C1549543;C0030193;C2926613;C0008031;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C1549543;C0030193;C2926613;C0008031;C0741025|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMS
null|Ethyl Methanesulfonate|Drug|false|false||EMSnull|EMSLR gene|Finding|false|false||EMSnull|Emergency Medical Services|Procedure|false|false||EMSnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletsnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitrate
null|isosorbide mononitrate|Drug|false|false||Isosorbide Mononitratenull|isosorbide|Drug|false|false||Isosorbide
null|isosorbide|Drug|false|false||Isosorbidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Atypical chest pain|Finding|false|false|C1527391;C0817096|Atypical Chest painnull|atypia morphology|Finding|false|false|C1527391;C0817096|Atypicalnull|Atypical|Modifier|false|false||Atypicalnull|Chest Pain|Finding|false|false|C1527391;C0817096|Chest painnull|null|Attribute|false|false|C1527391;C0817096|Chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C2598155;C2926613;C0741025;C0008031;C0741302;C0262384;C1549543;C0030193|Chest
null|Anterior thoracic region|Anatomy|false|false|C2598155;C2926613;C0741025;C0008031;C0741302;C0262384;C1549543;C0030193|Chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false|C1527391;C0817096|painnull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|dependent|Finding|false|false||dependentnull|Dependent - ability|Modifier|false|false||dependent
null|Conditional|Modifier|false|false||dependentnull|Apyrexial|Finding|false|false||Afebrilenull|Chest Pain|Finding|false|false|C1527391;C0817096|Chest painnull|null|Attribute|false|false|C1527391;C0817096|Chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|Chestnull|Chest|Anatomy|false|false|C1547311;C0008031;C2926613;C0741025;C1549543;C0030193;C0332296|Chest
null|Anterior thoracic region|Anatomy|false|false|C1547311;C0008031;C2926613;C0741025;C1549543;C0030193;C0332296|Chestnull|Pain-Free|Drug|false|false||pain freenull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Free of (attribute)|Finding|false|false|C1527391;C0817096|freenull|Empty (qualifier)|Modifier|false|false||freenull|Patient Condition Code - Stable|Finding|false|false|C1527391;C0817096|stablenull|Stable status|Modifier|false|false||stablenull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C2926613|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Myocardial Infarction|Disorder|false|false|C4037974;C0018787|heart attacknull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C1304680;C1261512;C0027051;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C1304680;C1261512;C0027051;C0153957;C0153500|heartnull|Attack (finding)|Finding|false|false|C4037974;C0018787|attack
null|Attack behavior|Finding|false|false|C4037974;C0018787|attacknull|Attack device|Device|false|false||attacknull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0741025;C0008031;C1549543;C0030193|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0741025;C0008031;C1549543;C0030193|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Only a Little|Finding|false|false||a little
null|A little bit|Finding|false|false||a littlenull|Little's Disease|Disorder|false|false||littlenull|Only a Little|Finding|false|false||littlenull|Smallest|LabModifier|false|false||little
null|Small|LabModifier|false|false||littlenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Several|LabModifier|false|false||Severalnull|Dosage|LabModifier|false|false||dosesnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Imdur|Drug|false|false||imdur
null|Imdur|Drug|false|false||imdurnull|Daily|Time|false|false||dailynull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Daily|Time|false|false||dailynull|atenolol|Drug|false|false||atenolol
null|atenolol|Drug|false|false||atenololnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Exercise stress test|Procedure|false|false|C4318744|stress test
null|Stress Test|Procedure|false|false|C4318744|stress testnull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false|C4318744|stressnull|W stress|Attribute|false|false||stressnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0015260;C3494508;C0022885;C0038435;C0039593;C0392366;C0456984|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Follow|Finding|false|false||adhere tonull|Fix|Phenomenon|false|false||adherenull|Diet, Healthy|Finding|false|false||healthy dietnull|Healthy|Modifier|false|false||healthynull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Daily|Time|false|false||dailynull|Additional|Finding|false|false||additionalnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C2926613;C0741025;C0008031|chest
null|Anterior thoracic region|Anatomy|false|false|C2926613;C0741025;C0008031|chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Breath|Finding|false|false||breathnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||return tonull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions