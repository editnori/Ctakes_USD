CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|true|false||MEDICINEnull|Medicine|Title|true|false||MEDICINEnull|Known|Modifier|true|false||Knownnull|Hypersensitivity|Finding|true|false||Allergiesnull|null|Attribute|true|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|true|false||Drug
null|Pharmacologic Substance|Drug|true|false||Drugnull|Drug problem|Finding|true|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial|Modifier|false|false||superficialnull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Structure of left lower leg|Anatomy|false|false||lower Left legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false||Left leg numbnessnull|Structure of left lower leg|Anatomy|false|false||Left leg
null|Left lower extremity|Anatomy|false|false||Left legnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Numbness in leg|Finding|false|false||leg numbnessnull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Evening|Time|false|false||eveningnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Last|Modifier|false|false||lastnull|Night time|Time|false|false||nightnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Gradual|Modifier|false|false||gradualnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Muscle Cramp|Finding|false|false||crampingnull|Cramping sensation quality|Modifier|false|false||crampingnull|Lateral|Modifier|false|false||lateralnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|BORNHOLM EYE DISEASE|Disorder|true|false||bednull|Bachelor of Education|Finding|true|false||bednull|Beds|Device|true|false||bednull|Patient Location - Bed|Modifier|true|false||bednull|Exertion|Finding|true|false||exertionnull|Muscle Weakness Lower Limb|Finding|true|false||leg weakness
null|Monoparesis of lower limb|Finding|true|false||leg weaknessnull|Leg|Anatomy|true|false||leg
null|Lower Extremity|Anatomy|true|false||legnull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Able (qualifier value)|Finding|true|false||ablenull|Ability|Subject|true|false||ablenull|Helping Behavior|Finding|true|false||assistancenull|Assisted (qualifier value)|Modifier|true|false||assistancenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Residual|Modifier|false|false||residualnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Lateral|Modifier|false|false||lateralnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Spine Problem|Finding|true|false||spinenull|Neuron spine|Anatomy|true|false||spine
null|Vertebral column|Anatomy|true|false||spinenull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|true|false||traumanull|trauma qualifier|Modifier|true|false||traumanull|Back Pain|Finding|true|false||back painnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Incontinence|Disorder|true|false||incontinencenull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Headache|Finding|true|false||headachenull|Visual changes|Finding|true|false||visual changesnull|Visual|Finding|true|false||visualnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Chest Pain|Finding|false|false||pain, chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Chest pressure|Finding|false|false||chest pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Palpitations|Finding|false|false||palpitationsnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dysuria|Finding|false|false||dysurianull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Hypertensive disease|Disorder|false|false||hypertensionnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Cerebellum|Anatomy|false|false||cerebellarnull|Medullary - body parts|Anatomy|false|false||medullary
null|Medulla Oblongata|Anatomy|false|false||medullary
null|Adrenal Medulla|Anatomy|false|false||medullarynull|Cerebrovascular accident|Disorder|false|false||strokenull|Stroke (heart beat)|Finding|false|false||strokenull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Circumflex|Modifier|false|false||circumflexnull|Peripheral Arterial Diseases|Disorder|false|false||peripheral arterial disease
null|Peripheral Vascular Diseases|Disorder|false|false||peripheral arterial diseasenull|Peripheral|Modifier|false|false||peripheralnull|Arteriopathic disease|Disorder|false|false||arterial diseasenull|Arteries|Anatomy|false|false||arterialnull|Arterial|Modifier|false|false||arterialnull|Disease|Disorder|false|false||diseasenull|Intermittent Claudication|Disorder|false|false||claudicationnull|Claudication (finding)|Finding|false|false||claudication
null|Lameness|Finding|false|false||claudicationnull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Terminal esophageal web|Disorder|false|false||esophageal ringsnull|Esophageal Diseases|Disorder|false|false||esophagealnull|Esophageal|Modifier|false|false||esophagealnull|Ring device|Device|false|false||ringsnull|ring form of protozoa|Entity|false|false||ringsnull|Niece|Subject|false|false||Niecenull|Sorting - Cell Movement|Finding|false|false||sort
null|Sorting (Cognition)|Finding|false|false||sortnull|Sorting|Event|false|false||sortnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Lung diseases|Disorder|false|false||lung diseasenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Disease|Disorder|false|false||diseasenull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Early|Time|true|false||earlynull|DFFB protein, human|Drug|true|false||CAD
null|DFFB protein, human|Drug|true|false||CADnull|Cold Hemagglutinin Disease|Disorder|true|false||CAD
null|Coronary heart disease|Disorder|true|false||CAD
null|Coronary Artery Disease|Disorder|true|false||CADnull|CAD gene|Finding|true|false||CAD
null|CALD1 wt Allele|Finding|true|false||CAD
null|B4GALNT2 gene|Finding|true|false||CAD
null|DFFB wt Allele|Finding|true|false||CAD
null|ACOD1 gene|Finding|true|false||CAD
null|DFFB gene|Finding|true|false||CADnull|cytarabine/daunorubicin protocol|Procedure|true|false||CAD
null|Computer Assisted Diagnosis|Procedure|true|false||CAD
null|Collision-Induced Dissociation|Procedure|true|false||CAD
null|CyADIC regimen|Procedure|true|false||CADnull|Caddo language|Entity|true|false||CADnull|Sudden Cardiac Death|Finding|true|false||sudden cardiac deathnull|Sudden (qualifier value)|Modifier|true|false||suddennull|Cardiac Death|Finding|true|false||cardiac deathnull|Cardiac attachment|Finding|true|false||cardiacnull|Heart|Anatomy|true|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|true|false||cardiacnull|Event Consequence - Death|Finding|true|false||death
null|Death (finding)|Finding|true|false||death
null|Cessation of life|Finding|true|false||deathnull|Known|Modifier|true|false||knownnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|true|false||historynull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|true|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Pleasant|Finding|false|false||Pleasantnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|true|false||Supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|true|false||rhythm
null|rhythmic process (biological)|Finding|true|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Minimal|Modifier|false|false||Minimal
null|Mild (qualifier value)|Modifier|false|false||Minimal
null|Minimum|Modifier|false|false||Minimalnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Obese abdomen|Finding|false|false||obese abdomennull|Obesity|Disorder|false|false||obesenull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|true|false||softnull|Soft|Modifier|true|false||softnull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Posterior part of right leg|Anatomy|false|false||right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Swollen calf|Finding|false|false||calf swellingnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Greater|LabModifier|false|false||greaternull|Posterior part of left leg|Anatomy|false|false||left calfnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swollen calf|Finding|false|false||calf swellingnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|CALF TENDERNESS|Finding|true|false||calf tendernessnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Palpation|Procedure|true|false||palpationnull|Thick|Modifier|false|false||Thicknull|Structure of nail of toe|Anatomy|false|false||toenailsnull|Dry Skin brand of emollient|Drug|false|false||dry skinnull|Xeroderma|Disorder|false|false||dry skinnull|Dry skin|Finding|false|false||dry skinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|Congenital hallux valgus|Disorder|false|false||Hallux valgus
null|Hallux Valgus|Disorder|false|false||Hallux valgus
null|Acquired hallux valgus|Disorder|false|false||Hallux valgusnull|Hallux structure|Anatomy|false|false||Halluxnull|Valgus deformity|Disorder|false|false||valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|physical examination (physical finding)|Finding|false|false||PHYSICAL EXAMnull|Physical Examination|Procedure|false|false||PHYSICAL EXAMnull|physical examination (physical finding)|Finding|false|false||PHYSICAL
null|Physical|Finding|false|false||PHYSICALnull|Physical Examination|Procedure|false|false||PHYSICALnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Tmax|LabModifier|false|false||Tmaxnull|Saturation of Peripheral Oxygen|Attribute|false|false||SpO2null|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Pleasant|Finding|false|false||Pleasantnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Passive joint movement of neck (finding)|Finding|false|false||Neck
null|Neck problem|Finding|false|false||Necknull|dendritic spine neck|Anatomy|false|false||Neck
null|Neck|Anatomy|false|false||Necknull|Supple|Finding|true|false||Supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|true|false||rhythm
null|rhythmic process (biological)|Finding|true|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|true|false||clear
null|Transparent (qualitative concept)|Modifier|true|false||clearnull|Auscultation|Procedure|true|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Malignant neoplasm of abdomen|Disorder|true|false||Abdomennull|Abdomen problem|Finding|true|false||Abdomennull|Abdomen|Anatomy|true|false||Abdomen
null|Abdominal Cavity|Anatomy|true|false||Abdomennull|Obese abdomen|Finding|false|false||obese abdomennull|Obesity|Disorder|false|false||obesenull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|true|false||softnull|Soft|Modifier|true|false||softnull|Protective muscle spasm|Finding|true|false||guardingnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|null|Finding|false|false||radial pulsenull|examination of radial pulses|Procedure|false|false||radial pulsenull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Pulse Wave Normal|Finding|false|false||pulse 2+null|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|null|Finding|false|false||radial pulsenull|examination of radial pulses|Procedure|false|false||radial pulsenull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Pulse Wave Decreased|Finding|false|false||pulse 1+null|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Posterior part of right leg|Anatomy|false|false||right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Swollen calf|Finding|false|false||calf swellingnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Posterior part of left leg|Anatomy|false|false||left calfnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Swollen calf|Finding|false|false||calf swellingnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|CALF TENDERNESS|Finding|true|false||calf tendernessnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Palpation|Procedure|true|false||palpationnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Palpation|Procedure|true|false||palpationnull|Table Cell Horizontal Align - left|Finding|true|false||leftnull|Left sided|Modifier|true|false||left
null|Left|Modifier|true|false||leftnull|Dorsal|Modifier|true|false||dorsalnull|Lateral|Modifier|false|false||lateralnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Skin callus|Disorder|false|false||callousnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Lateral to the left|Modifier|false|false||left lateralnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lateral|Modifier|false|false||lateralnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Thick toenails|Finding|false|false||Thick toenailsnull|Thick|Modifier|false|false||Thicknull|Structure of nail of toe|Anatomy|false|false||toenailsnull|Dry Skin brand of emollient|Drug|false|false||dry skinnull|Xeroderma|Disorder|false|false||dry skinnull|Dry skin|Finding|false|false||dry skinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|indurated|Finding|false|false||induratednull|Cone-Rod Dystrophy 2|Disorder|false|false||cordnull|Cord - Body Parts|Anatomy|false|false||cordnull|Cord Device|Device|false|false||cordnull|left antecubital fossa|Anatomy|false|false||left antecubital fossanull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital Fossa|Anatomy|false|false||antecubital fossanull|Antecubital|Anatomy|false|false||antecubitalnull|Fossa|Anatomy|false|false||fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Ruta graveolens preparation|Drug|false|false||RUE
null|Ruta graveolens preparation|Drug|false|false||RUEnull|Ruta graveolens|Entity|false|false||RUE
null|Ruta|Entity|false|false||RUEnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Flexor (Anatomical coordinate)|Anatomy|false|false||flexornull|Flexor <Diplocrepinae>|Entity|false|false||flexornull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Plantar (qualifier value)|Anatomy|false|false||plantar
null|Sole of Foot|Anatomy|false|false||plantarnull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Legal fine|Entity|false|false||finenull|Fine (qualifier value)|Modifier|false|false||finenull|Touch sensation|Finding|false|false||touch sensationnull|Touch sensation|Finding|false|false||touch
null|Touch Perception|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Laboratory test finding|Lab|false|false||LABSnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Packed red blood cells|Drug|false|false||pRBCs
null|Packed red blood cells|Drug|false|false||pRBCsnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Coffee ground vomiting|Finding|false|false||coffee ground emesis
null|Vomit contains coffee grounds (finding)|Finding|false|false||coffee ground emesisnull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Doppler studies|Procedure|false|false||dopplernull|Deep Vein Thrombosis|Disorder|false|false||Deep venous thrombosisnull|Deep Resection Margin|Attribute|false|false||Deepnull|Deep (qualifier value)|Modifier|false|false||Deepnull|Venous thrombosis after immobility|Finding|false|false||venous thrombosis
null|Venous Thrombosis|Finding|false|false||venous thrombosisnull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Thrombosis|Finding|false|false||thrombosisnull|Bilateral|Modifier|false|false||bilateralnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false||tibialnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Right sided|Modifier|false|false||right-sidednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Small amount|LabModifier|true|false||Small amountnull|Small|LabModifier|true|false||Smallnull|Amount class - Amount|Finding|true|false||amountnull|Quantity|LabModifier|true|false||amountnull|Hematin|Drug|true|false||hematin
null|Hematin|Drug|true|false||hematinnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Ulceration|Finding|true|false||ulceration
null|Ulcer|Finding|true|false||ulcerationnull|Hemorrhage|Finding|true|false||bleedingnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Diffuse|Modifier|false|false||Diffusenull|Erythema|Disorder|false|false||erythemanull|Superficial|Modifier|false|false||superficialnull|Ulcer|Finding|false|false||ulcerationsnull|Carcinoma in situ of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Gastritis|Disorder|false|false||gastritisnull|Hemorrhage|Finding|true|false||bleedingnull|Medium (Substance)|Drug|false|false||Medium
null|Culture Media|Drug|false|false||Mediumnull|A Medium Amount of Time|Finding|false|false||Medium
null|Communications Media|Finding|false|false||Medium
null|A Medium Amount|Finding|false|false||Mediumnull|Message Waiting Priority - Medium|Modifier|false|false||Medium
null|medium exposure|Modifier|false|false||Mediumnull|Medium|LabModifier|false|false||Mediumnull|Hiatal Hernia|Disorder|false|false||hiatal hernianull|Hernia|Disorder|false|false||hernianull|Erythema|Disorder|false|false||Erythemanull|Superficial|Modifier|false|false||superficialnull|Ulcer|Finding|false|false||ulcerationsnull|Duodenal ampulla|Anatomy|false|false||duodenal bulbnull|Duodenum|Anatomy|false|false||duodenalnull|anatomical bulb|Anatomy|false|false||bulb
null|Medulla Oblongata|Anatomy|false|false||bulbnull|plant bulb|Entity|false|false||bulbnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Duodenitis|Disorder|false|false||duodenitis
null|Acute Enteritis of the Mouse Intestinal Tract|Disorder|false|false||duodenitisnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|III (suffix)|Modifier|false|false||thirdnull|Third|LabModifier|false|false||thirdnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Malignant neoplasm of duodenum|Disorder|false|false||duodenum
null|Benign neoplasm of duodenum|Disorder|false|false||duodenumnull|Duodenum|Anatomy|false|false||duodenumnull|Left upper extremity|Anatomy|false|false||Left upper extremitynull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Upper Extremity|Anatomy|false|false||upper extremitynull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Limb structure|Anatomy|false|false||extremitynull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Deep vein thrombosis of lower limb|Disorder|true|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|true|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|true|false||deep veinnull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|true|false||deepnull|Venous Thrombosis|Finding|true|false||vein thrombosisnull|Veins|Anatomy|true|false||veinnull|Thrombosis|Finding|true|false||thrombosisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Limb structure|Anatomy|false|false||extremitynull|Probable diagnosis|Finding|false|false||Likely
null|Probably|Finding|false|false||Likelynull|Evolving|Finding|false|false||evolvingnull|Hematoma|Finding|false|false||hematomanull|left antecubital fossa|Anatomy|false|false||left antecubital fossanull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital Fossa|Anatomy|false|false||antecubital fossanull|Antecubital|Anatomy|false|false||antecubitalnull|Fossa|Anatomy|false|false||fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|CAT scan of head|Procedure|false|false||CT headnull|null|Attribute|false|false||CT headnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Infarction|Finding|true|false||infarctionnull|Hemorrhage|Finding|true|false||hemorrhagenull|Fracture|Disorder|false|false||fracturesnull|Fractured|Finding|false|false||fracturesnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|edetic acid|Drug|false|false||EDTA
null|edetic acid|Drug|false|false||EDTAnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|Provider|Finding|false|false||Providersnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial|Modifier|false|false||superficialnull|Lower extremity>Femoral artery|Anatomy|false|false||femoral artery
null|Structure of femoral artery|Anatomy|false|false||femoral arterynull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Structure of left lower leg|Anatomy|false|false||lower left legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false||left leg numbnessnull|Structure of left lower leg|Anatomy|false|false||left leg
null|Left lower extremity|Anatomy|false|false||left legnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Numbness in leg|Finding|false|false||leg numbnessnull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Bilateral|Modifier|false|false||bilateralnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Hemorrhage|Finding|false|false||bleedingnull|Event|Event|false|false||eventsnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||blood
null|In Blood|Finding|true|false||bloodnull|Rectal Dosage Form|Drug|true|false||rectalnull|Rectal Route of Administration|Finding|true|false||rectal
null|Rectal (intended site)|Finding|true|false||rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|true|false||rectalnull|rectal|Modifier|true|false||rectalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Left upper arm structure|Anatomy|false|false||left arm
null|Left arm|Anatomy|false|false||left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Hematoma|Finding|false|false||hematomanull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Hematoma|Finding|false|false||hematomanull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Diagnostic Service Section ID - Hematology|Finding|false|false||Hematologynull|diagnostic service sources hematology (procedure)|Procedure|false|false||Hematology
null|Hematology procedure|Procedure|false|false||Hematology
null|Hematologic Tests|Procedure|false|false||Hematologynull|hematology (field)|Title|false|false||Hematologynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Left upper arm structure|Anatomy|false|false||left arm
null|Left arm|Anatomy|false|false||left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Hematoma|Finding|false|false||hematomanull|Slow|Modifier|false|false||slowlynull|Recommendation|Finding|false|false||recommendationsnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Rehabilitation therapy|Procedure|false|false||rehabnull|More|LabModifier|false|false||morenull|Problem|Finding|false|false||problemnull|null|Attribute|false|false||problemnull|summary - ActRelationshipSubset|Finding|false|false||summary
null|Summary (document)|Finding|false|false||summarynull|Marketing basis - Transitional|Finding|false|false||transitionalnull|Transitional cell morphology|Modifier|false|false||transitionalnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Peripheral Vascular Diseases|Disorder|false|false||PVDnull|Pomalidomide/Bortezomib/Dexamethasone Regimen|Procedure|false|false||PVDnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Superficial femoral artery|Anatomy|false|false||superficial femoral arterynull|Superficial|Modifier|false|false||superficialnull|Lower extremity>Femoral artery|Anatomy|false|false||femoral artery
null|Structure of femoral artery|Anatomy|false|false||femoral arterynull|Femur|Anatomy|false|false||femoralnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Structure of left lower leg|Anatomy|false|false||lower Left legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|numbness of left leg|Finding|false|false||Left leg numbnessnull|Structure of left lower leg|Anatomy|false|false||Left leg
null|Left lower extremity|Anatomy|false|false||Left legnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Numbness in leg|Finding|false|false||leg numbnessnull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Numbness|Finding|false|false||numbness
null|Hypesthesia|Finding|false|false||numbnessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Evening|Time|false|false||eveningnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Bilateral|Modifier|false|false||bilateralnull|Structure of posterior tibial vein|Anatomy|false|false||posterior tibial veinsnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Tibial vein structure|Anatomy|false|false||tibial veinsnull|Bone structure of tibia|Anatomy|false|false||tibialnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Bilateral|Modifier|false|false||Bilateralnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Clinical NEC (not elsewhere classified in LNC)|Finding|true|false||clinicalnull|Clinical|Modifier|true|false||clinicalnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Admission activity|Procedure|true|false||admission
null|Hospital admission|Procedure|true|false||admissionnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Bilateral|Modifier|false|false||bilateralnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Therapeutic brand of coal tar|Drug|false|false||therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||therapeutic
null|Therapeutic|Finding|false|false||therapeuticnull|Therapeutic procedure|Procedure|false|false||therapeuticnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Coagulation tissue factor induced.INR goal|Attribute|false|false||INR goalnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Due to|Finding|false|false||Due
null|Due|Finding|false|false||Duenull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Diagnostic Service Section ID - Hematology|Finding|true|false||hematologynull|diagnostic service sources hematology (procedure)|Procedure|true|false||hematology
null|Hematology procedure|Procedure|true|false||hematology
null|Hematologic Tests|Procedure|true|false||hematologynull|hematology (field)|Title|true|false||hematologynull|Further|Modifier|true|false||furthernull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Cardiologists|Subject|false|false||cardiologistnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Appropriate|Modifier|false|false||appropriatenull|Screening for cancer|Procedure|false|false||cancer screeningnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|Screening for cancer|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|research subject screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Encounter due to Screening for malignant neoplasm of breast|Finding|false|false||mammogramnull|Mammography|Procedure|false|false||mammogramnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|3 Months|Time|false|false||3 monthsnull|month|Time|false|false||monthsnull|Upper gastrointestinal hemorrhage|Finding|false|false||Upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||Upper GInull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Episode of|Time|false|false||episodenull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Coffee|Drug|false|false||coffeenull|Coffea <Coffeeae>|Entity|false|false||coffeenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Packed red blood cells|Drug|false|false||pRBCs
null|Packed red blood cells|Drug|false|false||pRBCsnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Gastritis|Disorder|false|false||gastritisnull|Superficial|Modifier|false|false||superficialnull|Superficial ulcer|Disorder|false|false||erosionsnull|Erosion lesion|Finding|false|false||erosionsnull|Hemorrhage|Finding|true|false||bleedingnull|Incidental Findings|Finding|false|false||Incidental findingnull|Incidental|Finding|false|false||Incidentalnull|Experimental Finding|Finding|false|false||finding
null|Signs and Symptoms|Finding|false|false||finding
null|Finding|Finding|false|false||findingnull|Medium (Substance)|Drug|false|false||medium
null|Culture Media|Drug|false|false||mediumnull|A Medium Amount of Time|Finding|false|false||medium
null|Communications Media|Finding|false|false||medium
null|A Medium Amount|Finding|false|false||mediumnull|Message Waiting Priority - Medium|Modifier|false|false||medium
null|medium exposure|Modifier|false|false||mediumnull|Medium|LabModifier|false|false||mediumnull|Hiatal Hernia|Disorder|false|false||hiatal hernianull|Hernia|Disorder|false|false||hernianull|Feces|Finding|false|false||Stoolnull|Stool seat|Device|false|false||Stoolnull|Antigens|Drug|false|false||antigennull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|week|Time|false|false||weeksnull|High dose|LabModifier|false|false||high dosenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Antecubital|Anatomy|false|false||antecubitalnull|Hematoma|Finding|false|false||hematomanull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Antecubital|Anatomy|false|false||antecubitalnull|Hematoma|Finding|false|false||hematomanull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|diagnostic service sources phlebotomy|Finding|false|false||phlebotomynull|Phlebotomy, therapeutic (separate procedure)|Procedure|false|false||phlebotomy
null|Venous blood sampling|Procedure|false|false||phlebotomy
null|Venesection|Procedure|false|false||phlebotomynull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin, porcine|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparin
null|heparin|Drug|false|false||Heparinnull|Hematoma|Finding|false|false||hematomanull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Stage level 4|Finding|false|false||Stage IVnull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Initially|Time|false|false||initiallynull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Daily|Time|false|false||dailynull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Has patient|Finding|false|false||Patient hasnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Rectal examination|Procedure|false|false||Rectal examnull|Rectal Dosage Form|Drug|false|false||Rectalnull|Rectal Route of Administration|Finding|false|false||Rectal
null|Rectal (intended site)|Finding|false|false||Rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||Rectalnull|rectal|Modifier|false|false||Rectalnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|EPO protein, human|Drug|false|false||EPO
null|epoetin alfa|Drug|false|false||EPO
null|epoetin alfa|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|Erythropoietin|Drug|false|false||EPO
null|EPO protein, human|Drug|false|false||EPOnull|EPO gene|Finding|false|false||EPO
null|TIMP1 wt Allele|Finding|false|false||EPO
null|EPX gene|Finding|false|false||EPO
null|TIMP1 gene|Finding|false|false||EPO
null|Exclusive Provider Organization Plan|Finding|false|false||EPOnull|Esperanto Language|Entity|false|false||EPOnull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|Adverse Event Probably Related to Intervention|Modifier|false|false||likely relatednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Slow|Modifier|false|false||slownull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Gastritis|Disorder|false|false||gastritisnull|Duodenitis|Disorder|false|false||duodenitis
null|Acute Enteritis of the Mouse Intestinal Tract|Disorder|false|false||duodenitisnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Hemorrhage|Finding|true|false||bleedingnull|iron studies|Procedure|false|false||Iron studiesnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Scientific Study|Procedure|false|false||studiesnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|BID protein, human|Drug|false|false||bid
null|BID protein, human|Drug|false|false||bidnull|Body integrity dysphoria|Disorder|false|false||bidnull|BID gene|Finding|false|false||bidnull|Twice a day|Time|false|false||bidnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Daily|Time|false|false||dailynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Circumflex|Modifier|false|false||circumflexnull|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Disorder|false|false||Pernull|Per - dosing instruction fragment|Finding|false|false||Per
null|PER1 gene|Finding|false|false||Per
null|Follow|Finding|false|false||Per
null|PER1 wt Allele|Finding|false|false||Pernull|PER (body structure)|Anatomy|false|false||Pernull|Per (qualifier)|Modifier|false|false||Pernull|Discussion (procedure)|Procedure|false|false||discussionsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cardiologists|Subject|false|false||cardiologistnull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Initially|Time|false|false||initiallynull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Daily|Time|false|false||dailynull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|Hypertensive disease|Disorder|false|false||HTNnull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Numerous|LabModifier|false|false||multiplenull|Bleeding episodes|Finding|false|false||bleeding episodesnull|Hemorrhage|Finding|false|false||bleedingnull|Episode of|Time|false|false||episodesnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|carvedilol|Drug|false|false||carvedilol
null|carvedilol|Drug|false|false||carvedilolnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Daily|Time|false|false||dailynull|Acute hemorrhage|Finding|false|false||acute bleednull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hemorrhage|Finding|false|false||bleednull|Structure of subparietal sulcus|Anatomy|false|false||SBPsnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Daily|Time|false|false||dailynull|Daily|Time|false|false||dailynull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Bedtime (qualifier value)|Time|false|false||bedtime
null|Once a day, at bedtime|Time|false|false||bedtimenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Screening - procedure intent|Finding|false|false||screening
null|Special screening finding|Finding|false|false||screening
null|Aspects of disease screening|Finding|false|false||screeningnull|research subject screening|Procedure|false|false||screening
null|Disease Screening|Procedure|false|false||screening
null|Screening|Procedure|false|false||screening
null|Screening for cancer|Procedure|false|false||screening
null|Screening procedure|Procedure|false|false||screeningnull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|Last|Modifier|false|false||lastnull|Encounter due to Screening for malignant neoplasm of breast|Finding|false|false||mammogramnull|Mammography|Procedure|false|false||mammogramnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Course|Time|false|false||coursenull|High dose|LabModifier|false|false||high dosenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|End date|Time|false|false||end datenull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Gastritis|Disorder|false|false||gastritisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|hypertensive agents|Drug|false|false||hypertension medicationsnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Daily|Time|false|false||dailynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|nifedipine|Drug|false|false||nifedipine
null|nifedipine|Drug|false|false||nifedipinenull|Daily|Time|false|false||dailynull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Hemorrhage|Finding|false|false||bleednull|Structure of subparietal sulcus|Anatomy|false|false||SBPsnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Cardiovascular system|Anatomy|false|false||cardiologynull|cardiology (field)|Title|false|false||cardiologynull|Cardiology service|Entity|false|false||cardiologynull|Arylsulfatase A, human|Drug|false|false||ASA
null|Arylsulfatase A, human|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASA
null|aspirin|Drug|false|false||ASAnull|ARSA gene|Finding|false|false||ASAnull|MDF Attribute Type - Address|Finding|false|false||address
null|Address (property)|Finding|false|false||address
null|Address|Finding|false|false||address
null|Value type - Address|Finding|false|false||address
null|Addresses (publication format)|Finding|false|false||address
null|Address Data Type|Finding|false|false||addressnull|null|Attribute|false|false||addressnull|Patient's home|Device|false|false||patient's homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|home environment (history)|Finding|false|false||home environmentnull|Home environment|Modifier|false|false||home environmentnull|Address type - Home|Finding|false|false||home
null|Visit User Code - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Home environment|Modifier|false|false||home
null|Person location type - Home|Modifier|false|false||homenull|Environment|Modifier|false|false||environmentnull|At increased risk for falls|Finding|false|false||fall risknull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Risk|Finding|false|false||risknull|Recent|Time|false|false||recentnull|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||trip
null|triptorelin|Drug|false|false||tripnull|TRAIP wt Allele|Finding|false|false||trip
null|TRAIP gene|Finding|false|false||trip
null|PIK3IP1 gene|Finding|false|false||trip
null|LRRFIP1 gene|Finding|false|false||tripnull|Tripping|Phenomenon|false|false||tripnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Class - Outpatient|Finding|false|false||outpatient
null|Referral category - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Rehabilitation therapy|Procedure|false|false||rehabnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|ranitidine|Drug|false|false||Ranitidine
null|ranitidine|Drug|false|false||Ranitidinenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Reflux|Finding|false|false||refluxnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Dinner|Finding|false|false||Dinnernull|With dinner|Time|false|false||Dinnernull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|allopurinol|Drug|false|false||Allopurinol
null|allopurinol|Drug|false|false||Allopurinolnull|Transaction counts and value totals - day|Finding|false|false||DAY
null|Precision - day|Finding|false|false||DAYnull|Land Dayak Languages|Entity|false|false||DAYnull|day|Time|false|false||DAY
null|Daily|Time|false|false||DAYnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|carvedilol|Drug|false|false||Carvedilol
null|carvedilol|Drug|false|false||Carvedilolnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Dinner|Finding|false|false||Dinnernull|With dinner|Time|false|false||Dinnernull|lisinopril|Drug|false|false||Lisinopril
null|lisinopril|Drug|false|false||Lisinoprilnull|Daily|Time|false|false||DAILYnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|nifedipine|Drug|false|false||NIFEdipine
null|nifedipine|Drug|false|false||NIFEdipinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|Neuropathic pain|Finding|false|false||neuropathic pain
null|Neuralgia|Finding|false|false||neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Every twelve hours|Time|false|false||Q12Hnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Constipation|Finding|false|false||constipationnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Deep Vein Thrombosis|Disorder|false|false||Deep vein thrombosis (DVT)null|Deep vein thrombosis of lower limb|Disorder|false|false||Deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||Deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||Deep veinnull|Deep Resection Margin|Attribute|false|false||Deepnull|Deep (qualifier value)|Modifier|false|false||Deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Deep Vein Thrombosis|Disorder|false|false||DVT
null|Deep thrombophlebitis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Upper gastrointestinal hemorrhage|Finding|false|false||Upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||Upper GInull|Upper Surface|Modifier|false|false||Upper
null|Upper|Modifier|false|false||Uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|Left arm|Anatomy|false|false||L armnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Hematoma|Finding|false|false||hematomanull|Superficial Thrombophlebitis|Disorder|false|false||Superficial thrombophlebitisnull|Superficial|Modifier|false|false||Superficialnull|Thrombophlebitis|Finding|false|false||thrombophlebitisnull|Antecubital Fossa|Anatomy|false|false||antecubital fossanull|Antecubital|Anatomy|false|false||antecubitalnull|Fossa|Anatomy|false|false||fossanull|Fossa <Euplerinae>|Entity|false|false||fossa
null|Cryptoprocta ferox|Entity|false|false||fossanull|Chronic Kidney Diseases|Disorder|false|false||Chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Kidney Diseases|Disorder|false|false||kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Disease|Disorder|false|false||diseasenull|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Peripheral Vascular Diseases|Disorder|false|false||Peripheral vascular diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false||vascular diseasenull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Disease|Disorder|false|false||diseasenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes mellitus type IInull|Diabetes Mellitus|Disorder|false|false||Diabetes mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Coronary Artery Disease|Disorder|false|false||Coronary artery disease
null|Coronary Arteriosclerosis|Disorder|false|false||Coronary artery diseasenull|Coronary artery|Anatomy|false|false||Coronary arterynull|Heart|Anatomy|false|false||Coronarynull|Coronary|Modifier|false|false||Coronarynull|Arteriopathic disease|Disorder|false|false||artery diseasenull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Disease|Disorder|false|false||diseasenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Swelling of lower limb|Finding|false|false||leg swellingnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Diagnostic tests|Procedure|false|false||Diagnostic testsnull|diagnostic tests device|Device|false|false||Diagnostic testsnull|Diagnostic agents|Drug|false|false||Diagnosticnull|Location Service Code - Diagnostic|Finding|false|false||Diagnostic
null|Diagnostic|Finding|false|false||Diagnosticnull|Diagnostic dental procedure|Procedure|false|false||Diagnostic
null|Diagnosis|Procedure|false|false||Diagnosticnull|Tests (qualifier value)|Finding|false|false||testsnull|Laboratory Procedures|Procedure|false|false||testsnull|Deep vein thrombosis of lower limb|Disorder|false|false||deep vein thrombosis
null|Deep Vein Thrombosis|Disorder|false|false||deep vein thrombosisnull|Structure of deep vein|Anatomy|false|false||deep veinnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Venous Thrombosis|Finding|false|false||vein thrombosisnull|Veins|Anatomy|false|false||veinnull|Thrombosis|Finding|false|false||thrombosisnull|Blood Clot|Finding|false|false||blood clots
null|Thrombus|Finding|false|false||blood clotsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Blood Clot|Finding|false|false||clotsnull|Leg|Anatomy|false|false||legsnull|null|Attribute|false|false||legsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Thinning Weight Loss|Finding|false|false||thinningnull|Decreased thickness|Modifier|false|false||thinningnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleedingnull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleedingnull|Hemorrhage|Finding|false|false||bleedingnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Left upper arm structure|Anatomy|false|false||left arm
null|Left arm|Anatomy|false|false||left armnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Hematoma|Finding|false|false||hematomanull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Own|Finding|false|false||ownnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Blood Clot|Finding|false|false||blood clots
null|Thrombus|Finding|false|false||blood clotsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Blood Clot|Finding|false|false||clotsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Upper gastrointestinal hemorrhage|Finding|false|false||upper GI bleednull|Upper gastrointestinal tract series|Procedure|false|false||upper GInull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Gastrointestinal Hemorrhage|Finding|false|false||GI bleednull|Hemorrhage|Finding|false|false||bleednull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|week|Time|false|false||weeksnull|clopidogrel|Drug|true|false||Clopidogrel
null|clopidogrel|Drug|true|false||Clopidogrelnull|Plavix|Drug|true|false||Plavix
null|Plavix|Drug|true|false||Plavixnull|Cardiologists|Subject|false|false||cardiologistnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions