 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Event|Event|Allergies|244,253|false|false|false|||Attending
Finding|Functional Concept|Allergies|244,253|false|false|false|C1999232|Attending (action)|Attending
Disorder|Disease or Syndrome|Chief Complaint|279,288|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|Chief Complaint|279,288|false|false|false|||Pneumonia
Event|Event|Chief Complaint|289,299|false|false|false|||identified
Finding|Classification|Chief Complaint|303,313|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Chief Complaint|303,313|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Chief Complaint|314,317|false|false|false|||CXR
Procedure|Diagnostic Procedure|Chief Complaint|314,317|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Classification|Chief Complaint|321,326|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|327,335|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|327,335|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|339,357|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|348,357|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|348,357|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|348,357|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|348,357|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|348,357|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|History of Present Illness|399,402|true|false|false|||PMH
Finding|Finding|History of Present Illness|399,402|true|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|History of Present Illness|406,412|false|false|false|C0004096|Asthma|Asthma
Event|Event|History of Present Illness|406,412|false|false|false|||Asthma
Disorder|Disease or Syndrome|History of Present Illness|414,418|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|414,418|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|414,418|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|414,418|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Hazardous or Poisonous Substance|History of Present Illness|420,427|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Immunologic Factor|History of Present Illness|420,427|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Organic Chemical|History of Present Illness|420,427|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Pharmacologic Substance|History of Present Illness|420,427|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Attribute|Clinical Attribute|History of Present Illness|420,431|false|false|false|C4522050||tobacco use
Finding|Finding|History of Present Illness|420,431|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Finding|Individual Behavior|History of Present Illness|420,431|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Event|Event|History of Present Illness|428,431|false|false|false|||use
Finding|Functional Concept|History of Present Illness|428,431|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|History of Present Illness|428,431|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|History of Present Illness|440,444|false|false|false|||days
Disorder|Disease or Syndrome|History of Present Illness|449,453|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|History of Present Illness|449,453|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|History of Present Illness|449,453|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|History of Present Illness|449,453|false|false|false|||cold
Finding|Organism Function|History of Present Illness|449,453|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|History of Present Illness|449,453|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|449,453|false|false|false|C0010412|Cold Therapy|cold
Event|Event|History of Present Illness|461,469|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|461,469|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|461,469|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|474,479|false|false|false|||noted
Finding|Intellectual Product|History of Present Illness|495,502|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|495,502|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Sign or Symptom|History of Present Illness|495,508|false|false|false|C0010201|Chronic Cough|chronic cough
Drug|Organic Chemical|History of Present Illness|503,508|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|503,508|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|503,508|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|503,508|false|false|false|C0010200|Coughing|cough
Drug|Biomedical or Dental Material|History of Present Illness|512,520|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|512,520|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|512,520|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|523,528|false|false|false|||worse
Finding|Finding|History of Present Illness|523,528|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|History of Present Illness|523,528|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Event|Event|History of Present Illness|543,548|false|false|false|||noted
Drug|Organic Chemical|History of Present Illness|558,563|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|558,563|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|558,563|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|558,563|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|572,582|false|false|false|||productive
Event|Event|History of Present Illness|591,597|false|false|false|||sputum
Finding|Body Substance|History of Present Illness|591,597|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|History of Present Illness|591,597|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|History of Present Illness|610,618|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|610,618|false|false|false|C0043144|Wheezing|wheezing
Attribute|Clinical Attribute|History of Present Illness|623,633|false|false|false|C2979880||subjective
Finding|Finding|History of Present Illness|623,633|false|false|false|C2266644|subjective (symptom)|subjective
Event|Event|History of Present Illness|634,640|false|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|634,640|false|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|655,659|true|false|false|||take
Event|Event|History of Present Illness|664,675|true|false|false|||temperature
Procedure|Health Care Activity|History of Present Illness|664,675|true|false|false|C0886414|Body temperature measurement|temperature
Event|Event|History of Present Illness|686,691|false|false|false|||noted
Drug|Biomedical or Dental Material|History of Present Illness|697,705|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|697,705|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|697,705|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|706,709|false|false|false|||DOE
Finding|Sign or Symptom|History of Present Illness|706,709|false|false|false|C0231807|Dyspnea on exertion|DOE
Event|Event|History of Present Illness|711,720|false|false|false|||increased
Finding|Intellectual Product|History of Present Illness|724,728|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|History of Present Illness|724,748|false|false|false|C4054523|Mildly Short of Breath|mild shortness of breath
Event|Event|History of Present Illness|729,738|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|729,748|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|729,748|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Finding|History of Present Illness|729,756|false|false|false|C0743330|Rest Dyspnea|shortness of breath at rest
Event|Event|History of Present Illness|742,748|false|false|false|||breath
Finding|Body Substance|History of Present Illness|742,748|false|false|false|C0225386|Breath|breath
Finding|Functional Concept|History of Present Illness|749,756|false|false|false|C0443144|At rest (qualifier value)|at rest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|752,756|false|false|false|C1742913|REST protein, human|rest
Drug|Biologically Active Substance|History of Present Illness|752,756|false|false|false|C1742913|REST protein, human|rest
Event|Event|History of Present Illness|752,756|false|false|false|||rest
Finding|Daily or Recreational Activity|History of Present Illness|752,756|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Gene or Genome|History of Present Illness|752,756|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Molecular Function|History of Present Illness|752,756|false|false|false|C0035253;C1419346;C1622890|REST gene;Rest;site-specific telomere resolvase activity|rest
Finding|Finding|History of Present Illness|774,778|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|774,778|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|774,778|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|779,785|false|false|false|||period
Finding|Organism Function|History of Present Illness|779,785|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|History of Present Illness|779,785|false|false|false|C2347804|Clinical Trial Period|period
Drug|Organic Chemical|History of Present Illness|795,802|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|History of Present Illness|795,802|false|false|false|C0699142|Tylenol|tylenol
Event|Event|History of Present Illness|795,802|false|false|false|||tylenol
Drug|Organic Chemical|History of Present Illness|807,817|false|false|false|C0723110|Robitussin|robitussin
Drug|Pharmacologic Substance|History of Present Illness|807,817|false|false|false|C0723110|Robitussin|robitussin
Event|Event|History of Present Illness|807,817|false|false|false|||robitussin
Finding|Idea or Concept|History of Present Illness|821,825|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Finding|History of Present Illness|821,832|false|false|false|C0541990|good effect|good effect
Event|Event|History of Present Illness|826,832|false|false|false|||effect
Event|Event|History of Present Illness|838,844|true|false|false|||denied
Event|Event|History of Present Illness|849,851|true|false|false|||CP
Event|Event|History of Present Illness|857,862|false|false|false|||noted
Event|Event|History of Present Illness|872,876|false|false|false|||felt
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|881,886|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|History of Present Illness|881,886|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|History of Present Illness|881,886|false|false|false|||heart
Finding|Sign or Symptom|History of Present Illness|881,886|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|History of Present Illness|888,895|false|false|false|||flutter
Finding|Pathologic Function|History of Present Illness|888,895|false|false|false|C0016385|Cardiac Flutter|flutter
Finding|Finding|History of Present Illness|910,914|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|910,914|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|910,914|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|915,921|false|false|false|||period
Finding|Organism Function|History of Present Illness|915,921|false|false|false|C0025344|Menstruation|period
Procedure|Research Activity|History of Present Illness|915,921|false|false|false|C2347804|Clinical Trial Period|period
Event|Event|History of Present Illness|926,933|true|false|false|||changed
Event|Event|History of Present Illness|950,959|true|false|false|||orthopnea
Finding|Finding|History of Present Illness|950,959|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|950,959|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|989,993|true|false|false|C0221423|Illness (finding)|sick
Event|Event|History of Present Illness|994,1002|true|false|false|||contacts
Procedure|Health Care Activity|History of Present Illness|994,1002|true|false|false|C4036459|Contacts|contacts
Event|Event|History of Present Illness|1007,1013|true|false|false|||denied
Event|Event|History of Present Illness|1019,1030|true|false|false|||association
Finding|Conceptual Entity|History of Present Illness|1019,1030|true|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Mental Process|History of Present Illness|1019,1030|true|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Social Behavior|History of Present Illness|1019,1030|true|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Phenomenon|Phenomenon or Process|History of Present Illness|1019,1030|true|false|false|C0596306|Chemical Association|association
Event|Event|History of Present Illness|1034,1042|true|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|1034,1042|true|false|false|C0018681|Headache|headache
Finding|Sign or Symptom|History of Present Illness|1044,1048|true|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|History of Present Illness|1044,1055|true|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|History of Present Illness|1044,1055|true|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|History of Present Illness|1044,1055|true|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|History of Present Illness|1044,1055|true|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|History of Present Illness|1049,1055|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1049,1055|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|History of Present Illness|1049,1055|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|History of Present Illness|1049,1055|false|false|false|||throat
Finding|Body Substance|History of Present Illness|1049,1055|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|History of Present Illness|1049,1055|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|History of Present Illness|1057,1065|false|false|false|||sneezing
Event|Event|History of Present Illness|1067,1077|false|false|false|||rhinorrhea
Finding|Sign or Symptom|History of Present Illness|1067,1077|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Attribute|Clinical Attribute|History of Present Illness|1080,1086|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1080,1086|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1080,1086|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1088,1096|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1088,1096|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1098,1106|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1098,1106|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1098,1106|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Anatomy|Body Location or Region|History of Present Illness|1108,1117|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1108,1122|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1118,1122|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1118,1122|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1118,1122|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1118,1122|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Gene or Genome|History of Present Illness|1147,1150|false|false|false|C1417080;C1537681|MCRS1 gene;MED25 gene|P78
Anatomy|Cell|History of Present Illness|1173,1176|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1173,1176|false|false|false|||WBC
Event|Event|History of Present Illness|1181,1187|false|false|false|||normal
Event|Event|History of Present Illness|1196,1201|false|false|false|||noted
Event|Event|History of Present Illness|1210,1218|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|1210,1218|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|1222,1226|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|1222,1226|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1222,1226|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|1232,1235|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1232,1235|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1240,1250|false|false|false|||suggestive
Finding|Functional Concept|History of Present Illness|1240,1250|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|History of Present Illness|1240,1253|false|false|false|C0332299|Suggestive of|suggestive of
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1254,1257|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|1259,1262|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|History of Present Illness|1259,1262|false|false|false|||PNA
Event|Event|History of Present Illness|1270,1275|false|false|false|||given
Drug|Organic Chemical|History of Present Illness|1282,1298|false|false|false|C4519262|Methylprednisone|methylprednisone
Drug|Pharmacologic Substance|History of Present Illness|1282,1298|false|false|false|C4519262|Methylprednisone|methylprednisone
Event|Event|History of Present Illness|1282,1298|false|false|false|||methylprednisone
Drug|Organic Chemical|History of Present Illness|1306,1314|false|false|false|C0721336|Levaquin|levaquin
Drug|Pharmacologic Substance|History of Present Illness|1306,1314|false|false|false|C0721336|Levaquin|levaquin
Event|Event|History of Present Illness|1306,1314|false|false|false|||levaquin
Drug|Biomedical or Dental Material|History of Present Illness|1327,1331|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|History of Present Illness|1327,1331|false|false|false|||nebs
Drug|Organic Chemical|History of Present Illness|1333,1342|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|History of Present Illness|1333,1342|false|false|false|C0001927|albuterol|albuterol
Event|Event|History of Present Illness|1333,1342|false|false|false|||albuterol
Event|Event|History of Present Illness|1356,1360|false|false|false|||CHEM
Finding|Functional Concept|History of Present Illness|1356,1360|false|false|false|C0079107|chemical aspects|CHEM
Procedure|Laboratory Procedure|History of Present Illness|1356,1360|false|false|false|C0201682|Chemical procedure|CHEM
Event|Event|History of Present Illness|1370,1378|false|false|false|||negative
Finding|Classification|History of Present Illness|1370,1378|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1370,1378|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1370,1378|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|1404,1412|false|false|false|||decision
Finding|Mental Process|History of Present Illness|1404,1412|false|false|false|C0679006|Decision|decision
Procedure|Health Care Activity|History of Present Illness|1425,1430|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admit
Event|Event|History of Present Illness|1456,1463|false|false|false|||therapy
Finding|Finding|History of Present Illness|1456,1463|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|History of Present Illness|1456,1463|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1456,1463|false|false|false|C0087111|Therapeutic procedure|therapy
Disorder|Disease or Syndrome|Past Medical History|1491,1497|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|Past Medical History|1491,1497|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1498,1502|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1498,1502|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1498,1502|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1498,1502|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Hazardous or Poisonous Substance|Past Medical History|1503,1510|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|Past Medical History|1503,1510|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|Past Medical History|1503,1510|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|Past Medical History|1503,1510|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Attribute|Clinical Attribute|Past Medical History|1503,1514|false|false|false|C4522050||Tobacco use
Finding|Finding|Past Medical History|1503,1514|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Finding|Individual Behavior|Past Medical History|1503,1514|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco use
Event|Event|Past Medical History|1511,1514|false|false|false|||use
Finding|Functional Concept|Past Medical History|1511,1514|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Past Medical History|1511,1514|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Disorder|Disease or Syndrome|Past Medical History|1515,1542|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|Peripheral Arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1526,1534|false|false|false|C0003842|Arteries|Arterial
Disorder|Disease or Syndrome|Past Medical History|1526,1542|false|false|false|C0852949|Arteriopathic disease|Arterial disease
Disorder|Disease or Syndrome|Past Medical History|1535,1542|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|1535,1542|false|false|false|||disease
Event|Event|Past Medical History|1554,1560|false|false|false|||common
Finding|Functional Concept|Past Medical History|1554,1560|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Past Medical History|1554,1560|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1561,1566|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1561,1575|false|false|false|C0850459|iliac stents|iliac stenting
Event|Event|Past Medical History|1567,1575|false|false|false|||stenting
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1567,1575|false|false|false|C2348535|Stenting|stenting
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1576,1582|false|false|false|C0018792|Heart Atrium|ATRIAL
Disorder|Disease or Syndrome|Past Medical History|1576,1594|false|false|false|C0546959|Atrial tachycardia|ATRIAL TACHYCARDIA
Finding|Finding|Past Medical History|1576,1594|false|false|false|C2059391|continuous electrocardiogram atrial tachycardia|ATRIAL TACHYCARDIA
Event|Event|Past Medical History|1583,1594|false|false|false|||TACHYCARDIA
Finding|Finding|Past Medical History|1583,1594|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|TACHYCARDIA
Finding|Finding|Past Medical History|1598,1606|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|1598,1617|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|1607,1612|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1607,1612|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|1607,1617|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|1607,1617|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|1613,1617|false|true|false|C2598155||PAIN
Event|Event|Past Medical History|1613,1617|false|false|false|||PAIN
Finding|Functional Concept|Past Medical History|1613,1617|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|1613,1617|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Anatomy|Body Location or Region|Past Medical History|1621,1629|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1621,1641|false|false|false|C0263884|Cervical radiculitis|CERVICAL RADICULITIS
Disorder|Disease or Syndrome|Past Medical History|1630,1641|false|false|false|C0034544|Radiculitis|RADICULITIS
Event|Event|Past Medical History|1630,1641|false|false|false|||RADICULITIS
Anatomy|Body Location or Region|Past Medical History|1645,1653|false|false|false|C0027530|Neck|CERVICAL
Disorder|Disease or Syndrome|Past Medical History|1645,1665|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|CERVICAL SPONDYLOSIS
Disorder|Disease or Syndrome|Past Medical History|1654,1665|false|false|false|C0038019|Spondylosis|SPONDYLOSIS
Event|Event|Past Medical History|1654,1665|false|false|false|||SPONDYLOSIS
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1669,1677|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1669,1684|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Past Medical History|1669,1692|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1678,1684|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|1678,1684|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|1678,1692|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Past Medical History|1685,1692|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|1685,1692|false|false|false|||DISEASE
Finding|Sign or Symptom|Past Medical History|1696,1704|false|false|false|C0018681|Headache|HEADACHE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1708,1711|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1708,1711|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|1708,1711|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|1708,1711|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|1708,1711|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|1708,1711|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1708,1711|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1708,1723|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|1712,1723|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|1712,1723|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|1712,1723|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1712,1723|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Disorder|Disease or Syndrome|Past Medical History|1727,1741|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|1727,1741|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|1727,1741|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Disorder|Disease or Syndrome|Past Medical History|1745,1757|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|1745,1757|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|1761,1775|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|1761,1775|false|false|false|||OSTEOARTHRITIS
Disorder|Disease or Syndrome|Past Medical History|1779,1785|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|HERPES
Disorder|Disease or Syndrome|Past Medical History|1779,1792|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Virus|Past Medical History|1779,1792|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|HERPES ZOSTER
Disorder|Disease or Syndrome|Past Medical History|1786,1792|false|false|false|C0019360|Herpes zoster (disorder)|ZOSTER
Event|Event|Past Medical History|1786,1792|false|false|false|||ZOSTER
Drug|Hazardous or Poisonous Substance|Past Medical History|1796,1803|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Past Medical History|1796,1803|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Past Medical History|1796,1803|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Past Medical History|1796,1803|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1796,1809|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1804,1809|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Past Medical History|1804,1809|false|false|false|||ABUSE
Event|Event|Past Medical History|1804,1809|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Past Medical History|1804,1809|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1813,1819|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Past Medical History|1813,1832|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|1813,1832|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Past Medical History|1813,1832|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|1820,1832|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|1820,1832|false|false|false|||FIBRILLATION
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1836,1843|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|ANXIETY
Event|Event|Past Medical History|1836,1843|false|false|false|||ANXIETY
Finding|Sign or Symptom|Past Medical History|1836,1843|false|false|false|C0860603|Anxiety symptoms|ANXIETY
Finding|Intellectual Product|Past Medical History|1848,1864|false|false|false|C1314977|Gastrointestinal attachment|GASTROINTESTINAL
Finding|Pathologic Function|Past Medical History|1848,1873|false|false|false|C0017181|Gastrointestinal Hemorrhage|GASTROINTESTINAL BLEEDING
Finding|Pathologic Function|Past Medical History|1865,1873|false|false|false|C0019080|Hemorrhage|BLEEDING
Disorder|Disease or Syndrome|Past Medical History|1877,1891|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|1877,1891|false|false|false|||OSTEOARTHRITIS
Finding|Functional Concept|Past Medical History|1895,1910|false|false|false|C0333482|atherosclerotic|ATHEROSCLEROTIC
Disorder|Disease or Syndrome|Past Medical History|1895,1933|false|false|false|C0004153|Atherosclerosis|ATHEROSCLEROTIC CARDIOVASCULAR DISEASE
Anatomy|Body System|Past Medical History|1911,1925|false|false|false|C0007226;C3887460|Cardiovascular;Cardiovascular system|CARDIOVASCULAR
Disorder|Disease or Syndrome|Past Medical History|1911,1933|false|false|false|C0007222|Cardiovascular Diseases|CARDIOVASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|1926,1933|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|1926,1933|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|1937,1964|false|false|false|C0085096|Peripheral Vascular Diseases|PERIPHERAL VASCULAR DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1948,1956|false|false|false|C0005847|Blood Vessel|VASCULAR
Disorder|Disease or Syndrome|Past Medical History|1948,1964|false|false|false|C0042373|Vascular Diseases|VASCULAR DISEASE
Disorder|Disease or Syndrome|Past Medical History|1957,1964|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|1957,1964|false|false|false|||DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1968,1975|false|false|false|C0042027|Urinary tract|URINARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1968,1981|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|URINARY TRACT
Anatomy|Body System|Past Medical History|1968,1981|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|URINARY TRACT
Disorder|Disease or Syndrome|Past Medical History|1968,1991|false|false|false|C0042029|Urinary tract infection|URINARY TRACT INFECTION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1976,1981|false|false|false|C1185740|Tract|TRACT
Disorder|Disease or Syndrome|Past Medical History|1982,1991|false|false|false|C0009450|Communicable Diseases|INFECTION
Event|Event|Past Medical History|1982,1991|false|false|false|||INFECTION
Finding|Pathologic Function|Past Medical History|1982,1991|false|false|false|C3714514|Infection|INFECTION
Disorder|Disease or Syndrome|Past Medical History|1995,2003|false|false|false|C0086543|Cataract|CATARACT
Event|Event|Past Medical History|1995,2003|false|false|false|||CATARACT
Finding|Finding|Past Medical History|1995,2003|false|false|false|C1690964|cataract on exam (physical finding)|CATARACT
Finding|Finding|Past Medical History|1995,2011|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Finding|Intellectual Product|Past Medical History|1995,2011|false|false|false|C1548833;C2186377|Consent Type - Cataract Surgery;reported history of cataract surgery|CATARACT SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1995,2011|false|false|false|C0007389;C2939459|Cataract Extraction;Cataract surgery|CATARACT SURGERY
Event|Event|Past Medical History|2004,2011|false|false|false|||SURGERY
Finding|Finding|Past Medical History|2004,2011|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Past Medical History|2004,2011|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Past Medical History|2004,2011|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2004,2011|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Finding|Past Medical History|2018,2025|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Past Medical History|2018,2025|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Past Medical History|2018,2025|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2018,2025|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Finding|Functional Concept|Past Medical History|2037,2043|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Finding|Intellectual Product|Past Medical History|2037,2043|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|COMMON
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2037,2056|false|false|false|C1261084|Common iliac artery structure|COMMON ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2044,2049|false|false|false|C0020889|Bone structure of ilium|ILIAC
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2044,2056|false|false|false|C0020887|Structure of iliac artery|ILIAC ARTERY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2050,2056|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|2050,2056|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Event|Event|Past Medical History|2057,2065|false|false|false|||STENTING
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2057,2065|false|false|false|C2348535|Stenting|STENTING
Event|Event|Past Medical History|2071,2083|false|false|false|||BUNIONECTOMY
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2071,2083|false|false|false|C1542057|Silver bunionectomy|BUNIONECTOMY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2087,2090|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|HIP
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2087,2090|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Biologically Active Substance|Past Medical History|2087,2090|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Drug|Pharmacologic Substance|Past Medical History|2087,2090|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|HIP
Event|Event|Past Medical History|2087,2090|false|false|false|||HIP
Finding|Gene or Genome|Past Medical History|2087,2090|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2087,2090|false|false|false|C1292890|Procedure on hip|HIP
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2087,2102|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|HIP REPLACEMENT
Event|Event|Past Medical History|2091,2102|false|false|false|||REPLACEMENT
Finding|Functional Concept|Past Medical History|2091,2102|false|false|false|C0559956|Replacement|REPLACEMENT
Procedure|Health Care Activity|Past Medical History|2091,2102|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2091,2102|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|REPLACEMENT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2112,2120|false|false|false|C3841297|Cesarean|CESAREAN
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2112,2128|false|false|false|C0007876|Cesarean section|CESAREAN SECTION
Drug|Substance|Past Medical History|2121,2128|false|false|false|C1522472|section sample|SECTION
Event|Event|Past Medical History|2121,2128|false|false|false|||SECTION
Finding|Intellectual Product|Past Medical History|2121,2128|false|false|false|C1551341;C1552858|Act Class - Section;Html Link Type - section|SECTION
Procedure|Laboratory Procedure|Past Medical History|2121,2128|false|false|false|C0700320|Sectioning technique|SECTION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2132,2140|false|false|false|C0017067|Ganglia|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2132,2140|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION
Disorder|Anatomical Abnormality|Past Medical History|2132,2145|false|false|false|C0085648;C1258666|Myxoid cyst;Synovial Cyst|GANGLION CYST
Disorder|Anatomical Abnormality|Past Medical History|2141,2145|false|false|false|C0010709|Cyst|CYST
Event|Event|Past Medical History|2141,2145|false|false|false|||CYST
Finding|Body Substance|Past Medical History|2141,2145|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Intellectual Product|Past Medical History|2141,2145|false|false|false|C1546594;C1550626|SpecimenType - Cyst|CYST
Finding|Idea or Concept|Family Medical History|2185,2191|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2198,2201|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|2198,2201|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|2204,2210|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2204,2210|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|2221,2228|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2221,2228|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2221,2228|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2236,2243|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|2236,2243|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2236,2243|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|2253,2261|false|false|false|||Physical
Finding|Finding|Family Medical History|2253,2261|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|2253,2261|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|2253,2261|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|2267,2276|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|Family Medical History|2277,2285|false|false|false|||PHYSICAL
Finding|Finding|Family Medical History|2277,2285|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|2277,2285|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|2277,2285|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|2277,2290|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|2277,2290|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|Family Medical History|2286,2290|false|false|false|||EXAM
Finding|Functional Concept|Family Medical History|2286,2290|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|2286,2290|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|Family Medical History|2339,2342|false|false|false|||P71
Finding|Gene or Genome|Family Medical History|2339,2342|false|false|false|C1425481|ZNF398 gene|P71
Event|Event|Family Medical History|2357,2364|false|false|false|||GENERAL
Finding|Classification|Family Medical History|2357,2364|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|2357,2364|false|false|false|C3812897|General medical service|GENERAL
Event|Event|Family Medical History|2372,2380|false|false|false|||pleasant
Finding|Mental Process|Family Medical History|2372,2380|false|false|false|C2987187|Pleasant|pleasant
Event|Event|Family Medical History|2381,2387|false|false|false|||affect
Finding|Mental Process|Family Medical History|2381,2387|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Family Medical History|2381,2387|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|Family Medical History|2389,2392|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|2389,2392|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|2389,2392|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|2389,2392|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|2389,2392|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|2389,2392|false|false|false|||NAD
Finding|Finding|Family Medical History|2389,2392|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|2393,2398|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2400,2403|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|2400,2403|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|Family Medical History|2400,2403|false|false|false|||MMM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2408,2411|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|2408,2411|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|2408,2411|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|2408,2411|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|Family Medical History|2416,2419|true|false|false|||JVD
Finding|Finding|Family Medical History|2416,2419|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2420,2425|true|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|2420,2425|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|Family Medical History|2420,2425|true|false|false|||HEART
Finding|Sign or Symptom|Family Medical History|2420,2425|true|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|Family Medical History|2427,2430|true|false|false|||RRR
Event|Event|Family Medical History|2449,2456|true|false|false|||murmurs
Finding|Finding|Family Medical History|2449,2456|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|Family Medical History|2465,2469|true|false|false|||rubs
Finding|Finding|Family Medical History|2465,2469|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2471,2476|false|false|false|C0024109|Lung|LUNGS
Finding|Sign or Symptom|Family Medical History|2478,2498|false|false|false|C3666016|Coarse breath sounds|Coarse breath sounds
Finding|Body Substance|Family Medical History|2485,2491|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Family Medical History|2485,2498|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|Family Medical History|2492,2498|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|2492,2498|false|false|false|C0037709||sounds
Finding|Organism Function|Family Medical History|2508,2518|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Family Medical History|2508,2527|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Event|Event|Family Medical History|2519,2527|false|false|false|||wheezing
Finding|Sign or Symptom|Family Medical History|2519,2527|false|false|false|C0043144|Wheezing|wheezing
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2540,2543|true|false|false|C4281590|Structure of middle lobe of right lung|RML
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2544,2547|true|false|false|C1261075|Structure of right lower lobe of lung|RLL
Finding|Finding|Family Medical History|2544,2547|true|false|false|C5703311|Radiolucent Lines|RLL
Event|Event|Family Medical History|2548,2556|true|false|false|||crackles
Finding|Finding|Family Medical History|2548,2556|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|Family Medical History|2566,2569|true|false|false|||WOB
Disorder|Congenital Abnormality|Family Medical History|2574,2590|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2584,2590|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Family Medical History|2584,2590|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|Family Medical History|2592,2595|true|false|false|||use
Finding|Functional Concept|Family Medical History|2592,2595|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|2592,2595|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Attribute|Clinical Attribute|Family Medical History|2601,2605|true|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|Family Medical History|2601,2605|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|Family Medical History|2606,2614|true|false|false|||distress
Finding|Finding|Family Medical History|2606,2614|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|2606,2614|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|2615,2622|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|Family Medical History|2615,2622|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|Family Medical History|2615,2622|true|false|false|||ABDOMEN
Finding|Finding|Family Medical History|2615,2622|true|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|Family Medical History|2624,2628|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|2624,2628|false|false|false|||soft
Event|Event|Family Medical History|2630,2639|false|false|false|||nontender
Event|Event|Family Medical History|2641,2653|false|false|false|||nondistended
Disorder|Congenital Abnormality|Family Medical History|2672,2675|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|Family Medical History|2672,2675|false|false|false|||EXT
Finding|Gene or Genome|Family Medical History|2672,2675|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|Family Medical History|2677,2681|false|false|false|||Warm
Finding|Finding|Family Medical History|2677,2681|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|2677,2681|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|2688,2692|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|2693,2701|false|false|false|||perfused
Finding|Pathologic Function|Family Medical History|2706,2722|false|false|false|C0085649|Peripheral edema|peripheral edema
Attribute|Clinical Attribute|Family Medical History|2717,2722|false|false|false|C1717255||edema
Event|Event|Family Medical History|2717,2722|false|false|false|||edema
Finding|Pathologic Function|Family Medical History|2717,2722|false|false|false|C0013604|Edema|edema
Event|Event|Family Medical History|2730,2736|false|false|false|||calves
Anatomy|Body System|Family Medical History|2743,2747|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|Family Medical History|2743,2747|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|Family Medical History|2743,2747|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|Family Medical History|2743,2747|false|false|false|||SKIN
Finding|Body Substance|Family Medical History|2743,2747|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|Family Medical History|2743,2747|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|Family Medical History|2754,2758|true|false|false|||warm
Finding|Finding|Family Medical History|2754,2758|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|2754,2758|true|false|false|C0687712|warming process|warm
Event|Event|Family Medical History|2763,2769|true|false|false|||rashes
Finding|Sign or Symptom|Family Medical History|2763,2769|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2776,2781|true|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|Family Medical History|2796,2802|false|false|false|||speech
Finding|Organism Function|Family Medical History|2796,2802|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Family Medical History|2796,2802|false|false|false|C0846595|Speech assessment|speech
Disorder|Disease or Syndrome|Family Medical History|2804,2807|false|false|false|C0393702|Myoclonic Astatic Epilepsy|MAE
Event|Event|Family Medical History|2804,2807|false|false|false|||MAE
Finding|Gene or Genome|Family Medical History|2804,2807|false|false|false|C5960827|SLC6A1 wt Allele|MAE
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2804,2807|false|false|false|C0286540|MAV protocol|MAE
Finding|Body Substance|Family Medical History|2823,2832|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|2823,2832|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|2823,2832|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|2823,2832|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|Family Medical History|2833,2841|false|false|false|||PHYSICAL
Finding|Finding|Family Medical History|2833,2841|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|Family Medical History|2833,2841|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|Family Medical History|2833,2841|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|Family Medical History|2833,2846|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|Family Medical History|2833,2846|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|Family Medical History|2842,2846|false|false|false|||EXAM
Finding|Functional Concept|Family Medical History|2842,2846|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|Family Medical History|2842,2846|false|false|false|C0582103|Medical Examination|EXAM
Finding|Gene or Genome|Family Medical History|2903,2906|false|false|false|C1413957;C1418458|DDX17 gene;TWNK gene|P72
Finding|Intellectual Product|Family Medical History|2916,2919|false|false|false|C1548704|O29|O29
Event|Event|Family Medical History|2928,2935|false|false|false|||GENERAL
Finding|Classification|Family Medical History|2928,2935|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|2928,2935|false|false|false|C3812897|General medical service|GENERAL
Event|Event|Family Medical History|2943,2951|false|false|false|||pleasant
Finding|Mental Process|Family Medical History|2943,2951|false|false|false|C2987187|Pleasant|pleasant
Event|Event|Family Medical History|2952,2958|false|false|false|||affect
Finding|Mental Process|Family Medical History|2952,2958|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Family Medical History|2952,2958|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|Family Medical History|2960,2963|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|2960,2963|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|2960,2963|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|2960,2963|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|2960,2963|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|2960,2963|false|false|false|||NAD
Finding|Finding|Family Medical History|2960,2963|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|2964,2969|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2971,2974|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|2971,2974|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|Family Medical History|2971,2974|false|false|false|||MMM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2979,2982|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|2979,2982|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|2979,2982|true|false|false|||LAD
Finding|Gene or Genome|Family Medical History|2979,2982|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|Family Medical History|2987,2990|true|false|false|||JVD
Finding|Finding|Family Medical History|2987,2990|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2991,2996|true|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|2991,2996|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Event|Event|Family Medical History|2991,2996|true|false|false|||HEART
Finding|Sign or Symptom|Family Medical History|2991,2996|true|false|false|C0795691|HEART PROBLEM|HEART
Event|Event|Family Medical History|2998,3001|true|false|false|||RRR
Event|Event|Family Medical History|3020,3027|true|false|false|||murmurs
Finding|Finding|Family Medical History|3020,3027|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|Family Medical History|3036,3040|true|false|false|||rubs
Finding|Finding|Family Medical History|3036,3040|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3042,3047|false|false|false|C0024109|Lung|LUNGS
Finding|Sign or Symptom|Family Medical History|3049,3069|false|false|false|C3666016|Coarse breath sounds|Coarse breath sounds
Finding|Body Substance|Family Medical History|3056,3062|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Family Medical History|3056,3069|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|Family Medical History|3063,3069|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3063,3069|false|false|false|C0037709||sounds
Finding|Finding|Family Medical History|3079,3084|true|false|false|C3833383|Scant|scant
Finding|Organism Function|Family Medical History|3085,3095|true|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Family Medical History|3085,3102|true|false|false|C0231875|Expiratory wheezing|expiratory wheeze
Event|Event|Family Medical History|3096,3102|true|false|false|||wheeze
Finding|Sign or Symptom|Family Medical History|3096,3102|true|false|false|C0043144|Wheezing|wheeze
Event|Event|Family Medical History|3104,3106|true|false|false|||no
Event|Event|Family Medical History|3113,3116|true|false|false|||WOB
Disorder|Congenital Abnormality|Family Medical History|3121,3137|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|Family Medical History|3121,3141|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3131,3137|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Family Medical History|3131,3137|true|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|Family Medical History|3138,3141|true|false|false|||use
Finding|Functional Concept|Family Medical History|3138,3141|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|3138,3141|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Attribute|Clinical Attribute|Family Medical History|3147,3151|true|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|Family Medical History|3147,3151|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Event|Event|Family Medical History|3152,3160|true|false|false|||distress
Finding|Finding|Family Medical History|3152,3160|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|3152,3160|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|3161,3168|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|Family Medical History|3161,3168|true|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|Family Medical History|3161,3168|true|false|false|||ABDOMEN
Finding|Finding|Family Medical History|3161,3168|true|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|Family Medical History|3170,3174|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|3170,3174|false|false|false|||soft
Event|Event|Family Medical History|3176,3185|false|false|false|||nontender
Event|Event|Family Medical History|3187,3199|false|false|false|||nondistended
Disorder|Congenital Abnormality|Family Medical History|3218,3221|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|Family Medical History|3218,3221|false|false|false|||EXT
Finding|Gene or Genome|Family Medical History|3218,3221|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|Family Medical History|3223,3227|false|false|false|||Warm
Finding|Finding|Family Medical History|3223,3227|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3223,3227|false|false|false|C0687712|warming process|Warm
Finding|Finding|Family Medical History|3234,3238|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Family Medical History|3239,3247|false|false|false|||perfused
Finding|Pathologic Function|Family Medical History|3252,3268|false|false|false|C0085649|Peripheral edema|peripheral edema
Attribute|Clinical Attribute|Family Medical History|3263,3268|false|false|false|C1717255||edema
Event|Event|Family Medical History|3263,3268|false|false|false|||edema
Finding|Pathologic Function|Family Medical History|3263,3268|false|false|false|C0013604|Edema|edema
Event|Event|Family Medical History|3276,3282|false|false|false|||calves
Anatomy|Body System|Family Medical History|3289,3293|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|Family Medical History|3289,3293|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|Family Medical History|3289,3293|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|Family Medical History|3289,3293|false|false|false|||SKIN
Finding|Body Substance|Family Medical History|3289,3293|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|Family Medical History|3289,3293|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|Family Medical History|3300,3304|true|false|false|||warm
Finding|Finding|Family Medical History|3300,3304|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|Family Medical History|3300,3304|true|false|false|C0687712|warming process|warm
Event|Event|Family Medical History|3309,3315|true|false|false|||rashes
Finding|Sign or Symptom|Family Medical History|3309,3315|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Mental or Behavioral Dysfunction|Family Medical History|3322,3327|true|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|Family Medical History|3342,3348|false|false|false|||speech
Finding|Organism Function|Family Medical History|3342,3348|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Family Medical History|3342,3348|false|false|false|C0846595|Speech assessment|speech
Disorder|Disease or Syndrome|Family Medical History|3350,3353|false|false|false|C0393702|Myoclonic Astatic Epilepsy|MAE
Event|Event|Family Medical History|3350,3353|false|false|false|||MAE
Finding|Gene or Genome|Family Medical History|3350,3353|false|false|false|C5960827|SLC6A1 wt Allele|MAE
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3350,3353|false|false|false|C0286540|MAV protocol|MAE
Event|Event|Family Medical History|3400,3404|false|false|false|||LABS
Lab|Laboratory or Test Result|Family Medical History|3400,3404|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|3445,3450|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3445,3450|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3445,3450|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|3451,3454|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3459,3462|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3459,3462|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3459,3462|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3468,3471|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|3468,3471|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|3468,3471|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|3468,3471|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|3477,3480|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3477,3480|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|3486,3489|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|3486,3489|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|3486,3489|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3486,3489|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3486,3489|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3494,3497|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3494,3497|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|3494,3497|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|3494,3497|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3494,3497|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3494,3497|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|3503,3507|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|3503,3507|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|3522,3525|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3542,3547|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3542,3547|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3542,3547|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|3548,3551|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3557,3560|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3557,3560|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3557,3560|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3566,3569|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|3566,3569|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|3566,3569|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|3566,3569|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|3575,3578|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3575,3578|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|3585,3588|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|3585,3588|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|3585,3588|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3585,3588|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3585,3588|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3592,3595|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3592,3595|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|3592,3595|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|3592,3595|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3592,3595|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3592,3595|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|3601,3605|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|3601,3605|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|3620,3623|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3640,3645|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3640,3645|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3640,3645|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|Family Medical History|3661,3666|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|Family Medical History|3661,3666|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|Family Medical History|3661,3666|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|Family Medical History|3671,3674|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|Family Medical History|3671,3674|false|false|false|||Eos
Finding|Gene or Genome|Family Medical History|3671,3674|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|Family Medical History|3701,3706|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3701,3706|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3701,3706|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|3711,3714|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|3711,3714|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|3711,3714|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|Family Medical History|3736,3741|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3736,3741|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3736,3741|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|Family Medical History|3763,3764|false|false|false|||-
Drug|Inorganic Chemical|Family Medical History|3781,3785|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3781,3785|false|false|false|C0005367|Bicarbonates|HCO3
Event|Event|Family Medical History|3781,3785|false|false|false|||HCO3
Procedure|Laboratory Procedure|Family Medical History|3781,3785|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3810,3815|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3810,3815|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3810,3815|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3810,3823|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3810,3823|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3810,3823|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3816,3823|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3816,3823|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3816,3823|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|3816,3823|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|3816,3823|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3816,3823|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3869,3873|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3869,3873|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3869,3873|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3898,3903|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3898,3903|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3898,3903|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3904,3910|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|Family Medical History|3904,3910|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|Family Medical History|3927,3932|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3927,3932|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3927,3932|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3927,3940|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Family Medical History|3933,3940|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Family Medical History|3933,3940|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Family Medical History|3933,3940|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Family Medical History|3933,3940|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Family Medical History|3933,3940|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Family Medical History|3933,3940|false|false|false|||Calcium
Finding|Physiologic Function|Family Medical History|3933,3940|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Family Medical History|3933,3940|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|Family Medical History|3974,3979|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|3974,3979|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|3974,3979|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Family Medical History|3974,3987|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|Family Medical History|3980,3987|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|Family Medical History|3980,3987|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|Family Medical History|3980,3987|false|false|false|||Lactate
Procedure|Laboratory Procedure|Family Medical History|3980,3987|false|false|false|C0202115|Lactic acid measurement|Lactate
Event|Event|Family Medical History|4003,4008|false|false|false|||MICRO
Finding|Conceptual Entity|Family Medical History|4003,4008|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|Family Medical History|4003,4008|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|Family Medical History|4003,4008|false|false|false|C0085672|Microbiology procedure|MICRO
Event|Event|Family Medical History|4037,4047|false|false|false|||Urinalysis
Procedure|Laboratory Procedure|Family Medical History|4037,4047|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|Urinalysis
Finding|Body Substance|Family Medical History|4061,4066|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|Family Medical History|4061,4066|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|Family Medical History|4061,4066|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|Family Medical History|4061,4072|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|Family Medical History|4067,4072|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|Family Medical History|4067,4072|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|Family Medical History|4073,4076|false|false|false|||NEG
Finding|Finding|Family Medical History|4073,4076|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|Family Medical History|4077,4084|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|Family Medical History|4077,4084|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|Family Medical History|4077,4084|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|Family Medical History|4085,4088|false|false|false|||NEG
Finding|Finding|Family Medical History|4085,4088|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4089,4096|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|Family Medical History|4089,4096|false|false|false|C0033684|Proteins|Protein
Event|Event|Family Medical History|4089,4096|false|false|false|||Protein
Finding|Conceptual Entity|Family Medical History|4089,4096|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|Family Medical History|4089,4096|false|false|false|C0202202|Protein measurement|Protein
Event|Event|Family Medical History|4097,4099|false|false|false|||TR
Drug|Biologically Active Substance|Family Medical History|4101,4108|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|4101,4108|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|4101,4108|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|4101,4108|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|4101,4108|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|4101,4108|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|Family Medical History|4109,4112|false|false|false|||NEG
Finding|Finding|Family Medical History|4109,4112|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|Family Medical History|4113,4119|false|false|false|C0022634|Ketones|Ketone
Event|Event|Family Medical History|4120,4123|false|false|false|||NEG
Finding|Finding|Family Medical History|4120,4123|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|Family Medical History|4132,4135|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|Family Medical History|4144,4147|false|false|false|C5848551|Neg - answer|NEG
Event|Event|Family Medical History|4161,4164|false|false|false|||NEG
Finding|Finding|Family Medical History|4161,4164|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|Family Medical History|4177,4182|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|Family Medical History|4177,4182|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|Family Medical History|4177,4182|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|Family Medical History|4177,4186|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE RBC
Anatomy|Cell|Family Medical History|4183,4186|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|4183,4186|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|4183,4186|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|Family Medical History|4189,4192|true|false|false|C0023516|Leukocytes|WBC
Drug|Food|Family Medical History|4209,4214|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Immunologic Factor|Family Medical History|4209,4214|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Indicator, Reagent, or Diagnostic Aid|Family Medical History|4209,4214|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Drug|Pharmacologic Substance|Family Medical History|4209,4214|true|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|Yeast
Event|Event|Family Medical History|4209,4214|true|false|false|||Yeast
Event|Event|Family Medical History|4215,4219|true|false|false|||NONE
Disorder|Disease or Syndrome|Family Medical History|4221,4224|true|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4221,4224|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|Family Medical History|4221,4224|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|Family Medical History|4221,4224|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|Family Medical History|4221,4224|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|Family Medical History|4221,4224|true|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|Family Medical History|4221,4224|true|false|false|||Epi
Finding|Gene or Genome|Family Medical History|4221,4224|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|Family Medical History|4221,4224|true|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|Family Medical History|4221,4224|true|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Disorder|Disease or Syndrome|Family Medical History|4228,4233|true|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|Family Medical History|4228,4233|true|false|false|||Blood
Finding|Body Substance|Family Medical History|4228,4233|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|Family Medical History|4274,4281|false|false|false|||STUDIES
Procedure|Research Activity|Family Medical History|4274,4281|false|false|false|C0947630|Scientific Study|STUDIES
Event|Event|Family Medical History|4311,4314|false|false|false|||EKG
Finding|Intellectual Product|Family Medical History|4311,4314|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Family Medical History|4311,4314|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|Family Medical History|4316,4321|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|Family Medical History|4316,4321|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|Family Medical History|4316,4321|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|Family Medical History|4316,4321|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|Family Medical History|4316,4328|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|Family Medical History|4322,4328|false|false|false|||rhythm
Finding|Finding|Family Medical History|4322,4328|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|4322,4328|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4343,4349|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Family Medical History|4343,4365|false|false|false|C0033036|Atrial Premature Complexes|atrial premature beats
Finding|Finding|Family Medical History|4350,4359|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Finding|Pathologic Function|Family Medical History|4350,4359|false|false|false|C0151526;C4018905|Premature Birth;Too early|premature
Disorder|Disease or Syndrome|Family Medical History|4350,4365|false|false|false|C0340464|Premature Cardiac Complex|premature beats
Event|Event|Family Medical History|4360,4365|false|false|false|||beats
Finding|Functional Concept|Family Medical History|4367,4371|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Disease or Syndrome|Family Medical History|4373,4392|false|false|false|C0006384|Bundle-Branch Block|bundle-branch block
Drug|Chemical Viewed Structurally|Family Medical History|4380,4386|false|false|false|C1881507|Macromolecular Branch|branch
Drug|Biomedical or Dental Material|Family Medical History|4387,4392|false|false|false|C1706085|Block Dosage Form|block
Event|Event|Family Medical History|4387,4392|false|false|false|||block
Finding|Body Substance|Family Medical History|4387,4392|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|Family Medical History|4387,4392|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|Family Medical History|4387,4392|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|Family Medical History|4408,4436|false|false|false|C3279217|Repolarization abnormalities|repolarization abnormalities
Disorder|Congenital Abnormality|Family Medical History|4423,4436|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Family Medical History|4423,4436|false|false|false|||abnormalities
Finding|Functional Concept|Family Medical History|4423,4436|false|false|false|C0000769|teratologic|abnormalities
Event|Event|Family Medical History|4483,4489|false|false|false|||rhythm
Finding|Finding|Family Medical History|4483,4489|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Family Medical History|4483,4489|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Anatomy|Body Space or Junction|Family Medical History|4498,4503|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Family Medical History|4498,4503|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Family Medical History|4498,4503|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Family Medical History|4498,4503|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|Family Medical History|4506,4509|false|false|false|||CXR
Procedure|Diagnostic Procedure|Family Medical History|4506,4509|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Functional Concept|Family Medical History|4517,4522|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4517,4534|false|false|false|C4281590|Structure of middle lobe of right lung|Right middle lobe
Finding|Intellectual Product|Family Medical History|4523,4529|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4523,4534|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4530,4534|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Family Medical History|4530,4534|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Family Medical History|4535,4542|false|false|false|||opacity
Finding|Finding|Family Medical History|4535,4542|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Family Medical History|4535,4542|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Disorder|Disease or Syndrome|Family Medical History|4559,4568|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Family Medical History|4559,4568|false|false|false|||pneumonia
Event|Event|Hospital Course|4650,4653|false|false|false|||PMH
Finding|Finding|Hospital Course|4650,4653|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|Hospital Course|4657,4663|false|false|false|C0004096|Asthma|Asthma
Event|Event|Hospital Course|4657,4663|false|false|false|||Asthma
Disorder|Disease or Syndrome|Hospital Course|4665,4669|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4665,4669|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|4665,4669|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|4665,4669|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4671,4674|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4671,4674|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|4671,4674|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|4671,4674|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|4671,4674|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|4671,4674|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|4671,4674|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4671,4674|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Hazardous or Poisonous Substance|Hospital Course|4676,4683|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Immunologic Factor|Hospital Course|4676,4683|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Organic Chemical|Hospital Course|4676,4683|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Pharmacologic Substance|Hospital Course|4676,4683|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Attribute|Clinical Attribute|Hospital Course|4676,4687|false|false|false|C4522050||tobacco use
Finding|Finding|Hospital Course|4676,4687|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Finding|Individual Behavior|Hospital Course|4676,4687|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Event|Event|Hospital Course|4684,4687|false|false|false|||use
Finding|Functional Concept|Hospital Course|4684,4687|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|4684,4687|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Hospital Course|4693,4702|false|false|false|||presented
Event|Event|Hospital Course|4717,4726|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|4717,4736|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|4717,4736|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|4730,4736|false|false|false|C0225386|Breath|breath
Finding|Finding|Hospital Course|4741,4757|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|Hospital Course|4752,4757|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|4752,4757|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|4752,4757|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|4752,4757|false|false|false|C0010200|Coughing|cough
Finding|Body Substance|Hospital Course|4762,4768|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|4762,4768|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|Hospital Course|4780,4785|false|false|false|||found
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4794,4797|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Event|Event|Hospital Course|4798,4805|false|false|false|||opacity
Finding|Finding|Hospital Course|4798,4805|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Hospital Course|4798,4805|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|Hospital Course|4809,4812|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|4809,4812|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Classification|Hospital Course|4816,4826|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4816,4826|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|4842,4850|false|false|false|||referred
Event|Event|Hospital Course|4870,4876|false|false|false|||ISSUES
Disorder|Disease or Syndrome|Hospital Course|4907,4935|false|false|false|C0694549|Community-Acquired Pneumonia|Community Acquired Pneumonia
Disorder|Disease or Syndrome|Hospital Course|4926,4935|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|Hospital Course|4926,4935|false|false|false|||Pneumonia
Event|Event|Hospital Course|4939,4948|false|false|false|||presented
Finding|Classification|Hospital Course|4952,4962|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4952,4962|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body System|Hospital Course|4963,4973|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Activity|Hospital Course|4974,4985|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|4974,4985|false|false|false|||appointment
Event|Event|Hospital Course|5000,5009|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|5000,5019|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|5000,5019|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|5013,5019|false|false|false|C0225386|Breath|breath
Finding|Finding|Hospital Course|5024,5040|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|Hospital Course|5035,5040|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|5035,5040|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|5035,5040|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|5035,5040|false|false|false|C0010200|Coughing|cough
Finding|Body Substance|Hospital Course|5045,5051|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|5045,5051|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|Hospital Course|5063,5071|false|false|false|||referred
Finding|Intellectual Product|Hospital Course|5075,5087|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Hospital Course|5075,5087|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Hospital Course|5083,5087|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|5083,5087|false|false|false|||care
Finding|Finding|Hospital Course|5083,5087|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|5083,5087|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Hospital Course|5119,5122|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|5119,5122|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|5129,5135|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5136,5139|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Event|Event|Hospital Course|5140,5147|false|false|false|||opacity
Finding|Finding|Hospital Course|5140,5147|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Hospital Course|5140,5147|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Event|Event|Hospital Course|5151,5154|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|5151,5154|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|5168,5178|false|false|false|||underlying
Anatomy|Body Location or Region|Hospital Course|5179,5183|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5179,5183|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|5179,5183|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|5179,5183|false|false|false|C0740941|Lung Problem|lung
Event|Event|Hospital Course|5184,5193|false|false|false|||pathology
Finding|Functional Concept|Hospital Course|5184,5193|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|5184,5193|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|5184,5193|false|false|false|C0919386|Pathology procedure|pathology
Disorder|Disease or Syndrome|Hospital Course|5195,5199|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5195,5199|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5195,5199|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5195,5199|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Hazardous or Poisonous Substance|Hospital Course|5217,5224|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Immunologic Factor|Hospital Course|5217,5224|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Organic Chemical|Hospital Course|5217,5224|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Pharmacologic Substance|Hospital Course|5217,5224|true|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Attribute|Clinical Attribute|Hospital Course|5217,5228|false|false|false|C4522050||tobacco use
Finding|Finding|Hospital Course|5217,5228|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Finding|Individual Behavior|Hospital Course|5217,5228|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|tobacco use
Event|Event|Hospital Course|5225,5228|false|false|false|||use
Finding|Functional Concept|Hospital Course|5225,5228|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|5225,5228|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Hospital Course|5269,5277|false|false|false|||admitted
Finding|Functional Concept|Hospital Course|5290,5298|false|false|false|C1548602;C1704686|Initiate (source type);Initiation|initiate
Finding|Idea or Concept|Hospital Course|5290,5298|false|false|false|C1548602;C1704686|Initiate (source type);Initiation|initiate
Drug|Antibiotic|Hospital Course|5299,5310|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|5299,5310|false|false|false|||antibiotics
Drug|Organic Chemical|Hospital Course|5311,5319|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|5311,5319|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|5311,5319|false|false|false|||steroids
Event|Event|Hospital Course|5324,5330|false|false|false|||ensure
Event|Event|Hospital Course|5340,5348|false|false|false|||remained
Event|Event|Hospital Course|5361,5367|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|5361,5367|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5376,5379|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Event|Event|Hospital Course|5380,5393|false|false|false|||opacification
Event|Event|Hospital Course|5398,5408|false|false|false|||suggestive
Finding|Functional Concept|Hospital Course|5398,5408|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|5398,5411|false|false|false|C0332299|Suggestive of|suggestive of
Disorder|Congenital Abnormality|Hospital Course|5412,5415|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|5412,5415|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|5412,5415|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|5412,5415|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5412,5415|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Disorder|Disease or Syndrome|Hospital Course|5417,5421|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5417,5421|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5417,5421|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5417,5421|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5422,5427|false|false|false|||flare
Finding|Finding|Hospital Course|5422,5427|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Finding|Sign or Symptom|Hospital Course|5422,5427|false|false|false|C1517205;C3540542|Exacerbation of cGVHD;Flare|flare
Event|Event|Hospital Course|5438,5451|false|false|false|||consideration
Finding|Finding|Hospital Course|5438,5451|false|false|false|C0518609|Consideration|consideration
Finding|Finding|Hospital Course|5458,5466|false|false|false|C0277797|Apyrexial|afebrile
Attribute|Clinical Attribute|Hospital Course|5467,5473|false|false|false|C5889824||status
Event|Event|Hospital Course|5467,5473|false|false|false|||status
Finding|Idea or Concept|Hospital Course|5467,5473|false|false|false|C1546481|What subject filter - Status|status
Anatomy|Cell|Hospital Course|5485,5488|false|false|false|C0023516|Leukocytes|WBC
Event|Event|Hospital Course|5490,5494|false|false|false|||Exam
Finding|Functional Concept|Hospital Course|5490,5494|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|Hospital Course|5490,5494|false|false|false|C0582103|Medical Examination|Exam
Event|Event|Hospital Course|5496,5507|false|false|false|||significant
Finding|Idea or Concept|Hospital Course|5496,5507|false|false|false|C0750502|Significant|significant
Finding|Finding|Hospital Course|5512,5520|false|false|false|C0277797|Apyrexial|afebrile
Attribute|Clinical Attribute|Hospital Course|5521,5527|false|false|false|C5889824||status
Event|Event|Hospital Course|5521,5527|false|false|false|||status
Finding|Idea or Concept|Hospital Course|5521,5527|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Hospital Course|5529,5539|false|false|false|||saturation
Phenomenon|Natural Phenomenon or Process|Hospital Course|5529,5539|false|false|false|C0522534|Saturated|saturation
Drug|Biomedical or Dental Material|Hospital Course|5555,5563|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|5555,5563|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|5555,5563|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Sign or Symptom|Hospital Course|5577,5597|false|false|false|C3666016|Coarse breath sounds|coarse breath sounds
Finding|Body Substance|Hospital Course|5584,5590|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Hospital Course|5584,5597|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|Hospital Course|5591,5597|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|Hospital Course|5591,5597|false|false|false|C0037709||sounds
Finding|Organism Function|Hospital Course|5610,5620|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|Hospital Course|5610,5629|false|false|false|C0231875|Expiratory wheezing|expiratory wheezing
Event|Event|Hospital Course|5621,5629|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5621,5629|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|5639,5646|false|false|false|||treated
Drug|Organic Chemical|Hospital Course|5650,5658|false|false|false|C0721336|Levaquin|Levaquin
Drug|Pharmacologic Substance|Hospital Course|5650,5658|false|false|false|C0721336|Levaquin|Levaquin
Event|Event|Hospital Course|5672,5679|false|false|false|||planned
Drug|Organic Chemical|Hospital Course|5693,5701|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|5693,5701|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|5693,5701|false|false|false|||steroids
Event|Event|Hospital Course|5703,5711|false|false|false|||recieved
Drug|Organic Chemical|Hospital Course|5716,5732|false|false|false|C4519262|Methylprednisone|methylprednisone
Drug|Pharmacologic Substance|Hospital Course|5716,5732|false|false|false|C4519262|Methylprednisone|methylprednisone
Finding|Intellectual Product|Hospital Course|5733,5737|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|5741,5747|false|false|false|||course
Event|Event|Hospital Course|5751,5753|false|false|false|||PO
Drug|Hormone|Hospital Course|5755,5765|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|5755,5765|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|5755,5765|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|5755,5765|false|false|false|||prednisone
Event|Event|Hospital Course|5786,5796|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5786,5796|false|false|false|C0087111|Therapeutic procedure|treatments
Attribute|Clinical Attribute|Hospital Course|5801,5808|false|false|false|C3854129||symptom
Finding|Sign or Symptom|Hospital Course|5801,5808|false|false|false|C1457887|Symptoms|symptom
Drug|Organic Chemical|Hospital Course|5809,5815|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|Hospital Course|5809,5815|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|Hospital Course|5809,5815|false|false|false|||relief
Finding|Finding|Hospital Course|5809,5815|false|false|false|C0564405|Feeling relief|relief
Finding|Intellectual Product|Hospital Course|5829,5837|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|Hospital Course|5838,5847|false|false|false|||stability
Event|Event|Hospital Course|5857,5867|false|false|false|||discharged
Event|Event|Hospital Course|5868,5872|false|false|false|||home
Finding|Idea or Concept|Hospital Course|5868,5872|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5868,5872|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5868,5872|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|5882,5892|false|false|false|||outpatient
Finding|Classification|Hospital Course|5882,5892|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|5882,5892|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|5900,5903|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5900,5903|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|5900,5903|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5900,5903|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|5900,5903|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|5900,5903|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|5900,5903|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|5900,5903|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|5900,5903|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|5900,5903|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|5900,5903|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Intellectual Product|Hospital Course|5927,5931|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Hospital Course|5942,5946|false|false|false|||need
Event|Event|Hospital Course|5950,5958|false|false|false|||complete
Event|Event|Hospital Course|5959,5965|false|false|false|||course
Drug|Antibiotic|Hospital Course|5969,5980|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|Hospital Course|5969,5980|false|false|false|||Antibiotics
Drug|Organic Chemical|Hospital Course|5985,5993|false|false|false|C0038317|Steroids|Steroids
Drug|Pharmacologic Substance|Hospital Course|5985,5993|false|false|false|C0038317|Steroids|Steroids
Event|Event|Hospital Course|5985,5993|false|false|false|||Steroids
Event|Event|Hospital Course|6003,6013|false|false|false|||instructed
Event|Event|Hospital Course|6017,6025|false|false|false|||continue
Finding|Classification|Hospital Course|6030,6040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|6030,6040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|6041,6045|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6041,6045|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6041,6045|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6041,6045|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|6046,6055|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|6046,6055|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6046,6055|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6046,6055|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6046,6055|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6046,6063|false|false|false|C0040808|Treatment Protocols|treatment regimen
Event|Event|Hospital Course|6056,6063|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|6056,6063|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6056,6063|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|Hospital Course|6068,6077|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6068,6077|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6068,6077|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6080,6087|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|6080,6087|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|6080,6087|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6124,6132|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6124,6139|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Hospital Course|6124,6147|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6133,6139|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Hospital Course|6133,6139|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Hospital Course|6133,6147|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Hospital Course|6140,6147|false|false|false|C0012634|Disease|Disease
Event|Event|Hospital Course|6140,6147|false|false|false|||Disease
Event|Event|Hospital Course|6163,6170|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|6163,6170|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6163,6170|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|6163,6170|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6163,6173|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|6174,6177|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6174,6177|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|6174,6177|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|6174,6177|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|6174,6177|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|6174,6177|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|6174,6177|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6174,6177|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Location or Region|Hospital Course|6200,6205|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6200,6205|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6200,6210|true|true|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6200,6210|true|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6206,6210|true|false|false|C2598155||pain
Event|Event|Hospital Course|6206,6210|true|false|false|||pain
Finding|Functional Concept|Hospital Course|6206,6210|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6206,6210|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|6224,6239|true|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|6224,6239|true|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Hospital Course|6244,6247|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|6244,6247|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|6244,6247|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|Hospital Course|6252,6261|false|false|false|||unchanged
Finding|Finding|Hospital Course|6252,6261|false|false|false|C0442739||unchanged
Event|Event|Hospital Course|6296,6305|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|6309,6313|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6309,6313|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6309,6313|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|6314,6321|false|false|false|||dosages
Drug|Organic Chemical|Hospital Course|6325,6331|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|6325,6331|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|6325,6331|false|false|false|||plavix
Drug|Organic Chemical|Hospital Course|6334,6341|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|6334,6341|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|6334,6341|false|false|false|||aspirin
Event|Event|Hospital Course|6353,6364|false|false|false|||mononitrate
Drug|Organic Chemical|Hospital Course|6369,6378|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6369,6378|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|6369,6378|false|false|false|||diltiazem
Disorder|Disease or Syndrome|Hospital Course|6381,6393|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|6381,6393|false|false|false|||Hypertension
Event|Event|Hospital Course|6409,6416|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|6409,6416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6409,6416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|6409,6416|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6409,6419|false|false|false|C0262926|Medical History|history of
Finding|Finding|Hospital Course|6409,6432|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|Hospital Course|6420,6432|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|6420,6432|false|false|false|||hypertension
Event|Event|Hospital Course|6441,6450|false|false|false|||continued
Event|Event|Hospital Course|6459,6463|false|false|false|||home
Finding|Idea or Concept|Hospital Course|6459,6463|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6459,6463|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6459,6463|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6469,6488|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|6469,6488|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Hospital Course|6469,6488|false|false|false|||hydrochlorothiazide
Disorder|Disease or Syndrome|Hospital Course|6492,6500|false|false|false|C0017601|Glaucoma|Glaucoma
Event|Event|Hospital Course|6492,6500|false|false|false|||Glaucoma
Event|Event|Hospital Course|6508,6517|false|false|false|||continued
Drug|Organic Chemical|Hospital Course|6521,6532|false|false|false|C0090306|latanoprost|latanoprost
Drug|Pharmacologic Substance|Hospital Course|6521,6532|false|false|false|C0090306|latanoprost|latanoprost
Drug|Biomedical or Dental Material|Hospital Course|6533,6538|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|Hospital Course|6533,6538|false|false|false|||drops
Disorder|Disease or Syndrome|Hospital Course|6546,6549|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|Hospital Course|6546,6549|false|false|false|||bed
Finding|Intellectual Product|Hospital Course|6546,6549|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|Hospital Course|6553,6567|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Hospital Course|6553,6567|false|false|false|||Hyperlipidemia
Finding|Finding|Hospital Course|6553,6567|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Event|Event|Hospital Course|6575,6584|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|6588,6592|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6588,6592|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6588,6592|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6598,6609|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|6598,6609|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Hospital Course|6598,6609|false|false|false|||simvastatin
Finding|Idea or Concept|Hospital Course|6612,6624|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Event|Event|Hospital Course|6666,6670|false|false|false|||need
Event|Event|Hospital Course|6674,6682|false|false|false|||continue
Drug|Organic Chemical|Hospital Course|6683,6691|false|false|false|C0721336|Levaquin|Levaquin
Drug|Pharmacologic Substance|Hospital Course|6683,6691|false|false|false|C0721336|Levaquin|Levaquin
Event|Event|Hospital Course|6692,6697|false|false|false|||750mg
Drug|Organic Chemical|Hospital Course|6707,6715|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|6707,6715|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|6707,6715|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|6707,6715|false|false|false|||complete
Finding|Functional Concept|Hospital Course|6707,6715|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6707,6715|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6719,6722|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6719,6722|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6723,6729|false|false|false|||course
Finding|Idea or Concept|Hospital Course|6731,6734|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Finding|Intellectual Product|Hospital Course|6731,6734|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Event|Event|Hospital Course|6754,6758|false|false|false|||need
Event|Event|Hospital Course|6762,6770|false|false|false|||continue
Drug|Hormone|Hospital Course|6771,6781|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|6771,6781|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|6771,6781|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|6796,6804|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|6796,6804|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|6796,6804|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|6796,6804|false|false|false|||complete
Finding|Functional Concept|Hospital Course|6796,6804|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6796,6804|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6808,6811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6808,6811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6812,6818|false|false|false|||course
Finding|Idea or Concept|Hospital Course|6820,6823|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Finding|Intellectual Product|Hospital Course|6820,6823|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|Day
Event|Event|Hospital Course|6843,6847|false|false|false|||need
Event|Event|Hospital Course|6851,6852|false|false|false|||f
Disorder|Disease or Syndrome|Hospital Course|6858,6861|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6858,6861|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|6858,6861|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6858,6861|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|6858,6861|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|6858,6861|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|6858,6861|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|6858,6861|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|6858,6861|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|6858,6861|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|6858,6861|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|6880,6888|false|false|false|||response
Finding|Finding|Hospital Course|6880,6888|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Hospital Course|6880,6888|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Hospital Course|6880,6888|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Classification|Hospital Course|6904,6911|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|Hospital Course|6904,6911|false|false|false|C3812897|General medical service|general
Attribute|Clinical Attribute|Hospital Course|6904,6918|false|false|false|C4018875||general health
Finding|Finding|Hospital Course|6904,6918|false|false|false|C0424575|General health|general health
Finding|Idea or Concept|Hospital Course|6912,6918|false|false|false|C0018684|Health|health
Procedure|Health Care Activity|Hospital Course|6912,6923|false|false|false|C0086388|Health Care|health care
Procedure|Health Care Activity|Hospital Course|6912,6935|false|false|false|C0262500|Health maintenance|health care maintenance
Event|Activity|Hospital Course|6919,6923|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|6919,6923|false|false|false|||care
Finding|Finding|Hospital Course|6919,6923|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|6919,6923|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Health Care Activity|Hospital Course|6919,6935|false|false|false|C0741961|CARE MAINTENANCE|care maintenance
Event|Activity|Hospital Course|6924,6935|false|false|false|C0024501|Maintenance|maintenance
Event|Event|Hospital Course|6924,6935|false|false|false|||maintenance
Event|Event|Hospital Course|6947,6951|false|false|false|||need
Event|Event|Hospital Course|6955,6958|false|false|false|||use
Event|Event|Hospital Course|6969,6979|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6969,6979|false|false|false|C0087111|Therapeutic procedure|treatments
Finding|Finding|Hospital Course|6980,6987|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Hospital Course|6983,6987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6983,6987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6983,6987|false|false|false|C1553498|home health encounter|home
Finding|Functional Concept|Hospital Course|6993,7004|false|false|false|C0231220|Symptomatic|symptomatic
Finding|Idea or Concept|Hospital Course|6993,7011|false|false|false|C3242309|symptomatic relief|symptomatic relief
Drug|Organic Chemical|Hospital Course|7005,7011|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|Hospital Course|7005,7011|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|Hospital Course|7005,7011|false|false|false|||relief
Finding|Finding|Hospital Course|7005,7011|false|false|false|C0564405|Feeling relief|relief
Finding|Idea or Concept|Hospital Course|7020,7024|false|false|false|C1552851|next - HtmlLinkType|next
Disorder|Disease or Syndrome|Hospital Course|7034,7043|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|7044,7050|false|false|false|||clears
Event|Occupational Activity|Hospital Course|7052,7056|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|7052,7056|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|Hospital Course|7052,7063|false|false|false|C0742531|CODE STATUS|Code Status
Attribute|Clinical Attribute|Hospital Course|7057,7063|false|false|false|C5889824||Status
Event|Event|Hospital Course|7057,7063|false|false|false|||Status
Finding|Idea or Concept|Hospital Course|7057,7063|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Hospital Course|7065,7069|false|false|false|||FULL
Event|Event|Hospital Course|7071,7080|false|false|false|||confirmed
Event|Activity|Hospital Course|7088,7095|false|false|false|C3812666|Personal Contact|Contact
Event|Event|Hospital Course|7088,7095|false|false|false|||Contact
Finding|Functional Concept|Hospital Course|7088,7095|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Idea or Concept|Hospital Course|7088,7095|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Finding|Intellectual Product|Hospital Course|7088,7095|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|Contact
Phenomenon|Phenomenon or Process|Hospital Course|7088,7095|false|false|false|C0392367|Physical contact|Contact
Attribute|Clinical Attribute|Hospital Course|7127,7138|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7127,7138|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|7127,7138|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|7127,7138|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|7127,7151|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|7142,7151|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|7142,7151|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|7170,7180|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|7170,7180|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|7170,7185|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|7181,7185|false|false|false|||list
Finding|Intellectual Product|Hospital Course|7181,7185|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|7189,7197|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|7202,7210|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|7202,7210|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|7202,7210|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|7202,7210|false|false|false|||complete
Finding|Functional Concept|Hospital Course|7202,7210|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7202,7210|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|7215,7224|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|7215,7224|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7232,7235|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|7232,7235|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|7232,7235|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|7232,7235|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|7232,7235|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7243,7246|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|7243,7246|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|7243,7246|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|7243,7246|false|false|false|||NEB
Finding|Cell Function|Hospital Course|7243,7246|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|7243,7246|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|7254,7257|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|7258,7267|false|false|false|||shortness
Finding|Body Substance|Hospital Course|7272,7278|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|7283,7292|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|7283,7292|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|7293,7300|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|7315,7318|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|7319,7328|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|7319,7338|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|7319,7338|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|7332,7338|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|7343,7352|false|false|false|C1121854|Symbicort|Symbicort
Drug|Pharmacologic Substance|Hospital Course|7343,7352|false|false|false|C1121854|Symbicort|Symbicort
Event|Event|Hospital Course|7343,7352|false|false|false|||Symbicort
Drug|Organic Chemical|Hospital Course|7354,7364|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|7354,7364|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|7354,7375|false|false|false|C1276807|budesonide / formoterol|budesonide-formoterol
Drug|Organic Chemical|Hospital Course|7365,7375|false|false|false|C0060657|formoterol|formoterol
Drug|Pharmacologic Substance|Hospital Course|7365,7375|false|false|false|C0060657|formoterol|formoterol
Event|Event|Hospital Course|7365,7375|false|false|false|||formoterol
Finding|Functional Concept|Hospital Course|7400,7410|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|7400,7410|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7411,7414|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7411,7414|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7411,7414|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7411,7414|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7411,7414|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7419,7430|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|7419,7430|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|7450,7459|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|7450,7459|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|7460,7468|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7460,7468|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|7469,7476|false|false|false|||Release
Finding|Functional Concept|Hospital Course|7469,7476|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7469,7476|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7469,7476|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|7497,7508|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|7497,7508|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|7497,7508|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|7497,7519|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|7497,7519|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|7509,7519|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7520,7525|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|7520,7525|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|7520,7525|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|7520,7525|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|7520,7525|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|7520,7525|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|7528,7532|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|7542,7545|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7546,7551|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|7546,7551|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|7546,7551|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|7546,7551|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Event|Event|Hospital Course|7546,7551|false|false|false|||nasal
Finding|Finding|Hospital Course|7546,7551|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|7546,7551|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Event|Event|Hospital Course|7553,7563|false|false|false|||congestion
Finding|Pathologic Function|Hospital Course|7553,7563|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Hospital Course|7568,7587|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|7568,7587|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|7607,7617|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|7607,7617|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|7607,7629|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|7607,7629|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|7618,7629|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|7631,7639|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7631,7639|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|7640,7647|false|false|false|||Release
Finding|Functional Concept|Hospital Course|7640,7647|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7640,7647|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7640,7647|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|7669,7680|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|7669,7680|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|7688,7693|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|7703,7707|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|7703,7707|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|7708,7712|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|7708,7712|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7708,7716|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|7708,7716|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|7713,7716|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7713,7716|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|7713,7716|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|7713,7716|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|7713,7716|false|false|false|||EYE
Finding|Body Substance|Hospital Course|7713,7716|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|7713,7716|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|7713,7716|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|7725,7736|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|7725,7736|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|Hospital Course|7757,7769|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|7757,7769|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|7757,7769|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|7757,7769|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|7757,7772|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Hospital Course|7757,7772|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|Hospital Course|7770,7772|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7783,7786|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7783,7786|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7783,7786|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|7783,7786|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|7783,7786|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|7792,7802|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|7792,7802|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|7792,7802|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|7792,7810|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|7792,7810|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|7803,7810|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|7803,7810|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|7803,7810|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|7813,7816|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|7813,7816|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|7813,7816|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|7813,7816|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7813,7816|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|7831,7844|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7831,7844|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|7831,7844|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7831,7844|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|7859,7862|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|7863,7867|false|false|false|C2598155||pain
Event|Event|Hospital Course|7863,7867|false|false|false|||pain
Finding|Functional Concept|Hospital Course|7863,7867|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7863,7867|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|7873,7880|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|7873,7880|false|false|false|C0004057|aspirin|Aspirin
Drug|Inorganic Chemical|Hospital Course|7901,7908|false|false|false|C0719084|CalCarb|Calcarb
Event|Event|Hospital Course|7901,7908|false|false|false|||Calcarb
Drug|Organic Chemical|Hospital Course|7918,7925|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|7918,7925|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|7918,7925|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|7918,7927|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|7918,7927|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|7918,7927|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|7918,7927|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|7918,7927|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|Hospital Course|7929,7936|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|7929,7936|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|7929,7936|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|7929,7936|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|7929,7936|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|7929,7936|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|7929,7936|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|7929,7936|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|7929,7946|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|7929,7946|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|7937,7946|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|7937,7946|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|7937,7946|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Hospital Course|7937,7946|false|false|false|||carbonate
Drug|Organic Chemical|Hospital Course|7947,7954|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|7947,7954|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|7947,7954|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|7947,7954|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|7947,7957|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|7947,7957|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|7947,7957|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|7971,7975|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|7971,7975|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|7971,7975|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|7971,7975|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7987,7990|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|7987,7990|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|7987,7990|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|7987,7990|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|Hospital Course|7987,7990|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|7987,7990|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|7987,7990|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|7987,8000|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|7987,8000|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|7987,8000|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7991,7996|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|7991,7996|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|7991,7996|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|7991,7996|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|7991,7996|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|7991,7996|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|7991,7996|false|false|false|||liver
Finding|Finding|Hospital Course|7991,7996|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|7991,7996|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|7997,8000|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|7997,8000|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|7997,8000|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|7997,8000|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Space or Junction|Hospital Course|8016,8020|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8016,8020|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8016,8020|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8016,8020|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8021,8024|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8021,8024|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8021,8024|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8021,8024|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8021,8024|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8030,8043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|8030,8043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|8030,8043|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|8030,8043|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|8046,8054|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|8046,8054|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|8057,8060|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|8057,8060|false|false|false|||TAB
Event|Event|Hospital Course|8074,8083|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|8074,8083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8074,8083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8074,8083|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8074,8083|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8074,8095|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8084,8095|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8084,8095|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8084,8095|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8084,8095|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8100,8113|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8100,8113|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|8100,8113|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8100,8113|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8128,8131|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8132,8136|false|false|false|C2598155||pain
Event|Event|Hospital Course|8132,8136|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8132,8136|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8132,8136|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|8141,8150|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8141,8150|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8158,8161|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8158,8161|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8158,8161|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|8158,8161|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8158,8161|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8169,8172|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|8169,8172|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|8169,8172|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|8169,8172|false|false|false|||NEB
Finding|Cell Function|Hospital Course|8169,8172|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8169,8172|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|8180,8183|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8184,8193|false|false|false|||shortness
Finding|Body Substance|Hospital Course|8198,8204|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|8209,8216|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8209,8216|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8236,8247|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|8236,8247|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|8267,8276|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8267,8276|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8277,8285|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8286,8293|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8286,8293|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8286,8293|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8314,8325|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8314,8325|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|8314,8325|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|8314,8336|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|8314,8336|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|8326,8336|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8337,8342|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|8337,8342|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|8337,8342|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|8337,8342|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|8337,8342|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|8337,8342|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|8345,8349|false|false|false|||SPRY
Finding|Gene or Genome|Hospital Course|8359,8362|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8363,8368|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8363,8368|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8363,8368|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8363,8368|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Event|Event|Hospital Course|8363,8368|false|false|false|||nasal
Finding|Finding|Hospital Course|8363,8368|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8363,8368|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Event|Event|Hospital Course|8370,8380|false|false|false|||congestion
Finding|Pathologic Function|Hospital Course|8370,8380|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Hospital Course|8385,8404|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|8385,8404|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|8424,8434|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|8424,8434|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|8424,8446|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|8424,8446|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|8435,8446|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|8448,8456|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8448,8456|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8457,8464|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8457,8464|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8457,8464|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8457,8464|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8486,8497|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|8486,8497|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|8505,8510|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8520,8524|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8520,8524|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|8525,8529|false|false|false|||LEFT
Finding|Functional Concept|Hospital Course|8525,8529|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8525,8533|false|false|false|C0229090|Left eye structure|LEFT EYE
Procedure|Diagnostic Procedure|Hospital Course|8525,8533|false|false|false|C2141124|examination of left eye|LEFT EYE
Anatomy|Body Location or Region|Hospital Course|8530,8533|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8530,8533|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|EYE
Disorder|Disease or Syndrome|Hospital Course|8530,8533|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Disorder|Neoplastic Process|Hospital Course|8530,8533|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|EYE
Event|Event|Hospital Course|8530,8533|false|false|false|||EYE
Finding|Body Substance|Hospital Course|8530,8533|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Finding|Hospital Course|8530,8533|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Finding|Intellectual Product|Hospital Course|8530,8533|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|EYE
Drug|Organic Chemical|Hospital Course|8542,8555|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|8542,8555|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|8542,8555|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|8542,8555|false|false|false|||Multivitamins
Drug|Inorganic Chemical|Hospital Course|8558,8566|false|false|false|C0026162|Minerals|minerals
Event|Event|Hospital Course|8558,8566|false|false|false|||minerals
Drug|Biomedical or Dental Material|Hospital Course|8569,8572|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|8569,8572|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|8587,8598|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Pharmacologic Substance|Hospital Course|8587,8598|false|false|false|C0074554|simvastatin|Simvastatin
Drug|Organic Chemical|Hospital Course|8619,8631|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|8619,8631|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|8619,8631|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|8619,8631|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|8619,8634|false|false|false|C2241157|Theophylline ER|Theophylline ER
Drug|Pharmacologic Substance|Hospital Course|8619,8634|false|false|false|C2241157|Theophylline ER|Theophylline ER
Event|Event|Hospital Course|8632,8634|false|false|false|||ER
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8645,8648|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8645,8648|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8645,8648|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8645,8648|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8645,8648|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8654,8664|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|8654,8664|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|8654,8664|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|8654,8672|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|8654,8672|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|8665,8672|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|8665,8672|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|8665,8672|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|8675,8678|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|8675,8678|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|8675,8678|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|8675,8678|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8675,8678|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|8693,8702|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8693,8702|false|false|false|C0001927|albuterol|Albuterol
Finding|Functional Concept|Hospital Course|8703,8710|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Gene or Genome|Hospital Course|8725,8728|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|8729,8738|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|8729,8748|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|8729,8748|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|8742,8748|false|false|false|C0225386|Breath|breath
Drug|Inorganic Chemical|Hospital Course|8754,8761|false|false|false|C0719084|CalCarb|Calcarb
Event|Event|Hospital Course|8754,8761|false|false|false|||Calcarb
Drug|Organic Chemical|Hospital Course|8771,8778|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|8771,8778|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|8771,8778|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|8771,8780|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|8771,8780|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|8771,8780|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|8771,8780|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|8771,8780|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Biologically Active Substance|Hospital Course|8782,8789|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|8782,8789|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|8782,8789|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|8782,8789|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|8782,8789|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|8782,8789|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|8782,8789|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|8782,8789|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|8782,8799|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|8782,8799|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|8790,8799|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|8790,8799|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|8790,8799|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Hospital Course|8790,8799|false|false|false|||carbonate
Drug|Organic Chemical|Hospital Course|8800,8807|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|8800,8807|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|8800,8807|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|8800,8807|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|8800,8810|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|8800,8810|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|8800,8810|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|8824,8828|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8824,8828|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8824,8828|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8824,8828|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8840,8843|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|8840,8843|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|8840,8843|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|8840,8843|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Finding|Finding|Hospital Course|8840,8843|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|8840,8843|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|8840,8843|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|8840,8853|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|8840,8853|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|8840,8853|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8844,8849|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|8844,8849|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|8844,8849|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|8844,8849|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|8844,8849|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|8844,8849|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|8844,8849|false|false|false|||liver
Finding|Finding|Hospital Course|8844,8849|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|8844,8849|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|8850,8853|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|8850,8853|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|8850,8853|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|8850,8853|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Space or Junction|Hospital Course|8869,8873|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8869,8873|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8869,8873|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8869,8873|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8874,8877|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8874,8877|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8874,8877|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8874,8877|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8874,8877|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8883,8892|false|false|false|C1121854|Symbicort|Symbicort
Drug|Pharmacologic Substance|Hospital Course|8883,8892|false|false|false|C1121854|Symbicort|Symbicort
Event|Event|Hospital Course|8883,8892|false|false|false|||Symbicort
Drug|Organic Chemical|Hospital Course|8894,8904|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|8894,8904|false|false|false|C0054201|budesonide|budesonide
Drug|Pharmacologic Substance|Hospital Course|8894,8915|false|false|false|C1276807|budesonide / formoterol|budesonide-formoterol
Drug|Organic Chemical|Hospital Course|8905,8915|false|false|false|C0060657|formoterol|formoterol
Drug|Pharmacologic Substance|Hospital Course|8905,8915|false|false|false|C0060657|formoterol|formoterol
Event|Event|Hospital Course|8905,8915|false|false|false|||formoterol
Event|Event|Hospital Course|8940,8950|false|false|false|||INHALATION
Finding|Functional Concept|Hospital Course|8940,8950|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|INHALATION
Finding|Organism Function|Hospital Course|8940,8950|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|INHALATION
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8951,8954|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8951,8954|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8951,8954|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8951,8954|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8951,8954|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8960,8968|false|false|false|C0719218|Cepastat|Cepastat
Drug|Pharmacologic Substance|Hospital Course|8960,8968|false|false|false|C0719218|Cepastat|Cepastat
Drug|Organic Chemical|Hospital Course|8970,8976|false|false|false|C0031428;C0070570|Phenols;phenol|Phenol
Drug|Pharmacologic Substance|Hospital Course|8970,8976|false|false|false|C0031428;C0070570|Phenols;phenol|Phenol
Drug|Biomedical or Dental Material|Hospital Course|8978,8985|false|false|false|C0991564|Oral Lozenge|Lozenge
Event|Event|Hospital Course|8988,8991|false|false|false|||LOZ
Finding|Gene or Genome|Hospital Course|8999,9002|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9003,9007|false|false|false|||sore
Finding|Sign or Symptom|Hospital Course|9003,9007|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|Hospital Course|9003,9014|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|Hospital Course|9003,9014|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|Hospital Course|9003,9014|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|Hospital Course|9003,9014|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|Hospital Course|9008,9014|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9008,9014|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Hospital Course|9008,9014|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Hospital Course|9008,9014|false|false|false|||throat
Finding|Body Substance|Hospital Course|9008,9014|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Hospital Course|9008,9014|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Hospital Course|9016,9018|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|9020,9026|false|false|false|C0031428;C0070570|Phenols;phenol|phenol
Drug|Pharmacologic Substance|Hospital Course|9020,9026|false|false|false|C0031428;C0070570|Phenols;phenol|phenol
Drug|Organic Chemical|Hospital Course|9028,9036|false|false|false|C0719218|Cepastat|Cepastat
Drug|Pharmacologic Substance|Hospital Course|9028,9036|false|false|false|C0719218|Cepastat|Cepastat
Event|Event|Hospital Course|9028,9036|false|false|false|||Cepastat
Drug|Biomedical or Dental Material|Hospital Course|9048,9056|false|false|false|C0991564|Oral Lozenge|lozenges
Event|Event|Hospital Course|9048,9056|false|false|false|||lozenges
Event|Event|Hospital Course|9070,9076|false|false|false|||needed
Event|Event|Hospital Course|9082,9086|false|false|false|||sore
Finding|Sign or Symptom|Hospital Course|9082,9086|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|Hospital Course|9082,9093|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|Hospital Course|9082,9093|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|Hospital Course|9082,9093|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|Hospital Course|9082,9093|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|Hospital Course|9087,9093|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9087,9093|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Hospital Course|9087,9093|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Hospital Course|9087,9093|false|false|false|||throat
Finding|Body Substance|Hospital Course|9087,9093|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Hospital Course|9087,9093|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Drug|Biomedical or Dental Material|Hospital Course|9104,9111|false|false|false|C0991564|Oral Lozenge|Lozenge
Event|Event|Hospital Course|9112,9119|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9112,9119|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|Hospital Course|9127,9139|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Organic Chemical|Hospital Course|9127,9139|false|false|false|C0282386|levofloxacin|Levofloxacin
Drug|Pharmacologic Substance|Hospital Course|9155,9163|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|9155,9163|false|false|false|||Duration
Event|Event|Hospital Course|9167,9171|false|false|false|||Days
Drug|Antibiotic|Hospital Course|9177,9189|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|9177,9189|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|9177,9189|false|false|false|||levofloxacin
Drug|Biomedical or Dental Material|Hospital Course|9199,9205|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9209,9217|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9212,9217|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9212,9217|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|9234,9240|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9241,9248|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9241,9248|false|false|false|C0807726|refill|Refills
Drug|Hormone|Hospital Course|9256,9266|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|9256,9266|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|9256,9266|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|9282,9290|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|9282,9290|false|false|false|||Duration
Event|Event|Hospital Course|9294,9298|false|false|false|||Days
Drug|Hormone|Hospital Course|9304,9314|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|9304,9314|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|9304,9314|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|9304,9314|false|false|false|||prednisone
Drug|Biomedical or Dental Material|Hospital Course|9323,9329|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9333,9341|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9336,9341|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9336,9341|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|9357,9363|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9357,9363|false|false|false|||Tablet
Event|Event|Hospital Course|9365,9372|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9365,9372|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|9379,9388|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9379,9388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9379,9388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9379,9388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9379,9388|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9379,9400|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9379,9400|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9389,9400|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|9389,9400|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|9389,9400|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|9402,9406|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|9402,9406|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9402,9406|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9402,9406|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|9409,9418|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9409,9418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9409,9418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9409,9418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9409,9418|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9409,9428|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9419,9428|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|9419,9428|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|9419,9428|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9419,9428|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9419,9428|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|9430,9458|false|false|false|C0694549|Community-Acquired Pneumonia|Community Acquired Pneumonia
Disorder|Disease or Syndrome|Hospital Course|9449,9458|false|false|false|C0032285|Pneumonia|Pneumonia
Event|Event|Hospital Course|9449,9458|false|false|false|||Pneumonia
Disorder|Disease or Syndrome|Hospital Course|9459,9463|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|9459,9463|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|9459,9463|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|9459,9463|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|9464,9470|false|false|false|C0004096|Asthma|Asthma
Event|Event|Hospital Course|9464,9470|false|false|false|||Asthma
Event|Event|Discharge Condition|9495,9504|false|false|false|||Discharge
Finding|Body Substance|Discharge Condition|9495,9504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Discharge Condition|9495,9504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Discharge Condition|9495,9504|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Discharge Condition|9495,9504|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Discharge Condition|9505,9514|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|Discharge Condition|9505,9514|false|false|false|C0012634|Disease|Condition
Event|Event|Discharge Condition|9505,9514|false|false|false|||Condition
Finding|Conceptual Entity|Discharge Condition|9505,9514|false|false|false|C1705253|Logical Condition|Condition
Event|Event|Discharge Condition|9516,9522|false|false|false|||Stable
Finding|Intellectual Product|Discharge Condition|9516,9522|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Mental Process|Discharge Condition|9523,9529|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9523,9536|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9523,9536|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9530,9536|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9530,9536|false|false|false|C1546481|What subject filter - Status|Status
Drug|Biomedical or Dental Material|Discharge Condition|9544,9552|false|false|false|C0168634|BaseLine dental cement|Baseline
Event|Event|Discharge Condition|9544,9552|false|false|false|||Baseline
Finding|Idea or Concept|Discharge Condition|9544,9552|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Event|Event|Discharge Condition|9554,9564|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|9554,9564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9554,9564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9554,9564|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9554,9564|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Classification|Discharge Condition|9554,9571|false|false|false|C1550332|Ambulatory Status|Ambulatory Status
Attribute|Clinical Attribute|Discharge Condition|9565,9571|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9565,9571|false|false|false|C1546481|What subject filter - Status|Status
Drug|Biomedical or Dental Material|Discharge Condition|9573,9581|false|false|false|C0168634|BaseLine dental cement|Baseline
Event|Event|Discharge Condition|9573,9581|false|false|false|||Baseline
Finding|Idea or Concept|Discharge Condition|9573,9581|false|false|false|C1552824|baseline - TableCellVerticalAlign|Baseline
Event|Event|Discharge Instructions|9628,9636|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|9628,9636|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9628,9636|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|9644,9648|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|9644,9648|false|false|false|||care
Finding|Finding|Discharge Instructions|9644,9648|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9644,9648|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9644,9651|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|9671,9683|false|false|false|||hospitalized
Event|Event|Discharge Instructions|9716,9724|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|9729,9736|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|Discharge Instructions|9737,9746|false|false|false|||treatment
Finding|Conceptual Entity|Discharge Instructions|9737,9746|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Discharge Instructions|9737,9746|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Discharge Instructions|9737,9746|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9737,9746|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|Discharge Instructions|9750,9759|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|9750,9759|false|false|false|||pneumonia
Event|Event|Discharge Instructions|9764,9770|false|false|false|||ensure
Event|Event|Discharge Instructions|9786,9796|false|false|false|||responding
Finding|Finding|Discharge Instructions|9797,9801|false|false|false|C5575035|Well (answer to question)|well
Drug|Antibiotic|Discharge Instructions|9809,9820|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|9809,9820|false|false|false|||antibiotics
Event|Event|Discharge Instructions|9833,9840|false|false|false|||history
Finding|Conceptual Entity|Discharge Instructions|9833,9840|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Discharge Instructions|9833,9840|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Discharge Instructions|9833,9840|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Discharge Instructions|9833,9843|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Discharge Instructions|9845,9849|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|9845,9849|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Discharge Instructions|9845,9849|false|false|false|||COPD
Finding|Gene or Genome|Discharge Instructions|9845,9849|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Discharge Instructions|9850,9856|false|false|false|C0004096|Asthma|Asthma
Event|Event|Discharge Instructions|9850,9856|false|false|false|||Asthma
Event|Event|Discharge Instructions|9875,9884|false|false|false|||responded
Event|Event|Discharge Instructions|9891,9895|false|false|false|||well
Finding|Finding|Discharge Instructions|9891,9895|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|9904,9916|false|false|false|||Antiobiotics
Drug|Organic Chemical|Discharge Instructions|9918,9926|false|false|false|C0038317|Steroids|Steroids
Drug|Pharmacologic Substance|Discharge Instructions|9918,9926|false|false|false|C0038317|Steroids|Steroids
Event|Event|Discharge Instructions|9918,9926|false|false|false|||Steroids
Event|Event|Discharge Instructions|9942,9952|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9942,9952|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|Discharge Instructions|9964,9976|false|false|false|||administered
Attribute|Clinical Attribute|Discharge Instructions|9989,9998|false|false|false|C5885990||breathing
Event|Event|Discharge Instructions|9989,9998|false|false|false|||breathing
Finding|Finding|Discharge Instructions|9989,9998|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|9989,9998|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|9989,9998|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|9989,9998|false|false|false|C1160636|respiratory system process|breathing
Event|Event|Discharge Instructions|10003,10009|false|false|false|||stable
Finding|Intellectual Product|Discharge Instructions|10003,10009|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|10024,10034|false|false|false|||responding
Event|Event|Discharge Instructions|10052,10062|false|false|false|||treatments
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10052,10062|false|false|false|C0087111|Therapeutic procedure|treatments
Event|Event|Discharge Instructions|10073,10083|false|false|false|||discharged
Event|Event|Discharge Instructions|10088,10092|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|10088,10092|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10088,10092|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10088,10092|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|10117,10125|false|false|false|||vigilant
Finding|Finding|Discharge Instructions|10117,10125|false|false|false|C0043012;C5240704|Vigilant (finding);Wakefulness|vigilant
Finding|Mental Process|Discharge Instructions|10117,10125|false|false|false|C0043012;C5240704|Vigilant (finding);Wakefulness|vigilant
Event|Event|Discharge Instructions|10136,10140|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10136,10140|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10151,10159|false|false|false|||continue
Drug|Antibiotic|Discharge Instructions|10164,10175|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|10164,10175|false|false|false|||antibiotics
Drug|Organic Chemical|Discharge Instructions|10178,10186|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Discharge Instructions|10178,10186|false|false|false|C0038317|Steroids|steroids
Event|Event|Discharge Instructions|10178,10186|false|false|false|||steroids
Event|Event|Discharge Instructions|10208,10214|false|false|false|||listed
Drug|Pharmacologic Substance|Discharge Instructions|10223,10233|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10223,10233|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10223,10233|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10234,10238|false|false|false|||page
Finding|Intellectual Product|Discharge Instructions|10234,10238|false|false|false|C1704732|Page (document)|page
Procedure|Laboratory Procedure|Discharge Instructions|10234,10238|false|false|false|C0013862|Polyacrylamide Gel Electrophoresis|page
Event|Event|Discharge Instructions|10259,10263|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|10259,10263|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|10267,10270|false|false|false|||see
Finding|Idea or Concept|Discharge Instructions|10288,10292|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Finding|Discharge Instructions|10288,10304|false|false|false|C1272171|Next appointment|next appointment
Event|Activity|Discharge Instructions|10293,10304|false|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|10293,10304|false|false|false|||appointment
Event|Event|Discharge Instructions|10308,10314|false|false|false|||ensure
Disorder|Disease or Syndrome|Discharge Instructions|10325,10334|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|10325,10334|false|false|false|||pneumonia
Event|Event|Discharge Instructions|10340,10348|false|false|false|||resolved
Procedure|Health Care Activity|Discharge Instructions|10352,10360|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10361,10373|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10361,10373|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10361,10373|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

