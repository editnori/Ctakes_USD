 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Organic Chemical|Allergies|183,193|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Allergies|183,193|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Allergies|183,193|false|false|false|||omeprazole
Drug|Biologically Active Substance|Allergies|196,202|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|196,202|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|196,202|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Event|Allergies|196,202|false|false|false|||Iodine
Drug|Inorganic Chemical|Allergies|207,213|false|false|false|C0021966|Iodides|Iodide
Event|Event|Allergies|207,213|false|false|false|||Iodide
Event|Activity|Allergies|214,224|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|214,224|false|false|false|C0332256|Containing (qualifier value)|Containing
Event|Event|Allergies|225,233|false|false|false|||Products
Drug|Hazardous or Poisonous Substance|Allergies|237,250|false|false|false|C0018533|Hallucinogens|hallucinogens
Drug|Pharmacologic Substance|Allergies|237,250|false|false|false|C0018533|Hallucinogens|hallucinogens
Event|Event|Allergies|237,250|false|false|false|||hallucinogens
Event|Event|Allergies|253,262|false|false|false|||Attending
Finding|Functional Concept|Allergies|253,262|false|false|false|C1999232|Attending (action)|Attending
Finding|Functional Concept|Chief Complaint|288,292|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|Chief Complaint|288,296|false|false|false|C0524471|Left hip region structure|Left hip
Finding|Sign or Symptom|Chief Complaint|288,301|false|false|false|C2141922|Pain of left hip joint|Left hip pain
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|293,296|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Chief Complaint|293,296|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Chief Complaint|293,296|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Chief Complaint|293,296|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Chief Complaint|293,296|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|293,296|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Chief Complaint|293,301|false|false|false|C1716793||hip pain
Finding|Sign or Symptom|Chief Complaint|293,301|false|false|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Chief Complaint|297,301|false|false|false|C2598155||pain
Event|Event|Chief Complaint|297,301|false|false|false|||pain
Finding|Functional Concept|Chief Complaint|297,301|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|297,301|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Classification|Chief Complaint|305,310|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|311,319|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|311,319|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|323,341|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|332,341|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|332,341|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|332,341|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|332,341|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|332,341|false|false|false|C0184661|Interventional procedure|Procedure
Attribute|Clinical Attribute|Chief Complaint|343,349|false|false|false|C5889824||Status
Event|Event|Chief Complaint|343,349|false|false|false|||Status
Finding|Idea or Concept|Chief Complaint|343,349|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Chief Complaint|355,359|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Chief Complaint|360,364|false|false|false|||CRPP
Event|Event|History of Present Illness|405,411|false|false|false|||REASON
Finding|Idea or Concept|History of Present Illness|405,411|false|false|false|C0392360|Indication of (contextual qualifier)|REASON
Finding|Idea or Concept|History of Present Illness|405,415|false|false|false|C0392360|Indication of (contextual qualifier)|REASON FOR
Event|Event|History of Present Illness|416,423|false|false|false|||CONSULT
Procedure|Health Care Activity|History of Present Illness|416,423|false|false|false|C0009818|Consultation|CONSULT
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|425,430|false|false|false|C0015811;C4299098|Femur;Lower extremity>Femur|Femur
Disorder|Injury or Poisoning|History of Present Illness|425,439|false|false|false|C0015802|Femoral Fractures|Femur fracture
Disorder|Injury or Poisoning|History of Present Illness|431,439|false|false|false|C0016658|Fracture|fracture
Event|Event|History of Present Illness|431,439|false|false|false|||fracture
Disorder|Disease or Syndrome|History of Present Illness|441,444|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|441,444|false|false|false|||HPI
Finding|Finding|History of Present Illness|441,444|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|441,444|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|457,465|false|false|false|||presents
Finding|Idea or Concept|History of Present Illness|475,480|false|false|false|C1552828|Table Frame - above|above
Disorder|Injury or Poisoning|History of Present Illness|481,489|false|false|false|C0016658|Fracture|fracture
Event|Event|History of Present Illness|481,489|false|false|false|||fracture
Event|Event|History of Present Illness|494,504|false|false|false|||mechanical
Finding|Functional Concept|History of Present Illness|494,504|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|494,504|false|false|false|C0699886|Mechanical Treatments|mechanical
Event|Event|History of Present Illness|505,509|false|false|false|||fall
Finding|Finding|History of Present Illness|505,509|false|false|false|C0085639|Falls|fall
Event|Event|History of Present Illness|532,539|false|false|false|||walking
Drug|Immunologic Factor|History of Present Illness|550,553|false|false|false|C1443014|Dog antigen|dog
Event|Event|History of Present Illness|550,553|false|false|false|||dog
Procedure|Laboratory Procedure|History of Present Illness|550,553|false|false|false|C2097312|allergy testing dog|dog
Event|Event|History of Present Illness|554,560|false|false|false|||pulled
Event|Event|History of Present Illness|564,569|false|false|false|||leash
Event|Event|History of Present Illness|574,578|false|false|false|||fell
Finding|Idea or Concept|History of Present Illness|589,598|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|History of Present Illness|589,598|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Attribute|Clinical Attribute|History of Present Illness|599,603|false|false|false|C2598155||pain
Event|Event|History of Present Illness|599,603|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|599,603|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|599,603|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|618,626|false|false|false|||movement
Finding|Organism Function|History of Present Illness|618,626|false|false|false|C0026649|Movement|movement
Event|Event|History of Present Illness|628,634|false|false|false|||Denies
Anatomy|Body Location or Region|History of Present Illness|635,639|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|635,639|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|History of Present Illness|635,639|true|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|635,639|true|false|false|C0876917|Procedure on head|Head
Event|Event|History of Present Illness|640,646|true|false|false|||strike
Event|Occupational Activity|History of Present Illness|640,646|true|false|false|C0038452|Strikes, Employee|strike
Event|Event|History of Present Illness|648,651|true|false|false|||LOC
Disorder|Disease or Syndrome|History of Present Illness|655,660|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|655,660|true|false|false|||blood
Finding|Body Substance|History of Present Illness|655,660|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Pharmacologic Substance|History of Present Illness|655,669|true|false|false|C0003280|Anticoagulants|blood thinners
Drug|Hazardous or Poisonous Substance|History of Present Illness|661,669|true|false|false|C0556614|Thinners|thinners
Event|Event|History of Present Illness|661,669|true|false|false|||thinners
Event|Event|History of Present Illness|671,677|false|false|false|||Denies
Event|Event|History of Present Illness|678,686|true|false|false|||numbness
Finding|Finding|History of Present Illness|678,686|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|678,686|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|History of Present Illness|690,698|true|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|690,698|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|706,717|true|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Disease or Syndrome|Past Medical History|746,750|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|746,750|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|756,776|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|Past Medical History|756,776|false|false|false|||Hypercholesterolemia
Finding|Finding|Past Medical History|756,776|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|782,788|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Past Medical History|782,788|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|Past Medical History|782,788|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Past Medical History|782,788|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Past Medical History|782,788|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Past Medical History|782,795|false|false|false|C0392525;C5779632|NEPHROLITHIASIS, CALCIUM OXALATE, 1;Nephrolithiasis|Kidney stones
Finding|Body Substance|Past Medical History|782,795|false|false|false|C0022650|Kidney Calculi|Kidney stones
Event|Event|Past Medical History|789,795|false|false|false|||stones
Finding|Body Substance|Past Medical History|789,795|false|false|false|C0006736|Calculi|stones
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|801,813|false|false|false|C0026264|Mitral Valve|Mitral valve
Disorder|Disease or Syndrome|Past Medical History|801,822|false|false|false|C0026267|Mitral Valve Prolapse Syndrome|Mitral valve prolapse
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|808,813|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|Past Medical History|814,822|false|false|false|C0033377|Ptosis|prolapse
Event|Event|Past Medical History|814,822|false|false|false|||prolapse
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|828,835|false|false|false|C0042149|Uterus|Uterine
Disorder|Neoplastic Process|Past Medical History|828,844|false|false|false|C0042133|Uterine Fibroids|Uterine fibroids
Disorder|Neoplastic Process|Past Medical History|836,844|false|false|false|C0023267;C0042133|Fibroid Tumor;Uterine Fibroids|fibroids
Event|Event|Past Medical History|836,844|false|false|false|||fibroids
Disorder|Disease or Syndrome|Past Medical History|850,862|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|Past Medical History|850,862|false|false|false|||Osteoporosis
Finding|Finding|Past Medical History|850,862|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|Past Medical History|868,876|false|false|false|C0149931|Migraine Disorders|Migraine
Disorder|Disease or Syndrome|Past Medical History|868,886|false|false|false|C0149931|Migraine Disorders|Migraine headaches
Event|Event|Past Medical History|877,886|false|false|false|||headaches
Finding|Sign or Symptom|Past Medical History|877,886|false|false|false|C0018681|Headache|headaches
Disorder|Disease or Syndrome|Family Medical History|928,931|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|928,931|false|false|false|||HTN
Event|Event|Family Medical History|934,940|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|934,940|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|934,940|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Disorder|Mental or Behavioral Dysfunction|Family Medical History|945,953|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Family Medical History|945,953|false|false|false|||Dementia
Event|Event|Family Medical History|956,962|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|956,962|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|956,962|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|General Exam|984,991|false|false|false|||General
Finding|Classification|General Exam|984,991|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|984,991|false|false|false|C3812897|General medical service|General
Finding|Finding|General Exam|993,997|true|false|false|C5575035|Well (answer to question)|Well
Event|Event|General Exam|998,1007|true|false|false|||appearing
Finding|Finding|General Exam|1015,1035|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|1021,1026|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|1027,1035|true|false|false|||distress
Finding|Finding|General Exam|1027,1035|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|1027,1035|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Functional Concept|General Exam|1038,1042|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|1038,1058|false|false|false|C0230416|Left lower extremity|Left Lower extremity
Anatomy|Body Location or Region|General Exam|1043,1048|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|General Exam|1043,1048|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|1043,1058|false|false|false|C0023216|Lower Extremity|Lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|1049,1058|false|false|false|C0015385|Limb structure|extremity
Anatomy|Body System|General Exam|1062,1066|true|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|1062,1066|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|1062,1066|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|1062,1066|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|1062,1066|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|1067,1073|true|false|false|||intact
Finding|Finding|General Exam|1067,1073|true|false|false|C1554187|Gender Status - Intact|intact
Disorder|Anatomical Abnormality|General Exam|1079,1088|true|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Disorder|Congenital Abnormality|General Exam|1079,1088|true|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Event|Event|General Exam|1079,1088|true|false|false|||deformity
Finding|Finding|General Exam|1079,1088|true|false|false|C2117111||deformity
Attribute|Clinical Attribute|General Exam|1090,1095|true|false|false|C1717255||edema
Event|Event|General Exam|1090,1095|true|false|false|||edema
Finding|Pathologic Function|General Exam|1090,1095|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|1097,1107|true|false|false|||ecchymosis
Finding|Finding|General Exam|1097,1107|true|false|false|C0013491;C3812660|Ecchymosis;Skin Bruise|ecchymosis
Finding|Pathologic Function|General Exam|1097,1107|true|false|false|C0013491;C3812660|Ecchymosis;Skin Bruise|ecchymosis
Disorder|Disease or Syndrome|General Exam|1109,1117|true|false|false|C0041834|Erythema|erythema
Event|Event|General Exam|1109,1117|true|false|false|||erythema
Event|Event|General Exam|1119,1129|false|false|false|||induration
Finding|Pathologic Function|General Exam|1119,1129|false|false|false|C0332534|Induration|induration
Disorder|Disease or Syndrome|General Exam|1132,1136|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|1132,1136|false|false|false|||Soft
Anatomy|Body Location or Region|General Exam|1149,1154|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Anatomy|Body Part, Organ, or Organ Component|General Exam|1159,1162|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Functional Concept|General Exam|1171,1179|false|false|false|C0234226|Painless|painless
Event|Event|General Exam|1180,1183|false|false|false|||ROM
Finding|Finding|General Exam|1180,1183|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|General Exam|1180,1183|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|General Exam|1180,1183|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Anatomy|Body Location or Region|General Exam|1184,1188|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|1184,1188|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|1184,1188|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|1184,1188|false|false|false|C0562271|Examination of knee joint|knee
Anatomy|Body Location or Region|General Exam|1194,1199|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Anatomy|Body Space or Junction|General Exam|1194,1199|false|false|false|C0003086;C0003087;C4284979|Ankle;Ankle joint structure;Lower extremity>Ankle|ankle
Disorder|Disease or Syndrome|General Exam|1202,1207|false|false|false|C4049262|Febrile infection related epilepsy syndrome|Fires
Event|Event|General Exam|1202,1207|false|false|false|||Fires
Event|Event|General Exam|1202,1207|false|false|false|C0016141|fire disaster|Fires
Phenomenon|Natural Phenomenon or Process|General Exam|1202,1207|false|false|false|C0700614|Fire (physical force)|Fires
Event|Event|General Exam|1219,1220|false|false|false|||S
Event|Event|General Exam|1223,1225|false|false|false|||SP
Drug|Food|General Exam|1254,1260|false|false|false|C5890763||pulses
Event|Event|General Exam|1254,1260|false|false|false|||pulses
Finding|Physiologic Function|General Exam|1254,1260|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|1254,1260|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|1262,1265|false|false|false|||WWP
Finding|Body Substance|Hospital Course|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1295,1302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1303,1312|false|false|false|||presented
Finding|Finding|Hospital Course|1320,1329|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Hospital Course|1320,1329|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Hospital Course|1320,1329|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Hospital Course|1320,1329|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Hospital Course|1320,1329|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Hospital Course|1320,1329|false|false|false|C1553500|emergency encounter|emergency
Event|Event|Hospital Course|1330,1340|false|false|false|||department
Finding|Idea or Concept|Hospital Course|1330,1340|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Event|Event|Hospital Course|1350,1359|false|false|false|||evaluated
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1367,1385|false|false|false|C0162439;C1136201|Orthopedic Rehabilitation Surgery;Orthopedic Surgical Procedures|orthopedic surgery
Event|Event|Hospital Course|1378,1385|false|false|false|||surgery
Finding|Finding|Hospital Course|1378,1385|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|1378,1385|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|1378,1385|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1378,1385|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Body Substance|Hospital Course|1396,1403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1396,1403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1396,1403|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1408,1413|false|false|false|||found
Finding|Functional Concept|Hospital Course|1425,1429|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Anatomical Abnormality|Hospital Course|1430,1436|false|false|false|C0042282|Valgus deformity|valgus
Event|Event|Hospital Course|1430,1436|false|false|false|||valgus
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1446,1453|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1446,1458|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|Hospital Course|1446,1467|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|Hospital Course|1454,1458|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|1454,1458|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|1454,1458|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Hospital Course|1454,1467|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|Hospital Course|1459,1467|false|false|false|C0016658|Fracture|fracture
Event|Event|Hospital Course|1459,1467|false|false|false|||fracture
Event|Event|Hospital Course|1477,1485|false|false|false|||admitted
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1493,1511|false|false|false|C0162439;C1136201|Orthopedic Rehabilitation Surgery;Orthopedic Surgical Procedures|orthopedic surgery
Event|Event|Hospital Course|1504,1511|false|false|false|||surgery
Finding|Finding|Hospital Course|1504,1511|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|1504,1511|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|1504,1511|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1504,1511|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Occupational Activity|Hospital Course|1512,1519|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|1512,1519|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Finding|Body Substance|Hospital Course|1525,1532|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1525,1532|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1525,1532|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1538,1543|false|false|false|||taken
Finding|Finding|Hospital Course|1551,1560|false|false|false|C4738506|Operating|operating
Finding|Functional Concept|Hospital Course|1577,1581|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|Hospital Course|1589,1598|false|false|false|||reduction
Finding|Finding|Hospital Course|1589,1598|false|false|false|C0392756|Reduced|reduction
Phenomenon|Natural Phenomenon or Process|Hospital Course|1589,1598|false|false|false|C0301630|Reduction (chemical)|reduction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1589,1598|false|false|false|C1293152;C4551656|Reduction procedure;Surgical reduction|reduction
Finding|Functional Concept|Hospital Course|1604,1616|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|Hospital Course|1617,1624|false|false|false|||pinning
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1617,1624|false|false|false|C0021885|Intramedullary Nailing|pinning
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1628,1631|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|1628,1631|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|1628,1631|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|1628,1631|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Event|Event|Hospital Course|1628,1631|false|false|false|||hip
Finding|Gene or Genome|Hospital Course|1628,1631|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1628,1631|false|false|false|C1292890|Procedure on hip|hip
Finding|Body Substance|Hospital Course|1643,1650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1643,1650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1643,1650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1651,1660|false|false|false|||tolerated
Event|Event|Hospital Course|1662,1666|false|false|false|||well
Finding|Finding|Hospital Course|1662,1666|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|1677,1684|false|false|false|||details
Attribute|Clinical Attribute|Hospital Course|1692,1701|false|false|false|C0945766||procedure
Event|Event|Hospital Course|1692,1701|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|1692,1701|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|1692,1701|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1692,1701|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Hospital Course|1709,1712|false|false|false|||see
Event|Event|Hospital Course|1729,1737|false|false|false|||dictated
Finding|Intellectual Product|Hospital Course|1738,1754|false|false|false|C1269801|Operative report|operative report
Attribute|Clinical Attribute|Hospital Course|1748,1754|false|false|false|C4255046||report
Event|Event|Hospital Course|1748,1754|false|false|false|||report
Finding|Intellectual Product|Hospital Course|1748,1754|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Hospital Course|1748,1754|false|false|false|C0700287|Reporting|report
Finding|Body Substance|Hospital Course|1760,1767|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1760,1767|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1760,1767|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|1772,1777|false|false|false|||taken
Event|Event|Hospital Course|1798,1802|false|false|false|||PACU
Finding|Intellectual Product|Hospital Course|1806,1812|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|1813,1822|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|1813,1822|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|1813,1822|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|1813,1822|false|false|false|C1705253|Logical Condition|condition
Event|Event|Hospital Course|1833,1845|false|false|false|||satisfactory
Finding|Intellectual Product|Hospital Course|1833,1845|false|false|false|C1547307|Satisfactory - Patient Condition Code|satisfactory
Event|Activity|Hospital Course|1847,1855|false|false|false|C0237820||recovery
Event|Event|Hospital Course|1847,1855|false|false|false|||recovery
Finding|Organism Function|Hospital Course|1847,1855|false|false|false|C2004454|Recovery - healing process|recovery
Attribute|Clinical Attribute|Hospital Course|1861,1871|false|false|false|C2926599||anesthesia
Drug|Pharmacologic Substance|Hospital Course|1861,1871|false|false|false|C4049933|Anesthesia substance|anesthesia
Event|Event|Hospital Course|1861,1871|false|false|false|||anesthesia
Finding|Finding|Hospital Course|1861,1871|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Finding|Sign or Symptom|Hospital Course|1861,1871|false|false|false|C0278134;C2219802|Absence of sensation|anesthesia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1861,1871|false|false|false|C0002903;C0002912|Anesthesia procedures;Dental anesthesia|anesthesia
Event|Event|Hospital Course|1876,1887|false|false|false|||transferred
Anatomy|Anatomical Structure|Hospital Course|1895,1900|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|Hospital Course|1907,1914|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|1907,1914|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|1907,1914|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Substance|Hospital Course|1938,1944|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|1938,1944|false|false|false|||fluids
Finding|Body Substance|Hospital Course|1938,1944|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1938,1944|false|false|false|C0016286|Fluid Therapy|fluids
Attribute|Clinical Attribute|Hospital Course|1952,1956|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|1952,1956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1952,1956|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Hospital Course|1957,1968|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|1957,1968|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|1957,1968|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|1957,1968|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|1975,1985|false|false|false|||progressed
Finding|Daily or Recreational Activity|Hospital Course|1991,2003|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|1999,2003|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1999,2003|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1999,2003|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1999,2003|false|false|false|C0012159|Diet therapy|diet
Anatomy|Body Space or Junction|Hospital Course|2008,2012|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2008,2012|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2008,2012|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2008,2012|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|Hospital Course|2013,2024|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|2013,2024|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|2013,2024|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|2013,2024|false|false|false|C4284232|Medications|medications
Finding|Body Substance|Hospital Course|2040,2047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2040,2047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2040,2047|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Antibiotic|Hospital Course|2062,2073|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|2062,2073|false|false|false|||antibiotics
Event|Event|Hospital Course|2079,2094|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|2079,2094|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|2079,2094|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2079,2094|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Hospital Course|2099,2106|false|false|false|||routine
Finding|Idea or Concept|Hospital Course|2099,2106|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|Hospital Course|2099,2106|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|Hospital Course|2099,2106|false|false|false|C1979801|Routine coag|routine
Finding|Body Substance|Hospital Course|2112,2119|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2112,2119|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2112,2119|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2122,2126|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|2122,2126|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|2122,2126|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|2127,2138|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|2127,2138|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|2127,2138|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|2127,2138|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|2145,2154|false|false|false|||continued
Event|Event|Hospital Course|2171,2186|false|false|false|||hospitalization
Procedure|Health Care Activity|Hospital Course|2171,2186|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Body Substance|Hospital Course|2192,2199|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2192,2199|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2192,2199|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2200,2206|false|false|false|||worked
Event|Event|Hospital Course|2221,2231|false|false|false|||determined
Event|Event|Hospital Course|2237,2246|false|false|false|||discharge
Finding|Body Substance|Hospital Course|2237,2246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|2237,2246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|2237,2246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|2237,2246|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2237,2254|false|false|false|C0184713|Discharge to home|discharge to home
Event|Event|Hospital Course|2250,2254|false|false|false|||home
Finding|Idea or Concept|Hospital Course|2250,2254|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|2250,2254|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|2250,2254|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|2250,2268|false|false|false|C4534324|Home with services|home with services
Event|Event|Hospital Course|2260,2268|false|false|false|||services
Event|Occupational Activity|Hospital Course|2260,2268|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|2260,2268|false|false|false|C1704289|Clinical Service|services
Event|Event|Hospital Course|2274,2285|false|false|false|||appropriate
Finding|Idea or Concept|Hospital Course|2295,2303|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|2295,2310|false|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|2295,2310|false|false|false|C0489547|Hospital course|hospital course
Event|Event|Hospital Course|2304,2310|false|false|false|||course
Event|Event|Hospital Course|2326,2338|false|false|false|||unremarkable
Finding|Finding|Hospital Course|2348,2352|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|2348,2352|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|2348,2352|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|2356,2365|false|false|false|||discharge
Finding|Body Substance|Hospital Course|2356,2365|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|2356,2365|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|2356,2365|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|2356,2365|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|2370,2377|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2370,2377|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2370,2377|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|2380,2384|false|false|false|C2598155||pain
Event|Event|Hospital Course|2380,2384|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2380,2384|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2380,2384|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|2389,2393|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|2394,2404|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|2411,2415|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2411,2415|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2411,2415|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2411,2415|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|Hospital Course|2416,2427|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|2416,2427|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|2416,2427|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|2416,2427|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|2429,2438|false|false|false|||incisions
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2429,2438|false|false|false|C0184898|Surgical incisions|incisions
Event|Activity|Hospital Course|2444,2449|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|Hospital Course|2444,2449|false|false|false|||clean
Event|Event|Hospital Course|2454,2460|false|false|false|||intact
Finding|Finding|Hospital Course|2454,2460|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Body Substance|Hospital Course|2471,2478|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2471,2478|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2471,2478|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2483,2490|false|false|false|||voiding
Finding|Functional Concept|Hospital Course|2483,2490|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Finding|Organism Function|Hospital Course|2483,2490|false|false|false|C0042034;C4067975|Urination;Voids|voiding
Finding|Organism Function|Hospital Course|2491,2497|false|false|false|C0560560|Moving|moving
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2498,2504|false|false|false|C0021853|Intestines|bowels
Finding|Body Substance|Hospital Course|2524,2531|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2524,2531|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2524,2531|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2537,2550|false|false|false|||weightbearing
Event|Event|Hospital Course|2554,2563|false|false|false|||tolerated
Finding|Functional Concept|Hospital Course|2571,2575|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2571,2591|false|false|false|C0230416|Left lower extremity|left lower extremity
Anatomy|Body Location or Region|Hospital Course|2576,2581|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|2576,2581|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2576,2591|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2582,2591|false|false|false|C0015385|Limb structure|extremity
Event|Event|Hospital Course|2606,2616|false|false|false|||discharged
Drug|Organic Chemical|Hospital Course|2620,2627|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Hospital Course|2620,2627|false|false|false|C0728963|Lovenox|Lovenox
Anatomy|Body Location or Region|Hospital Course|2632,2635|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|2632,2635|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|2632,2635|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2632,2647|false|false|false|C0853245|DVT prophylaxis|DVT prophylaxis
Event|Event|Hospital Course|2636,2647|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2636,2647|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Body Substance|Hospital Course|2653,2660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2653,2660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2653,2660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|2667,2673|false|false|false|||follow
Event|Event|Hospital Course|2690,2697|false|false|false|||routine
Finding|Idea or Concept|Hospital Course|2690,2697|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|Hospital Course|2690,2697|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|Hospital Course|2690,2697|false|false|false|C1979801|Routine coag|routine
Event|Event|Hospital Course|2710,2720|false|false|false|||discussion
Finding|Social Behavior|Hospital Course|2710,2720|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2710,2720|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Body Substance|Hospital Course|2739,2746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2739,2746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2739,2746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|2761,2770|false|false|false|C0945731||diagnosis
Event|Event|Hospital Course|2761,2770|false|false|false|||diagnosis
Finding|Classification|Hospital Course|2761,2770|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|2761,2770|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|2761,2770|false|false|false|C0011900|Diagnosis|diagnosis
Event|Event|Hospital Course|2775,2783|false|false|false|||expected
Event|Event|Hospital Course|2800,2806|false|false|false|||course
Event|Event|Hospital Course|2817,2824|false|false|false|||reasons
Finding|Idea or Concept|Hospital Course|2817,2824|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Event|Event|Hospital Course|2828,2832|false|false|false|||call
Event|Event|Hospital Course|2837,2843|false|false|false|||office
Finding|Idea or Concept|Hospital Course|2837,2843|false|false|false|C1549636|Address type - Office|office
Event|Event|Hospital Course|2848,2854|false|false|false|||return
Finding|Idea or Concept|Hospital Course|2862,2870|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|2880,2889|false|false|false|||questions
Event|Event|Hospital Course|2895,2903|false|false|false|||answered
Finding|Body Substance|Hospital Course|2910,2917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|2910,2917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|2910,2917|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|2941,2953|false|false|false|C3263700||instructions
Event|Event|Hospital Course|2941,2953|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|2941,2953|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Attribute|Clinical Attribute|Hospital Course|2980,2992|false|false|false|C3263700||instructions
Event|Event|Hospital Course|2980,2992|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|2980,2992|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Event|Event|Hospital Course|3013,3019|false|false|false|||follow
Finding|Functional Concept|Hospital Course|3013,3019|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|3013,3019|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|3013,3022|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|3013,3022|false|false|false|C1522577|follow-up|follow-up
Procedure|Health Care Activity|Hospital Course|3013,3027|false|false|false|C3899107|Follow-Up Care|follow-up care
Event|Activity|Hospital Course|3023,3027|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|3023,3027|false|false|false|||care
Finding|Finding|Hospital Course|3023,3027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|3023,3027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Body Substance|Hospital Course|3034,3041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3034,3041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3034,3041|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3052,3061|false|false|false|||readiness
Finding|Finding|Hospital Course|3052,3061|false|false|false|C1318963|Readiness|readiness
Attribute|Clinical Attribute|Hospital Course|3052,3075|false|false|false|C1320402|Readiness for discharge|readiness for discharge
Finding|Finding|Hospital Course|3052,3075|false|false|false|C2314972|Ready for discharge|readiness for discharge
Event|Event|Hospital Course|3066,3075|false|false|false|||discharge
Finding|Body Substance|Hospital Course|3066,3075|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|3066,3075|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|3066,3075|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|3066,3075|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Hospital Course|3080,3091|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3080,3091|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|3080,3091|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|3080,3091|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|3080,3104|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|3095,3104|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|3095,3104|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|3123,3133|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|3123,3133|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|3123,3138|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|3134,3138|false|false|false|||list
Finding|Intellectual Product|Hospital Course|3134,3138|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|3142,3150|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|3155,3163|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|3155,3163|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|3155,3163|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|3155,3163|false|false|false|||complete
Finding|Functional Concept|Hospital Course|3155,3163|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|3155,3163|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3168,3175|false|false|false|C0733877|Lactaid|Lactaid
Drug|Enzyme|Hospital Course|3168,3175|false|false|false|C0733877|Lactaid|Lactaid
Drug|Pharmacologic Substance|Hospital Course|3168,3175|false|false|false|C0733877|Lactaid|Lactaid
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3177,3184|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Drug|Enzyme|Hospital Course|3177,3184|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Drug|Pharmacologic Substance|Hospital Course|3177,3184|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Event|Event|Hospital Course|3177,3184|false|false|false|||lactase
Finding|Gene or Genome|Hospital Course|3177,3184|false|false|false|C1416808|LCT gene|lactase
Anatomy|Body Space or Junction|Hospital Course|3197,3201|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|3197,3201|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|3197,3201|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|3197,3201|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|3202,3207|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|3208,3211|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biologically Active Substance|Hospital Course|3216,3223|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|3216,3223|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|3216,3223|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|3216,3223|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|3216,3223|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|3216,3223|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|3216,3223|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|3216,3223|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Organic Chemical|Hospital Course|3216,3231|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Pharmacologic Substance|Hospital Course|3216,3231|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Organic Chemical|Hospital Course|3224,3231|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Drug|Pharmacologic Substance|Hospital Course|3224,3231|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Event|Event|Hospital Course|3224,3231|false|false|false|||Citrate
Procedure|Laboratory Procedure|Hospital Course|3224,3231|false|false|false|C0201956|Citrate measurement|Citrate
Drug|Biologically Active Substance|Hospital Course|3237,3244|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|3237,3244|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|3237,3244|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|3237,3244|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|3237,3244|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|3237,3244|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|3237,3244|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|3237,3244|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|3237,3252|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|3237,3252|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|3245,3252|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|3245,3252|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|3245,3252|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|3245,3252|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|3253,3260|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|3253,3260|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|3253,3260|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|3253,3260|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|3253,3263|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|3253,3263|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|3253,3263|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|3282,3286|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|3282,3286|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|3282,3286|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|3282,3286|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|3287,3292|false|false|false|||DAILY
Event|Event|Hospital Course|3297,3306|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3297,3306|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3297,3318|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|3307,3318|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3307,3318|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|3307,3318|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|3307,3318|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|3324,3337|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|3324,3337|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|3324,3337|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|3324,3337|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|3353,3356|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|3357,3361|false|false|false|C2598155||Pain
Event|Event|Hospital Course|3357,3361|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|3357,3361|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|3357,3361|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|3364,3368|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|3369,3374|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|3369,3374|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|3381,3390|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|3381,3390|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|Hospital Course|3409,3412|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|3413,3425|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|3413,3425|false|false|false|C0009806|Constipation|Constipation
Drug|Organic Chemical|Hospital Course|3432,3440|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|3432,3440|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|3432,3440|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|3432,3447|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|3432,3447|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|3441,3447|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|3441,3447|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|3441,3447|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|3441,3447|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|3441,3447|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|3441,3447|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3458,3461|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3458,3461|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3458,3461|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|3458,3461|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|3458,3461|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|3468,3478|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|3468,3478|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|Hospital Course|3468,3478|false|false|false|||Enoxaparin
Drug|Organic Chemical|Hospital Course|3468,3485|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|3468,3485|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|3479,3485|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|3479,3485|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|3479,3485|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|3479,3485|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|3479,3485|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|3479,3485|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|Hospital Course|3495,3498|false|false|false|||QHS
Drug|Organic Chemical|Hospital Course|3504,3514|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|Hospital Course|3504,3514|false|false|false|C0206460|enoxaparin|enoxaparin
Event|Event|Hospital Course|3504,3514|false|false|false|||enoxaparin
Event|Event|Hospital Course|3576,3583|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|3576,3583|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|3592,3601|false|false|false|C0030049|oxycodone|OxyCODONE
Drug|Pharmacologic Substance|Hospital Course|3592,3601|false|false|false|C0030049|oxycodone|OxyCODONE
Event|Event|Hospital Course|3592,3601|false|false|false|||OxyCODONE
Procedure|Laboratory Procedure|Hospital Course|3592,3601|false|false|false|C0524222|Oxycodone measurement|OxyCODONE
Finding|Idea or Concept|Hospital Course|3603,3612|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|3603,3612|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|3603,3620|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|3613,3620|false|false|false|||Release
Finding|Functional Concept|Hospital Course|3613,3620|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|3613,3620|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3613,3620|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|3636,3639|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|3640,3644|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|3640,3644|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|3640,3644|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|3648,3656|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|3648,3656|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Event|Event|Hospital Course|3658,3660|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|3662,3671|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|3662,3671|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|3662,3671|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|3662,3671|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|3679,3685|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|3689,3697|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|3692,3697|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|3692,3697|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Gene or Genome|Hospital Course|3701,3704|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biomedical or Dental Material|Hospital Course|3715,3721|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|3715,3721|false|false|false|||Tablet
Event|Event|Hospital Course|3723,3730|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|3723,3730|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|3739,3744|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|3739,3744|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3755,3758|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3755,3758|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3755,3758|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|3755,3758|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|3755,3758|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|Hospital Course|3765,3772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|3765,3772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|3765,3772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|3765,3772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|3765,3772|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|3765,3772|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|3765,3772|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|3765,3772|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Organic Chemical|Hospital Course|3765,3780|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Pharmacologic Substance|Hospital Course|3765,3780|false|false|false|C0108101|calcium citrate|Calcium Citrate
Drug|Organic Chemical|Hospital Course|3773,3780|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Drug|Pharmacologic Substance|Hospital Course|3773,3780|false|false|false|C0008857;C0376259|Citrates;citrate|Citrate
Event|Event|Hospital Course|3773,3780|false|false|false|||Citrate
Procedure|Laboratory Procedure|Hospital Course|3773,3780|false|false|false|C0201956|Citrate measurement|Citrate
Drug|Biologically Active Substance|Hospital Course|3786,3793|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|3786,3793|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|3786,3793|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|3786,3793|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|3786,3793|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|3786,3793|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|3786,3793|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|3786,3793|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|3786,3801|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|3786,3801|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|3794,3801|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|3794,3801|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|3794,3801|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|3794,3801|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|3802,3809|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|3802,3809|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|3802,3809|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|3802,3809|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|3802,3812|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|3802,3812|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|3802,3812|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|3831,3835|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|3831,3835|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|3831,3835|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|3831,3835|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|3836,3841|false|false|false|||DAILY
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3848,3855|false|false|false|C0733877|Lactaid|Lactaid
Drug|Enzyme|Hospital Course|3848,3855|false|false|false|C0733877|Lactaid|Lactaid
Drug|Pharmacologic Substance|Hospital Course|3848,3855|false|false|false|C0733877|Lactaid|Lactaid
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3857,3864|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Drug|Enzyme|Hospital Course|3857,3864|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Drug|Pharmacologic Substance|Hospital Course|3857,3864|false|false|false|C0083183;C1256865|GLB1 protein, human;lactase|lactase
Event|Event|Hospital Course|3857,3864|false|false|false|||lactase
Finding|Gene or Genome|Hospital Course|3857,3864|false|false|false|C1416808|LCT gene|lactase
Anatomy|Body Space or Junction|Hospital Course|3877,3881|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|3877,3881|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|3877,3881|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|3877,3881|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|3882,3887|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|3888,3891|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|3898,3911|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|3898,3911|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|3898,3911|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|3898,3911|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|3914,3917|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|3914,3917|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|3934,3941|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|3934,3941|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|3934,3941|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|3934,3943|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|3934,3943|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|3934,3943|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|3934,3943|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|3934,3943|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|3942,3943|false|false|false|||D
Event|Event|Hospital Course|3948,3952|false|false|false|||UNIT
Event|Event|Hospital Course|3967,3976|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3967,3976|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3967,3976|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3967,3976|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3967,3976|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|3967,3988|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|3967,3988|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|3977,3988|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|3977,3988|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|3977,3988|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|3990,3994|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|3990,3994|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|3990,3994|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|3990,3994|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|4000,4007|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|4000,4007|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|4010,4018|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|4010,4018|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|4026,4035|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|4026,4035|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4026,4035|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4026,4035|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4026,4035|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|4026,4045|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|4036,4045|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|4036,4045|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|4036,4045|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|4036,4045|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|4036,4045|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|4047,4051|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Anatomical Abnormality|Hospital Course|4052,4058|false|false|false|C0042282|Valgus deformity|valgus
Event|Event|Hospital Course|4052,4058|false|false|false|||valgus
Disorder|Disease or Syndrome|Hospital Course|4059,4067|false|false|false|C0040456|Impacted tooth|impacted
Event|Event|Hospital Course|4059,4067|false|false|false|||impacted
Finding|Functional Concept|Hospital Course|4059,4067|false|false|false|C0333125|Impacted|impacted
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4068,4075|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4068,4080|false|false|false|C0015815|Structure of neck of femur|femoral neck
Disorder|Injury or Poisoning|Hospital Course|4068,4089|false|false|false|C0015806|Femoral Neck Fractures|femoral neck fracture
Anatomy|Body Location or Region|Hospital Course|4076,4080|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|4076,4080|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|4076,4080|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Disorder|Injury or Poisoning|Hospital Course|4076,4089|false|false|false|C0262414|Fracture of cervical spine|neck fracture
Disorder|Injury or Poisoning|Hospital Course|4081,4089|false|false|false|C0016658|Fracture|fracture
Event|Event|Hospital Course|4081,4089|false|false|false|||fracture
Disorder|Disease or Syndrome|Discharge Condition|4119,4122|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Discharge Condition|4119,4122|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Discharge Condition|4119,4122|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Discharge Condition|4119,4122|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Discharge Condition|4119,4122|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Discharge Condition|4119,4122|false|false|false|||NAD
Finding|Finding|Discharge Condition|4119,4122|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|Discharge Condition|4124,4125|false|false|false|||A
Event|Event|Discharge Condition|4130,4133|false|false|false|||LLE
Anatomy|Body Location or Region|Discharge Condition|4135,4143|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|Discharge Condition|4135,4143|false|false|false|C0332803|Surgical wound|Incision
Event|Event|Discharge Condition|4135,4143|false|false|false|||Incision
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|4135,4143|false|false|false|C0184898|Surgical incisions|Incision
Finding|Finding|Discharge Condition|4144,4148|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Condition|4149,4161|false|false|false|||approximated
Drug|Biomedical or Dental Material|Discharge Condition|4163,4171|false|false|false|C1705365|Dressing Dosage Form|Dressing
Event|Event|Discharge Condition|4163,4171|false|false|false|||Dressing
Finding|Daily or Recreational Activity|Discharge Condition|4163,4171|false|false|false|C0518459;C1305428|Ability to dress|Dressing
Finding|Finding|Discharge Condition|4163,4171|false|false|false|C0518459;C1305428|Ability to dress|Dressing
Procedure|Health Care Activity|Discharge Condition|4163,4171|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|Dressing
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|4163,4171|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|Dressing
Event|Activity|Discharge Condition|4172,4177|false|false|false|C1947930|Cleaning (activity)|clean
Disorder|Disease or Syndrome|Discharge Condition|4187,4192|false|false|false|C4049262|Febrile infection related epilepsy syndrome|Fires
Event|Event|Discharge Condition|4187,4192|false|false|false|||Fires
Event|Event|Discharge Condition|4187,4192|false|false|false|C0016141|fire disaster|Fires
Phenomenon|Natural Phenomenon or Process|Discharge Condition|4187,4192|false|false|false|C0700614|Fire (physical force)|Fires
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4208,4211|false|false|false|C1522376;C4283742|Ceramide Glucosyltransferase, human;GCLC protein, human|GCS
Drug|Enzyme|Family Medical History|4208,4211|false|false|false|C1522376;C4283742|Ceramide Glucosyltransferase, human;GCLC protein, human|GCS
Event|Event|Family Medical History|4208,4211|false|false|false|||GCS
Finding|Gene or Genome|Family Medical History|4208,4211|false|false|false|C1415097;C1421319;C1704697;C4283933|GCLC gene;GCLC wt Allele;UGCG gene;UGCG wt Allele|GCS
Event|Event|Family Medical History|4224,4237|false|false|false|||distributions
Attribute|Clinical Attribute|Family Medical History|4246,4251|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|Family Medical History|4246,4251|false|false|false|||pulse
Finding|Physiologic Function|Family Medical History|4246,4251|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|Family Medical History|4246,4251|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|Family Medical History|4246,4251|false|false|false|C0034107|Pulse taking|pulse
Attribute|Clinical Attribute|Discharge Instructions|4294,4306|false|false|false|C3263700||INSTRUCTIONS
Event|Event|Discharge Instructions|4294,4306|false|false|false|||INSTRUCTIONS
Finding|Intellectual Product|Discharge Instructions|4294,4306|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|INSTRUCTIONS
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4313,4332|false|false|false|C1136201|Orthopedic Surgical Procedures|ORTHOPAEDIC SURGERY
Event|Event|Discharge Instructions|4325,4332|false|false|false|||SURGERY
Finding|Finding|Discharge Instructions|4325,4332|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Discharge Instructions|4325,4332|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Discharge Instructions|4325,4332|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4325,4332|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Idea or Concept|Discharge Instructions|4353,4361|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4366,4384|false|false|false|C0162439;C1136201|Orthopedic Rehabilitation Surgery;Orthopedic Surgical Procedures|orthopedic surgery
Event|Event|Discharge Instructions|4377,4384|false|false|false|||surgery
Finding|Finding|Discharge Instructions|4377,4384|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|4377,4384|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|4377,4384|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4377,4384|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|4392,4398|false|false|false|||normal
Event|Event|Discharge Instructions|4403,4407|false|false|false|||feel
Finding|Mental Process|Discharge Instructions|4403,4407|false|false|false|C1527305|Feelings|feel
Finding|Finding|Discharge Instructions|4403,4413|false|false|false|C0849970;C3539029|Feel Tired question;Feeling tired|feel tired
Finding|Intellectual Product|Discharge Instructions|4403,4413|false|false|false|C0849970;C3539029|Feel Tired question;Feeling tired|feel tired
Event|Event|Discharge Instructions|4408,4413|false|false|false|||tired
Finding|Finding|Discharge Instructions|4408,4413|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|Discharge Instructions|4408,4413|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|Discharge Instructions|4408,4413|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|Discharge Instructions|4418,4424|false|false|false|||washed
Finding|Finding|Discharge Instructions|4430,4443|false|false|false|C0241311|post operative (finding)|after surgery
Event|Event|Discharge Instructions|4436,4443|false|false|false|||surgery
Finding|Finding|Discharge Instructions|4436,4443|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|4436,4443|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|4436,4443|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4436,4443|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|4454,4461|false|false|false|||feeling
Finding|Mental Process|Discharge Instructions|4454,4461|false|false|false|C1527305|Feelings|feeling
Event|Event|Discharge Instructions|4470,4477|false|false|false|||improve
Finding|Intellectual Product|Discharge Instructions|4505,4509|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Discharge Instructions|4514,4520|false|false|false|||Resume
Finding|Functional Concept|Discharge Instructions|4514,4520|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Idea or Concept|Discharge Instructions|4514,4520|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Finding|Intellectual Product|Discharge Instructions|4514,4520|false|false|false|C1550028;C1880201;C3242342|Curriculum Vitae;Resume - Remote control command;resume - DataOperation|Resume
Event|Activity|Discharge Instructions|4534,4544|false|false|false|C0441655|Activities|activities
Event|Event|Discharge Instructions|4534,4544|false|false|false|||activities
Finding|Finding|Discharge Instructions|4534,4544|false|false|false|C2239122|activities (history)|activities
Event|Event|Discharge Instructions|4548,4557|false|false|false|||tolerated
Event|Event|Discharge Instructions|4570,4576|false|false|false|||follow
Attribute|Clinical Attribute|Discharge Instructions|4583,4589|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|4583,4589|false|false|false|||weight
Finding|Finding|Discharge Instructions|4583,4589|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|4583,4589|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|4583,4589|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|4598,4609|false|false|false|||precautions
Finding|Conceptual Entity|Discharge Instructions|4598,4609|false|false|false|C1882442|Precaution|precautions
Disorder|Disease or Syndrome|Discharge Instructions|4626,4631|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Activity|Discharge Instructions|4634,4642|false|false|false|C0441655|Activities|ACTIVITY
Finding|Daily or Recreational Activity|Discharge Instructions|4634,4642|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|Discharge Instructions|4634,4642|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Attribute|Clinical Attribute|Discharge Instructions|4647,4653|false|false|false|C0944911||WEIGHT
Event|Event|Discharge Instructions|4647,4653|false|false|false|||WEIGHT
Finding|Finding|Discharge Instructions|4647,4653|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Finding|Sign or Symptom|Discharge Instructions|4647,4653|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|WEIGHT
Procedure|Health Care Activity|Discharge Instructions|4647,4653|false|false|false|C1305866|Weighing patient|WEIGHT
Event|Event|Discharge Instructions|4665,4678|false|false|false|||Weightbearing
Event|Event|Discharge Instructions|4682,4691|false|false|false|||tolerated
Finding|Functional Concept|Discharge Instructions|4692,4696|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4692,4712|false|false|false|C0230416|Left lower extremity|left lower extremity
Anatomy|Body Location or Region|Discharge Instructions|4697,4702|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Discharge Instructions|4697,4702|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4697,4712|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4703,4712|false|false|false|C0015385|Limb structure|extremity
Event|Event|Medications|4733,4737|false|false|false|||Take
Drug|Organic Chemical|Medications|4738,4745|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|4738,4745|false|false|false|C0699142|Tylenol|Tylenol
Drug|Amino Acid, Peptide, or Protein|Medications|4775,4780|false|false|false|C1743089|CLOCK protein, human|clock
Drug|Enzyme|Medications|4775,4780|false|false|false|C1743089|CLOCK protein, human|clock
Event|Event|Medications|4775,4780|false|false|false|||clock
Finding|Gene or Genome|Medications|4775,4780|false|false|false|C1413503|CLOCK gene|clock
Drug|Pharmacologic Substance|Medications|4794,4810|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|Medications|4803,4810|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Medications|4803,4810|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Pharmacologic Substance|Medications|4811,4821|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|4811,4821|false|false|false|||medication
Finding|Intellectual Product|Medications|4811,4821|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Medications|4833,4842|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Medications|4833,4842|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Medications|4833,4842|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Medications|4833,4842|false|false|false|C0524222|Oxycodone measurement|oxycodone
Event|Event|Medications|4846,4852|false|false|false|||needed
Attribute|Clinical Attribute|Medications|4867,4871|false|false|false|C2598155||pain
Event|Event|Medications|4867,4871|false|false|false|||pain
Finding|Functional Concept|Medications|4867,4871|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|4867,4871|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|4880,4884|false|false|false|||wean
Finding|Finding|Medications|4880,4884|false|false|false|C0043084|Weaning|wean
Drug|Pharmacologic Substance|Medications|4895,4905|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|4895,4905|false|false|false|||medication
Finding|Intellectual Product|Medications|4895,4905|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|Medications|4911,4915|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Medications|4939,4946|false|false|false|||example
Finding|Conceptual Entity|Medications|4939,4946|false|false|false|C1707959|Example|example
Event|Event|Medications|4958,4962|false|false|false|||wean
Event|Event|Medications|4969,4973|false|false|false|||Take
Drug|Biomedical or Dental Material|Medications|4976,4982|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|4976,4982|false|false|false|||tablet
Event|Event|Medications|5000,5006|false|false|false|||needed
Finding|Idea or Concept|Medications|5011,5014|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5011,5014|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5016,5020|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Medications|5023,5029|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|5023,5029|false|false|false|||tablet
Event|Event|Medications|5047,5053|false|false|false|||needed
Finding|Idea or Concept|Medications|5058,5061|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5058,5061|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5063,5067|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Medications|5070,5076|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|5070,5076|false|false|false|||tablet
Event|Event|Medications|5094,5100|false|false|false|||needed
Finding|Idea or Concept|Medications|5105,5108|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5105,5108|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5110,5114|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Medications|5117,5123|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|5117,5123|false|false|false|||tablet
Event|Event|Medications|5141,5147|false|false|false|||needed
Finding|Intellectual Product|Medications|5159,5163|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Medications|5166,5172|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|5166,5172|false|false|false|||tablet
Event|Event|Medications|5191,5197|false|false|false|||needed
Finding|Idea or Concept|Medications|5202,5205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5202,5205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5207,5211|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Medications|5214,5220|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Medications|5214,5220|false|false|false|||tablet
Finding|Intellectual Product|Medications|5221,5226|false|false|false|C1720374|Every - dosing instruction fragment|every
Event|Event|Medications|5245,5251|false|false|false|||needed
Finding|Idea or Concept|Medications|5256,5259|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5256,5259|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Medications|5263,5267|false|false|false|C1720594|Then - dosing instruction fragment|Then
Event|Event|Medications|5268,5276|false|false|false|||continue
Drug|Organic Chemical|Medications|5282,5289|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|5282,5289|false|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|5282,5289|false|false|false|||Tylenol
Attribute|Clinical Attribute|Medications|5294,5298|false|false|false|C2598155||pain
Event|Event|Medications|5294,5298|false|false|false|||pain
Finding|Functional Concept|Medications|5294,5298|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|5294,5298|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|5313,5317|true|false|false|||stop
Drug|Organic Chemical|Medications|5322,5329|true|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Medications|5322,5329|true|false|false|C0699142|Tylenol|Tylenol
Event|Event|Medications|5322,5329|true|false|false|||Tylenol
Drug|Hazardous or Poisonous Substance|Medications|5355,5363|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Medications|5355,5363|false|false|false|C0027415|Narcotics|narcotic
Event|Event|Medications|5355,5363|false|false|false|||narcotic
Drug|Pharmacologic Substance|Medications|5365,5375|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|5365,5375|false|false|false|||medication
Finding|Intellectual Product|Medications|5365,5375|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Functional Concept|Medications|5387,5392|false|false|false|C1442792|State|state
Event|Event|Medications|5393,5404|false|false|false|||regulations
Event|Governmental or Regulatory Activity|Medications|5393,5404|false|false|false|C0851285|Regulation|regulations
Event|Event|Medications|5413,5420|false|false|false|||limited
Finding|Intellectual Product|Medications|5428,5434|false|false|false|C1561574|Amount class - Amount|amount
Drug|Hazardous or Poisonous Substance|Medications|5439,5448|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Medications|5439,5448|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Medications|5456,5465|false|false|false|||prescribe
Event|Event|Medications|5498,5505|false|false|false|||contact
Event|Event|Medications|5510,5516|false|false|false|||office
Finding|Idea or Concept|Medications|5510,5516|false|false|false|C1549636|Address type - Office|office
Event|Event|Medications|5520,5523|false|false|false|||set
Event|Activity|Medications|5530,5541|false|false|false|C0003629|Appointments|appointment
Event|Event|Medications|5530,5541|false|false|false|||appointment
Event|Event|Medications|5561,5567|true|false|false|||refill
Event|Event|Medications|5573,5577|true|false|false|||type
Finding|Gene or Genome|Medications|5573,5577|true|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Medications|5573,5577|true|true|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Attribute|Clinical Attribute|Medications|5581,5585|true|false|false|C2598155||pain
Finding|Functional Concept|Medications|5581,5585|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|5581,5585|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Medications|5586,5596|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|5586,5596|true|false|false|||medication
Finding|Intellectual Product|Medications|5586,5596|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Medications|5606,5611|false|false|false|||phone
Finding|Idea or Concept|Medications|5606,5611|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Intellectual Product|Medications|5606,5611|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Drug|Hazardous or Poisonous Substance|Medications|5620,5628|false|false|false|C0027415|Narcotics|Narcotic
Drug|Pharmacologic Substance|Medications|5620,5628|false|false|false|C0027415|Narcotics|Narcotic
Attribute|Clinical Attribute|Medications|5629,5633|false|false|false|C2598155||pain
Event|Event|Medications|5629,5633|false|false|false|||pain
Finding|Functional Concept|Medications|5629,5633|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|5629,5633|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Medications|5629,5643|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|Medications|5629,5643|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|Medications|5629,5643|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|Medications|5634,5643|false|false|false|||relievers
Event|Event|Medications|5654,5666|false|false|false|||constipation
Finding|Sign or Symptom|Medications|5654,5666|false|false|false|C0009806|Constipation|constipation
Event|Event|Medications|5683,5688|false|false|false|||drink
Drug|Inorganic Chemical|Medications|5710,5715|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Medications|5710,5715|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Medications|5710,5715|false|false|false|||water
Finding|Intellectual Product|Medications|5710,5715|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Medications|5710,5715|false|false|false|C0020311|Hydrotherapy|water
Event|Event|Medications|5726,5734|false|false|false|||continue
Event|Event|Medications|5736,5745|false|false|false|||following
Anatomy|Body Part, Organ, or Organ Component|Medications|5750,5755|false|false|false|C0021853|Intestines|bowel
Procedure|Health Care Activity|Medications|5750,5763|false|false|false|C5979615|Bowel Regimen|bowel regimen
Event|Event|Medications|5756,5763|false|false|false|||regimen
Finding|Intellectual Product|Medications|5756,5763|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Medications|5756,5763|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|Medications|5767,5773|false|false|false|||stated
Drug|Pharmacologic Substance|Medications|5782,5792|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Medications|5782,5792|false|false|false|||medication
Finding|Intellectual Product|Medications|5782,5792|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Attribute|Clinical Attribute|Medications|5794,5806|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Medications|5794,5806|false|false|false|||prescription
Finding|Intellectual Product|Medications|5794,5806|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Medications|5794,5806|false|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|Medications|5794,5811|false|false|false|C2741652||prescription list
Finding|Intellectual Product|Medications|5794,5811|false|false|false|C3533331|Prescription list|prescription list
Event|Event|Medications|5807,5811|false|false|false|||list
Finding|Intellectual Product|Medications|5807,5811|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Disorder|Disease or Syndrome|Medications|5819,5823|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Event|Event|Medications|5819,5823|false|false|false|||meds
Finding|Intellectual Product|Medications|5819,5823|false|false|false|C4284232|Medications|meds
Drug|Organic Chemical|Medications|5825,5830|false|false|false|C3489575|sennosides, USP|senna
Drug|Pharmacologic Substance|Medications|5825,5830|false|false|false|C3489575|sennosides, USP|senna
Event|Event|Medications|5825,5830|false|false|false|||senna
Drug|Organic Chemical|Medications|5832,5838|false|false|false|C0282139|Colace|colace
Drug|Pharmacologic Substance|Medications|5832,5838|false|false|false|C0282139|Colace|colace
Event|Event|Medications|5832,5838|false|false|false|||colace
Drug|Organic Chemical|Medications|5840,5847|false|false|false|C0876088|Miralax|miralax
Drug|Pharmacologic Substance|Medications|5840,5847|false|false|false|C0876088|Miralax|miralax
Event|Event|Medications|5840,5847|false|false|false|||miralax
Drug|Hazardous or Poisonous Substance|Medications|5863,5870|true|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Medications|5863,5870|true|false|false|C0702263|Counter brand of Terbufos|counter
Event|Event|Medications|5863,5870|true|false|false|||counter
Event|Event|Medications|5882,5890|true|false|false|||obtained
Event|Event|Medications|5898,5906|true|false|false|||pharmacy
Finding|Intellectual Product|Medications|5898,5906|true|false|false|C1547997;C3244303|Diagnostic Service Section ID - Pharmacy;Pharmacy domain|pharmacy
Procedure|Health Care Activity|Medications|5898,5906|true|false|false|C0031321|Pharmaceutical Services|pharmacy
Event|Event|Medications|5921,5926|true|false|false|||drink
Drug|Organic Chemical|Medications|5927,5934|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Medications|5927,5934|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Medications|5927,5934|true|false|false|||alcohol
Finding|Intellectual Product|Medications|5927,5934|true|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|Medications|5936,5941|true|false|false|||drive
Finding|Functional Concept|Medications|5944,5949|true|false|false|C1513492|motor movement|motor
Drug|Biomedical or Dental Material|Medications|5950,5957|true|false|false|C0042444|Drug vehicle|vehicle
Event|Event|Medications|5950,5957|true|false|false|||vehicle
Event|Event|Medications|5962,5969|false|false|false|||operate
Finding|Functional Concept|Medications|5962,5969|false|false|false|C3242339|operate|operate
Disorder|Injury or Poisoning|Medications|5971,5980|false|false|false|C0337246|Contact with machinery|machinery
Event|Event|Medications|5971,5980|false|false|false|||machinery
Event|Event|Medications|5987,5993|false|false|false|||taking
Drug|Hazardous or Poisonous Substance|Medications|5994,6002|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Medications|5994,6002|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Medications|6003,6007|false|false|false|C2598155||pain
Event|Event|Medications|6003,6007|false|false|false|||pain
Finding|Functional Concept|Medications|6003,6007|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Medications|6003,6007|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Medications|6003,6017|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Organic Chemical|Medications|6003,6017|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Drug|Pharmacologic Substance|Medications|6003,6017|false|false|false|C0002771;C0722425|Analgesics;Pain Relieve brand of acetaminophen|pain relievers
Event|Event|Medications|6008,6017|false|false|false|||relievers
Event|Event|Medications|6032,6036|false|false|false|||take
Attribute|Clinical Attribute|Medications|6041,6052|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|6041,6052|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|6041,6052|false|false|false|||medications
Finding|Intellectual Product|Medications|6041,6052|false|false|false|C4284232|Medications|medications
Event|Event|Medications|6056,6066|false|false|false|||prescribed
Event|Event|Medications|6076,6086|false|false|false|||physicians
Event|Event|Medications|6090,6099|false|false|false|||discharge
Finding|Body Substance|Medications|6090,6099|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Medications|6090,6099|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Medications|6090,6099|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Medications|6090,6099|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Medications|6107,6115|false|false|false|||Continue
Finding|Idea or Concept|Medications|6120,6124|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Medications|6120,6124|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Medications|6120,6124|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Medications|6125,6136|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Medications|6125,6136|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Medications|6125,6136|false|false|false|||medications
Finding|Intellectual Product|Medications|6125,6136|false|false|false|C4284232|Medications|medications
Event|Event|Medications|6158,6168|false|false|false|||instructed
Event|Event|Medications|6172,6176|false|false|false|||stop
Attribute|Clinical Attribute|Medications|6185,6192|false|false|false|C5444295||surgeon
Event|Event|Medications|6201,6216|false|false|false|||ANTICOAGULATION
Finding|Finding|Medications|6201,6216|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Finding|Physiologic Function|Medications|6201,6216|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|ANTICOAGULATION
Procedure|Therapeutic or Preventive Procedure|Medications|6201,6216|false|false|false|C0003281|Anticoagulation Therapy|ANTICOAGULATION
Event|Event|Medications|6227,6231|false|false|false|||take
Drug|Organic Chemical|Medications|6233,6240|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Medications|6233,6240|false|false|false|C0728963|Lovenox|Lovenox
Event|Event|Medications|6233,6240|false|false|false|||Lovenox
Procedure|Health Care Activity|Medications|6261,6269|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|6270,6282|false|false|false|C3263700||Instructions
Event|Event|Medications|6270,6282|false|false|false|||Instructions
Finding|Intellectual Product|Medications|6270,6282|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

