CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Chest pressure|Finding|false|false||chest pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|PMH - past medical history|Finding|false|false||past medical history
null|Medical History|Finding|false|false||past medical historynull|Medical History|Finding|false|false||medical history ofnull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Chest pressure|Finding|false|false||chest pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Initially|Time|false|false||initiallynull|GLAUCOMA, NORMAL TENSION, SUSCEPTIBILITY TO|Finding|false|false||NTG
null|OPA1 wt Allele|Finding|false|false||NTG
null|OPA1 gene|Finding|false|false||NTGnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Short menstrual periods|Finding|false|false||short periodnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Radiating to|Finding|false|false||radiatednull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|Both upper arms|Anatomy|false|false||both armsnull|Alveolar rhabdomyosarcoma|Disorder|false|false||armsnull|Adherence to Refills and Medications Scale|Finding|false|false||arms
null|KIDINS220 gene|Finding|false|false||armsnull|Upper arm|Anatomy|false|false||armsnull|null|Attribute|false|false||armsnull|Increased sweating|Finding|false|false||diaphoresisnull|Associated with|Modifier|true|false||associatednull|Nausea|Finding|true|false||nauseanull|null|Attribute|true|false||nauseanull|Vomiting|Finding|true|false||vomitingnull|Lightheadedness|Finding|true|false||lightheadednessnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Dyspnea|Finding|false|false||SOBnull|Recent|Time|false|false||recentnull|Pneumonia|Disorder|false|false||pneumonianull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|week|Time|false|false||weeksnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|null|Finding|true|false||dyspnea
null|Dyspnea|Finding|true|false||dyspneanull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Very|Modifier|false|false||verynull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|New LBBB|Finding|false|false||new LBBBnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Elevation|Modifier|false|false||elevationsnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Catheterization|Procedure|false|false||cathnull|AML Lab Table|Finding|false|false||lab
null|LAT2 gene|Finding|false|false||lab
null|EWS Lab Table|Finding|false|false||labnull|Laboratory|Device|false|false||labnull|Labrador retriever|Entity|false|false||lab
null|Laboratory|Entity|false|false||labnull|Catheterization|Procedure|false|false||Cathnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Scalable Vector Graphics|Entity|false|false||SVGnull|Native (qualifier value)|Finding|false|false||Nativenull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Concern|Finding|false|false||concernnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Dissecting hemorrhage|Finding|false|false||dissectionnull|Tissue Dissection|Procedure|false|false||dissectionnull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Diminutive|Finding|false|false||diminutivenull|Septal|Modifier|false|false||septalnull|diagnosis aspects|Finding|false|false||diagnull|Diagnosis|Procedure|false|false||diagnull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Androgen Binding Protein|Drug|false|false||SBP
null|Androgen Binding Protein|Drug|false|false||SBPnull|CCHCR1 wt Allele|Finding|false|false||SBP
null|SHBG wt Allele|Finding|false|false||SBPnull|Systolic blood pressure measurement|Procedure|false|false||SBPnull|Systolic Pressure|Attribute|false|false||SBPnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Current (present time)|Time|false|false||currentlynull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pain-Free|Drug|false|false||pain freenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|null|Time|true|false||priornull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|true|false||historynull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|true|false||deepnull|Venous thrombosis after immobility|Finding|true|false||venous thrombosis
null|Venous Thrombosis|Finding|true|false||venous thrombosisnull|Veins|Anatomy|true|false||venousnull|Venous|Modifier|true|false||venousnull|Thrombosis|Finding|true|false||thrombosisnull|Pulmonary Embolism|Finding|false|false||pulmonary embolismnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Embolism|Finding|false|false||embolism
null|Embolus|Finding|false|false||embolismnull|Hemorrhage|Finding|false|false||bleedingnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Myalgia|Finding|false|false||myalgiasnull|Arthralgia|Finding|false|false||joint painsnull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Pain|Finding|false|false||painsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Hemoptysis|Finding|false|false||hemoptysisnull|null|Finding|false|false||black stools
null|Melena|Finding|false|false||black stoolsnull|Black - ethnic group (ethnic group)|Subject|false|false||black
null|Black race|Subject|false|false||black
null|African|Subject|false|false||blacknull|Black - Structured Product Labeling Color|Modifier|false|false||black
null|Black color|Modifier|false|false||blacknull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Red stools|Finding|false|false||red stoolsnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|Recent|Time|true|false||recentnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Rigor - Temperature-associated observation|Finding|true|false||rigorsnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Review of systems (procedure)|Procedure|false|false||review of systemsnull|null|Attribute|false|false||review of systems
null|null|Attribute|false|false||review of systemsnull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|System|Finding|false|false||systemsnull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea on exertion|Finding|false|false||dyspnea on exertionnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Exertion|Finding|false|false||exertionnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||paroxysmal nocturnal dyspneanull|Paroxysmal|Time|false|false||paroxysmalnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Ankle edema (finding)|Finding|false|false||ankle edemanull|Lower extremity>Ankle|Anatomy|false|false||ankle
null|Ankle|Anatomy|false|false||ankle
null|Ankle joint structure|Anatomy|false|false||anklenull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Palpitations|Finding|false|false||palpitationsnull|Presyncope or syncope|Finding|false|false||syncope or presyncopenull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Presyncope|Finding|false|false||presyncopenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|cardiac risk factors|Finding|false|false||CARDIAC RISK FACTORSnull|CARD.RISK|Finding|false|false||CARDIAC RISKnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|risk factors - observation list|Finding|false|false||RISK FACTORS
null|risk factors|Finding|false|false||RISK FACTORS
null|History of - risk factor|Finding|false|false||RISK FACTORSnull|null|Attribute|false|false||RISK FACTORSnull|Risk|Finding|false|false||RISKnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Cardiac attachment|Finding|true|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|History of present illness (finding)|Finding|false|false||HISTORY
null|History of previous events|Finding|false|false||HISTORY
null|Historical aspects qualifier|Finding|false|false||HISTORY
null|Medical History|Finding|false|false||HISTORY
null|Concept History|Finding|false|false||HISTORYnull|History|Subject|false|false||HISTORYnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Following|Time|false|false||subsequentnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Percutaneous Coronary Intervention|Procedure|false|false||PERCUTANEOUS CORONARY INTERVENTIONSnull|Percutaneous Route of Drug Administration|Finding|false|false||PERCUTANEOUSnull|Percutaneous|Modifier|false|false||PERCUTANEOUSnull|Heart|Anatomy|false|false||CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Nursing interventions|Procedure|false|false||INTERVENTIONS
null|Intervention regimes|Procedure|false|false||INTERVENTIONSnull|null|Attribute|false|false||INTERVENTIONSnull|Pacing up and down|Finding|true|false||PACINGnull|Disruptive, Impulse Control, and Conduct Disorders|Disorder|true|false||ICD
null|Type II Mucolipidosis|Disorder|true|false||ICDnull|International Classification of Diseases|Finding|true|false||ICD
null|GNPTAB wt Allele|Finding|true|false||ICDnull|Icd Regimen|Procedure|true|false||ICDnull|between lunch and dinner|Time|true|false||ICDnull|PMH - past medical history|Finding|true|false||PAST MEDICAL HISTORY
null|Medical History|Finding|true|false||PAST MEDICAL HISTORYnull|Medical History|Finding|true|false||MEDICAL HISTORYnull|Medical referral type|Finding|true|false||MEDICAL
null|Medical|Finding|true|false||MEDICAL
null|Medical school type|Finding|true|false||MEDICALnull|Medical service|Procedure|true|false||MEDICALnull|Medical History|Finding|true|false||HISTORY
null|History of previous events|Finding|true|false||HISTORY
null|Historical aspects qualifier|Finding|true|false||HISTORY
null|History of present illness (finding)|Finding|true|false||HISTORY
null|Concept History|Finding|true|false||HISTORYnull|History|Subject|true|false||HISTORYnull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Small|LabModifier|false|false||smallnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Infarction|Finding|false|false||infarctnull|Tablet Dosage Form|Drug|false|false||tabnull|Tablet Dosing Unit|LabModifier|false|false||tabnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Daily|Time|false|false||dailynull|Hypercholesterolemia|Disorder|false|false||hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||hypercholesterolemianull|Small|LabModifier|false|false||smallnull|macular|Modifier|false|false||Macularnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Malignant neoplasm of stomach|Disorder|false|false||stomach cancer
null|Stomach Carcinoma|Disorder|false|false||stomach cancernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Malignant Bone Neoplasm|Disorder|false|false||bone cancer
null|Osteosarcoma of bone|Disorder|false|false||bone cancernull|Specimen Type - Bone|Finding|false|false||bone
null|null|Finding|false|false||bonenull|Skeletal bone|Anatomy|false|false||bone
null|XXX bone|Anatomy|false|false||bonenull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Oriented to place|Finding|false|false||Orientednull|Orientation, Spatial|Modifier|false|false||Orientednull|Mood (psychological function)|Finding|false|false||Mood
null|mood (physical finding)|Finding|false|false||Mood
null|Mood (attribute)|Finding|false|false||Moodnull|null|Attribute|false|false||Moodnull|Appropriate|Modifier|false|false||appropriatenull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false||Scleranull|examination of sclera|Procedure|false|false||Scleranull|Sclera|Anatomy|false|false||Scleranull|Anicteric|Finding|false|false||anictericnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Malignant neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|true|false||Conjunctiva
null|Conjunctival Diseases|Disorder|true|false||Conjunctivanull|Specimen Type - Conjunctiva|Finding|true|false||Conjunctiva
null|null|Finding|true|false||Conjunctivanull|examination of conjunctiva|Procedure|true|false||Conjunctiva
null|Procedure on conjunctiva|Procedure|true|false||Conjunctivanull|Structure of palpebral conjunctiva|Anatomy|true|false||Conjunctiva
null|conjunctiva|Anatomy|true|false||Conjunctivanull|Pink color|Modifier|true|false||pinknull|Pallor of skin|Finding|true|false||pallornull|Cyanosis|Finding|true|false||cyanosisnull|Oral mucous membrane structure|Anatomy|true|false||oral mucosanull|Oral Dosage Form|Drug|true|false||oralnull|Oral Route of Administration|Finding|true|false||oral
null|Oral (intended site)|Finding|true|false||oralnull|Oral cavity|Anatomy|true|false||oralnull|Oral|Modifier|true|false||oralnull|null|Finding|true|false||mucosanull|Mucous Membrane|Anatomy|true|false||mucosanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||Supplenull|Jugular venous pressure|Finding|false|false||JVPnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Point of Maximum Impulse|Finding|false|false||PMI
null|TMEM11 gene|Finding|false|false||PMI
null|PMM2 wt Allele|Finding|false|false||PMI
null|PMM2 gene|Finding|false|false||PMI
null|MPI gene|Finding|false|false||PMInull|Prostate Mechanical Imager|Device|false|false||PMInull|Space of intercostal compartment|Anatomy|false|false||intercostal space
null|Structure of intercostal space|Anatomy|false|false||intercostal spacenull|Intercostal|Modifier|false|false||intercostalnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Midclavicular|Modifier|false|false||midclavicularnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false||linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Cardiac thrill (finding)|Finding|true|false||thrillsnull|hoist [device]|Device|true|false||liftsnull|Lung|Anatomy|false|false||LUNGSnull|Deformity of chest wall|Disorder|true|false||chest wall deformitiesnull|Chest wall structure|Anatomy|true|false||chest wall
null|Chest>Chest wall|Anatomy|true|false||chest wallnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Walls of a building|Device|true|false||wallnull|Congenital Abnormality|Disorder|true|false||deformitiesnull|deformities qualifier|Modifier|true|false||deformitiesnull|Congenital scoliosis|Disorder|true|false||scoliosis
null|null|Disorder|true|false||scoliosis
null|Acquired scoliosis|Disorder|true|false||scoliosisnull|Kyphosis deformity of spine|Disorder|true|false||kyphosis
null|Acquired kyphosis|Disorder|true|false||kyphosis
null|Congenital kyphosis|Disorder|true|false||kyphosisnull|kyphosis|Finding|true|false||kyphosisnull|Respiratory, thoracic and mediastinal disorders|Disorder|true|false||Respnull|Respiratory rate|Attribute|true|false||Respnull|Unlabored|Finding|true|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|true|false||muscle
null|Muscle Tissue|Anatomy|true|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Cancer/Testis Antigen|Drug|true|false||CTAnull|PCYT1A wt Allele|Finding|true|false||CTA
null|CERNA3 gene|Finding|true|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|true|false||CTAnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Wheezing|Finding|true|false||wheezesnull|Rhonchi|Finding|true|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Emotional tenderness|Finding|true|false||tenderness
null|Sore to touch|Finding|true|false||tendernessnull|Absence of Biallelic TCRgamma Deletion|Disorder|true|false||Abdnull|ABD (body structure)|Anatomy|true|false||Abd
null|Abdomen|Anatomy|true|false||Abdnull|Procedure on aorta|Procedure|true|false||aortanull|Chest+Abdomen>Aorta|Anatomy|true|false||aorta
null|Aorta|Anatomy|true|false||aortanull|Palpation|Procedure|true|false||palpationnull|Bruit|Finding|true|false||bruitsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Femur|Anatomy|false|false||Femoralnull|Foreskin of penis|Anatomy|false|false||sheathnull|Condoms, Male|Device|false|false||sheathnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pelvis>Groin|Anatomy|false|false||groin
null|Inguinal region|Anatomy|false|false||groin
null|Inguinal part of abdomen|Anatomy|false|false||groinnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|Stasis dermatitis|Disorder|true|false||stasis dermatitisnull|Stasis|Finding|true|false||stasisnull|Dermatitis|Disorder|true|false||dermatitisnull|Ulcer|Finding|true|false||ulcersnull|Scar Tissue|Finding|true|false||scars
null|Cicatrix|Finding|true|false||scarsnull|Xanthoma|Disorder|true|false||xanthomasnull|null|Drug|false|false||PULSESnull|Physiologic pulse|Finding|false|false||PULSESnull|Pulse taking|Procedure|false|false||PULSESnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Carotid Arteries|Anatomy|false|false||Carotidnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|New LBBB|Finding|false|false||new LBBBnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Left Bundle-Branch Block|Disorder|false|false||LBBBnull|null|Lab|false|false||LBBBnull|SULT1E1 wt Allele|Finding|false|false||STE
null|SULT1E1 gene|Finding|false|false||STEnull|Lead Device|Device|false|false||leadsnull|Telemetry|Procedure|false|false||TELEMETRYnull|null|Finding|false|false||NSR
null|Neutral Sidebent Rotated|Finding|false|false||NSRnull|Echocardiography|Procedure|false|false||ECHOCARDIOGRAMnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|Trophoblastic tumor, epithelioid|Disorder|false|false||ETTnull|Cardiac Catheterization Procedures|Procedure|false|false||CARDIAC CATHnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Catheterization|Procedure|false|false||CATHnull|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCA
null|levomefolate calcium|Drug|false|false||LMCAnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Occluded|Finding|false|false||Occluded
null|Obstruction|Finding|false|false||Occludednull|Difficult (qualifier value)|Finding|false|false||difficultnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Distal Resection Margin|Attribute|false|false||Distalnull|Distal (qualifier value)|Modifier|false|false||Distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Diffuse|Modifier|false|false||diffusenull|Diseased|Modifier|false|false||diseasednull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Methylcytosine Dioxygenase TET1|Drug|false|false||LCX
null|Methylcytosine Dioxygenase TET1|Drug|false|false||LCXnull|TET1 wt Allele|Finding|false|false||LCX
null|TET1 gene|Finding|false|false||LCXnull|Occluded|Finding|false|false||Occluded
null|Obstruction|Finding|false|false||Occludednull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Catheterization|Procedure|false|false||catheterizationnull|Multiple Pulmonary Nodules|Finding|false|false||multiple pulmonary nodulesnull|Numerous|LabModifier|false|false||multiplenull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|ST segment elevation myocardial infarction|Disorder|false|false||STEMInull|ST Elevation Myocardial Infarction by ECG Finding|Finding|false|false||STEMInull|Risk|Finding|false|false||risknull|Score|Finding|false|false||scorenull|Risk|Finding|false|false||risknull|14 days|Time|false|false||14 daysnull|day|Time|false|false||daysnull|Aspects of mortality statistics|LabModifier|false|false||mortality
null|Mortality Vital Statistics|LabModifier|false|false||mortalitynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Certification patient type - Urgent|Finding|false|false||urgent
null|Admission Type - Urgent|Finding|false|false||urgent
null|Triage Code - Urgent|Finding|false|false||urgent
null|Visit Priority Code - Urgent|Finding|false|false||urgentnull|Act Priority - urgent|Time|false|false||urgentnull|Urgent|Modifier|false|false||urgentnull|urgent - premium|LabModifier|false|false||urgentnull|null|Procedure|false|false||revascularizationnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Completely - dosing instruction fragment|Finding|false|false||completelynull|Complete|Modifier|false|false||completelynull|Occluded|Finding|false|false||occluded
null|Obstruction|Finding|false|false||occludednull|Burning Mouth Syndrome|Disorder|false|false||BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|Timing, LOINC Axis 3|Finding|false|false||timingnull|Timing|Time|false|false||timingnull|Scalable Vector Graphics|Entity|false|false||SVGnull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|year|Time|false|false||yearsnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Leukocyte adhesion deficiency type 1|Disorder|false|false||LAD
null|Leukocyte adhesion deficiency|Disorder|false|false||LADnull|ITGB2 wt Allele|Finding|false|false||LAD
null|DLD gene|Finding|false|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|false|false||LADnull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|ACSS2 protein, human|Drug|false|false||ACS
null|ACSS2 protein, human|Drug|false|false||ACSnull|Acrocallosal Syndrome|Disorder|false|false||ACS
null|Acute Chest Syndrome|Disorder|false|false||ACSnull|ACS - Activity Card Sort|Finding|false|false||ACS
null|American Community Survey|Finding|false|false||ACS
null|ACCS gene|Finding|false|false||ACS
null|CO-methylating acetyl-CoA synthase activity|Finding|false|false||ACS
null|PLA2G15 gene|Finding|false|false||ACS
null|ACSS2 wt Allele|Finding|false|false||ACS
null|ACSS2 gene|Finding|false|false||ACS
null|acetate-CoA ligase activity|Finding|false|false||ACSnull|anterior calcarine sulcus (human only)|Anatomy|false|false||ACSnull|Alternate Care Site|Device|false|false||ACSnull|American College of Surgeons|Entity|false|false||ACS
null|American Cancer Society|Entity|false|false||ACS
null|Alternate Care Site|Entity|false|false||ACSnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|eptifibatide|Drug|false|false||eptifibatide
null|eptifibatide|Drug|false|false||eptifibatidenull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||hrsnull|HARS1 wt Allele|Finding|false|false||hrs
null|HARS1 gene|Finding|false|false||hrs
null|HGS wt Allele|Finding|false|false||hrs
null|HGS gene|Finding|false|false||hrs
null|ATN1 wt Allele|Finding|false|false||hrs
null|SRSF5 gene|Finding|false|false||hrsnull|Hour|Time|false|false||hrsnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|captopril|Drug|false|false||captopril
null|captopril|Drug|false|false||captoprilnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Cardiac enzymes|Drug|false|false||Cardiac enzymes
null|Cardiac enzymes|Drug|false|false||Cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||Cardiac enzymesnull|null|Attribute|false|false||Cardiac enzymesnull|Cardiac attachment|Finding|false|false||Cardiacnull|Heart|Anatomy|false|false||Cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||Cardiacnull|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Peak level|Modifier|false|false||peaknull|Creatine Kinase MB Isoenzyme|Drug|false|false||CKMB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CKMBnull|Concern|Finding|false|false||concernnull|Acute heart failure|Disorder|false|false||acute heart failurenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Ischemic|Finding|false|false||ischemicnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|Radiolucent Lines|Finding|true|false||RLLnull|Structure of right lower lobe of lung|Anatomy|true|false||RLLnull|Pneumonia|Disorder|true|false||pneumonianull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|true|false||significantnull|Pulmonary Edema|Finding|true|false||pulmonary edemanull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|true|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|true|false||pulmonarynull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false||left ventricular systolic dysfunctionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|inferiority|Finding|false|false||inferiornull|Inferior|Modifier|false|false||inferiornull|Inferolateral|Modifier|false|false||inferolateralnull|Hypokinesia|Finding|false|false||hypokinesisnull|Initially|Time|false|false||Initiallynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Cardiac ventricular thrombosis|Disorder|false|false||ventricular thrombusnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Thrombus|Finding|false|false||thrombus
null|Blood Clot|Finding|false|false||thrombusnull|Thrombus <Thrombidae>|Entity|false|false||thrombusnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Bleeding risk|Finding|false|false||risk of bleedingnull|Risk|Finding|false|false||risk ofnull|Risk|Finding|false|false||risknull|Hemorrhage|Finding|false|false||bleedingnull|Benefit|LabModifier|false|false||benefitnull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|Hospitalization|Procedure|false|false||hospitalizationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Saturated|Phenomenon|false|false||saturationsnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Plain chest X-ray|Procedure|false|false||CXRnull|Radiolucent Lines|Finding|false|false||RLLnull|Structure of right lower lobe of lung|Anatomy|false|false||RLLnull|Pneumonia|Disorder|false|false||pneumonianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|metronidazole|Drug|false|false||metronidazole
null|metronidazole|Drug|false|false||metronidazolenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Radiolucent Lines|Finding|false|false||RLLnull|Structure of right lower lobe of lung|Anatomy|false|false||RLLnull|Pneumonia|Disorder|false|false||pneumonianull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Structure of right lower lobe of lung|Anatomy|false|false||right lower lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Extensive|Modifier|false|false||extensivenull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Diffuse|Modifier|false|false||diffusenull|null|Finding|false|false||lung nodulesnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Abnormality detected in sputum by cytology|Lab|false|false||sputum cytology positivenull|Sputum cytology (finding)|Finding|false|false||sputum cytologynull|Sputum Cytology Screening|Procedure|false|false||sputum cytologynull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Cytology--Technique|Procedure|false|false||cytology
null|Cytological Techniques|Procedure|false|false||cytologynull|Cytology|Title|false|false||cytologynull|cellular aspects|Modifier|false|false||cytologynull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|Initially|Time|false|false||initiallynull|combination - answer to question|Finding|false|false||combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Postobstructive pneumonia|Disorder|false|false||postobstructive pneumonianull|Pneumonia|Disorder|false|false||pneumonianull|Tumor Burden|Procedure|false|false||tumor burdennull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Burden|Finding|false|false||burdennull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Flagyl|Drug|false|false||flagyl
null|Flagyl|Drug|false|false||flagylnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Little's Disease|Disorder|false|false||littlenull|Only a Little|Finding|false|false||littlenull|Smallest|LabModifier|false|false||little
null|Small|LabModifier|false|false||littlenull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Improvement|Finding|false|false||improvementnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|Respiratory Status|Finding|false|false||Respiratory statusnull|null|Attribute|false|false||Respiratory statusnull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Flow|Phenomenon|false|false||flownull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Requirement|Finding|false|false||requirementnull|Oxygen nasal cannula|Device|false|false||nasal cannula
null|Nasal Cannula|Device|false|false||nasal cannulanull|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal brand of oxymetazoline|Drug|false|false||nasal
null|Nasal dosage form|Drug|false|false||nasalnull|Nasal Route of Administration|Finding|false|false||nasal
null|Nasal (intended site)|Finding|false|false||nasalnull|null|Anatomy|false|false||nasalnull|Specimen Type - Cannula|Finding|false|false||cannula
null|null|Finding|false|false||cannulanull|Body Parts - Cannula|Anatomy|false|false||cannulanull|Cannula device|Device|false|false||cannulanull|Calamus <grasshoppers>|Entity|false|false||cannulanull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Saturated|Phenomenon|false|false||saturationnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|masked - No information|Finding|false|false||mask
null|ANKHD1 gene|Finding|false|false||mask
null|STK26 gene|Finding|false|false||masknull|Protective Face Mask|Device|false|false||mask
null|Masks|Device|false|false||masknull|Helping Behavior|Finding|false|false||assistnull|Assisting (procedure)|Procedure|false|false||assistnull|American Stop Smoking Intervention for Cancer Prevention|Entity|false|false||assistnull|Assisted (qualifier value)|Modifier|false|false||assistnull|Alveolar ventilation function|Finding|false|false||oxygenation
null|Cell Respiration|Finding|false|false||oxygenationnull|null|Finding|false|false||Lung nodulesnull|Lung diseases|Disorder|false|false||Lungnull|Lung Problem|Finding|false|false||Lungnull|Chest>Lung|Anatomy|false|false||Lung
null|Lung|Anatomy|false|false||Lungnull|Carcinoma|Disorder|false|false||carcinomanull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Diffuse|Modifier|false|false||diffusenull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Abnormality detected in sputum by cytology|Lab|false|false||sputum cytology positivenull|Sputum cytology (finding)|Finding|false|false||sputum cytologynull|Sputum Cytology Screening|Procedure|false|false||sputum cytologynull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Cytology--Technique|Procedure|false|false||cytology
null|Cytological Techniques|Procedure|false|false||cytologynull|Cytology|Title|false|false||cytologynull|cellular aspects|Modifier|false|false||cytologynull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|THYROID DIAGNOSTIC RADIOPHARMACEUTICALS|Drug|false|false||thyroid
null|THYROID|Drug|false|false||thyroid
null|THYROID|Drug|false|false||thyroid
null|thyroid (USP)|Drug|false|false||thyroid
null|thyroid (USP)|Drug|false|false||thyroid
null|thyroid (USP)|Drug|false|false||thyroidnull|Thyroid Diseases|Disorder|false|false||thyroidnull|examination of thyroid|Procedure|false|false||thyroidnull|Thyroid Gland|Anatomy|false|false||thyroidnull|null|Time|false|false||priornull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Carcinoma|Disorder|false|false||carcinomanull|Extended Priority Codes - Routine|Finding|true|false||routine
null|Report priority - Routine|Finding|true|false||routine
null|Admission Type - Routine|Finding|true|false||routine
null|Level of Care - Routine|Finding|true|false||routine
null|Processing priority - Routine|Finding|true|false||routine
null|Referral priority - Routine|Finding|true|false||routinenull|Routine coag|Procedure|true|false||routinenull|Priority - Routine|Time|true|false||routinenull|Routine|Modifier|true|false||routinenull|Screening for cancer|Procedure|true|false||cancer screeningnull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|true|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Screening - procedure intent|Finding|true|false||screening
null|Special screening finding|Finding|true|false||screening
null|Aspects of disease screening|Finding|true|false||screeningnull|Screening for cancer|Procedure|true|false||screening
null|Disease Screening|Procedure|true|false||screening
null|research subject screening|Procedure|true|false||screening
null|Screening|Procedure|true|false||screening
null|Screening procedure|Procedure|true|false||screeningnull|Tissue diagnosis|Finding|true|false||tissue diagnosisnull|Tissue Specimen Code|Finding|true|false||tissuenull|Body tissue|Anatomy|true|false||tissuenull|Diagnosis Classification - Diagnosis|Finding|true|false||diagnosis
null|diagnosis aspects|Finding|true|false||diagnosisnull|Diagnosis|Procedure|true|false||diagnosisnull|null|Attribute|true|false||diagnosisnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Message Waiting Priority - High|Finding|true|false||high
null|high - ActExposureLevelCode|Finding|true|false||high
null|IPSS Risk Category High|Finding|true|false||high
null|IPSS-R Risk Category High|Finding|true|false||high
null|High (finding)|Finding|true|false||highnull|Observation Value - High|Modifier|true|false||high
null|High|Modifier|true|false||high
null|Abnormally high|Modifier|true|false||highnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Arylsulfatase A, human|Drug|false|false||asa
null|Arylsulfatase A, human|Drug|false|false||asa
null|aspirin|Drug|false|false||asa
null|aspirin|Drug|false|false||asanull|ARSA gene|Finding|false|false||asanull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Recent|Time|false|false||recentnull|Clinical act of insertion|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|null|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Imaging problem|Finding|true|false||imagingnull|Diagnostic Imaging|Procedure|true|false||imaging
null|Imaging Techniques|Procedure|true|false||imagingnull|Imaging Technology|Title|true|false||imagingnull|Problems with head|Disorder|true|false||headnull|Procedure on head|Procedure|true|false||headnull|Structure of head of caudate nucleus|Anatomy|true|false||head
null|Head|Anatomy|true|false||headnull|Head Device|Device|true|false||headnull|With staging|Finding|true|false||stagingnull|Venezuelan equine encephalitis virus subtype IIIA|Disorder|false|false||IIIanull|Multiple Pulmonary Nodules|Finding|true|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|true|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|true|false||pulmonarynull|Lung diseases|Disorder|true|false||lungnull|Lung Problem|Finding|true|false||lungnull|Chest>Lung|Anatomy|true|false||lung
null|Lung|Anatomy|true|false||lungnull|Obvious|Modifier|true|false||obviousnull|Distal Resection Margin|Attribute|true|false||distalnull|Distal (qualifier value)|Modifier|true|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|true|false||LADnull|Ladino Language|Entity|true|false||LADnull|Neoplasm Metastasis|Disorder|true|false||metastasis
null|Metastatic malignant neoplasm|Disorder|true|false||metastasisnull|Metastasis|Finding|true|false||metastasis
null|Metastatic Lesion|Finding|true|false||metastasisnull|Empiric|Modifier|false|false||Empiricnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Agent|Drug|false|false||agent
null|Pharmacologic Substance|Drug|false|false||agentnull|GDC Therapeutic Agent Terminology|Finding|false|false||agent
null|agent - RoleClass|Finding|false|false||agent
null|Protocol Agent|Finding|false|false||agentnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|pemetrexed|Drug|false|false||Pemetrexed
null|pemetrexed|Drug|false|false||Pemetrexednull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|dexamethasone|Drug|false|false||dexamethasone
null|dexamethasone|Drug|false|false||dexamethasonenull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Chronic Kidney Insufficiency|Disorder|false|false||Chronic renal insufficiencynull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Renal Insufficiency|Disorder|false|false||renal insufficiency
null|Kidney Failure|Disorder|false|false||renal insufficiencynull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Insufficiency|Finding|false|false||insufficiencynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|With glomerular filtration rate|Modifier|false|false||with GFRnull|RAPGEF5 gene|Finding|false|false||GFRnull|Glomerular Filtration Rate|LabModifier|false|false||GFRnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Renal function|Finding|false|false||renal functionnull|Kidney Function Tests|Procedure|false|false||renal functionnull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Mucomyst|Drug|false|false||mucomyst
null|Mucomyst|Drug|false|false||mucomystnull|null|Time|false|false||priornull|IV contrast|Drug|false|false||IV contrastnull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hyperkalemia|Finding|false|false||Hyperkalemia
null|Serum potassium level above reference range|Finding|false|false||Hyperkalemianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Transaction counts and value totals - day|Finding|true|false||day
null|Precision - day|Finding|true|false||daynull|Land Dayak Languages|Entity|true|false||daynull|day|Time|true|false||day
null|Daily|Time|true|false||daynull|null|Time|true|false||prior tonull|null|Time|true|false||priornull|Body Substance Discharge|Finding|true|false||discharge
null|Discharge Body Fluid|Finding|true|false||discharge
null|Body Fluid Discharge|Finding|true|false||discharge
null|null|Finding|true|false||dischargenull|Patient Discharge|Procedure|true|false||dischargenull|Electrocardiogram image|Finding|true|false||EKG
null|Electrocardiogram|Finding|true|false||EKGnull|Electrocardiography|Procedure|true|false||EKGnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Kayexalate|Drug|false|false||kayexalate
null|Kayexalate|Drug|false|false||kayexalatenull|Electrolytes|Drug|false|false||Electrolytes
null|Electrolytes|Drug|false|false||Electrolytes
null|Electrolyte [EPC]|Drug|false|false||Electrolytesnull|Daily|Time|false|false||dailynull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hypertensive disease|Disorder|false|false||HTNnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||Dailynull|ezetimibe / simvastatin|Drug|false|false||Ezetimibe-Simvastatinnull|ezetimibe|Drug|false|false||Ezetimibe
null|ezetimibe|Drug|false|false||Ezetimibenull|simvastatin|Drug|false|false||Simvastatin
null|simvastatin|Drug|false|false||Simvastatinnull|Vytorin|Drug|false|false||Vytorin
null|Vytorin|Drug|false|false||Vytorinnull|Daily|Time|false|false||dailynull|nifedipine|Drug|false|false||Nifedipine
null|nifedipine|Drug|false|false||Nifedipinenull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|/hour|Time|false|false||/hournull|Hour|Time|false|false||hournull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Sublingual Route of Administration|Finding|true|false||sublingual
null|Sublingual (intended site)|Finding|true|false||sublingualnull|Sublingual location|Modifier|true|false||sublingualnull|CIAO3 gene|Finding|true|false||PRNnull|As required|Time|true|false||PRN
null|Pro Re Nata|Time|true|false||PRNnull|Recent|Time|true|false||recentlynull|null|Time|true|false||priornull|propranolol|Drug|false|false||Propranolol
null|propranolol|Drug|false|false||Propranololnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|ST segment elevation myocardial infarction|Disorder|false|false||ST elevation myocardial infarctionnull|ST segment elevation (finding)|Finding|false|false||ST elevationnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Myocardial Infarction|Disorder|false|false||myocardial infarctionnull|null|Attribute|false|false||myocardial infarctionnull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false||infarctionnull|Carcinoma|Disorder|false|false||carcinomanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Requirement|Finding|false|false||requirementnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Chest pressure|Finding|false|false||chest pressurenull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Present|Finding|false|false||foundnull|Myocardial Infarction|Disorder|false|false||heart attacknull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Attack (finding)|Finding|false|false||attack
null|Attack behavior|Finding|false|false||attacknull|Attack device|Device|false|false||attacknull|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Disorder|false|false||cardiac catheterizationnull|Diagnostic Service Section ID - Cardiac Catheterization|Finding|false|false||cardiac catheterizationnull|Consent Type - Cardiac Catheterization|Procedure|false|false||cardiac catheterization
null|Cardiac Catheterization Procedures|Procedure|false|false||cardiac catheterizationnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Catheterization|Procedure|false|false||catheterizationnull|Bare metal stent|Device|false|false||bare metal stentnull|null|Modifier|false|false||barenull|Metal stent|Device|false|false||metal stentnull|Metals|Drug|false|false||metalnull|null|Device|false|false||stentnull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Lung|Anatomy|false|false||lungsnull|Sputum specimen|Finding|false|false||sputum samplenull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Specimen|Drug|false|false||samplenull|Nucleotide Sequence Sample Name|Finding|false|false||sample
null|Biospecimen|Finding|false|false||samplenull|Tumor cells, malignant|Anatomy|false|false||malignant cellsnull|Malignant (qualifier value)|Modifier|false|false||malignantnull|Cells|Anatomy|false|false||cellsnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Further|Modifier|false|false||furthernull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Every morning|Time|false|false||every morningnull|Morning|Time|false|false||morningnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|1 Month|Time|false|false||1 monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Ensure (product)|Drug|true|false||ensurenull|Malignant neoplasm of heart|Disorder|true|false||heart
null|benign neoplasm of heart|Disorder|true|false||heartnull|HEART PROBLEM|Finding|true|false||heartnull|Chest>Heart|Anatomy|true|false||heart
null|Heart|Anatomy|true|false||heartnull|null|Device|true|false||stentnull|Obstruction|Finding|true|false||blocked
null|Blocking|Finding|true|false||blockednull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions