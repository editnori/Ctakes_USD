CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Low Back Pain|Finding|false|false||Low back painnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Back Pain with Radiation|Finding|false|false||back pain with radiationnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Radiation Ionizing Radiotherapy|Procedure|false|false||radiation
null|Radiotherapy Research|Procedure|false|false||radiation
null|Radiation therapy (procedure)|Procedure|false|false||radiationnull|Electromagnetic Radiation|Phenomenon|false|false||radiation
null|Radiation|Phenomenon|false|false||radiationnull|Unit of radiation dose|LabModifier|false|false||radiationnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Decompression - action (qualifier value)|Finding|false|false||DECOMPRESSIONnull|Decompression|Procedure|false|false||DECOMPRESSION
null|Decompressive incision|Procedure|false|false||DECOMPRESSIONnull|external decompression|Phenomenon|false|false||DECOMPRESSIONnull|Fused structure|Finding|false|false||FUSIONnull|Fusion procedure|Procedure|false|false||FUSIONnull|Duraplasty|Procedure|false|false||DURAPLASTYnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aortic Aneurysm, Abdominal|Disorder|false|false||aneurysm, abdominal aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Aorta|Anatomy|false|false||aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Pallister W syndrome|Disorder|false|false||syndrome wnull|Syndrome|Disorder|false|false||syndromenull|Numerous|LabModifier|false|false||multiplenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Event|Event|false|false||eventnull|Bilateral|Modifier|false|false||bilateralnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|BRCA1 gene mutation|Disorder|false|false||BRCA1 mutationnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||mutationnull|Mutation|Finding|false|false||mutationnull|Malignant neoplasm of breast|Disorder|false|false||breast cancer
null|Breast Carcinoma|Disorder|false|false||breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|right-sided low back pain|Finding|false|false||right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false||lower back painnull|Lower back (surface region)|Anatomy|false|false||lower back
null|Lower back structure|Anatomy|false|false||lower backnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Radicular pain|Finding|false|false||radicular painnull|Dermatomal|Modifier|false|false||radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in right leg|Finding|false|false||right leg painnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Recent|Time|false|false||recentnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Background|Finding|false|false||backgroundnull|month|Time|false|false||monthsnull|Pain in right leg|Finding|false|false||right leg painnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Evidence of (contextual qualifier)|Finding|false|false||evidence ofnull|Evidence|Finding|false|false||evidencenull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|true|false||DVTnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|right trochanteric bursitis|Disorder|false|false||right trochanteric bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Injection of steroid|Procedure|false|false||steroid injectionnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Right tibia|Anatomy|false|false||right tibianull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Tibia pain|Finding|false|false||tibia painnull|Bone structure of tibia|Anatomy|false|false||tibianull|Tibia <Rostellariidae>|Entity|false|false||tibianull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT A
null|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT Anull|Nephrolithiasis|Disorder|false|false||nephrolithiasisnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Swelling|Finding|false|false||bulgenull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Narrow|Modifier|false|false||narrowing ofnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Spinal Canal|Anatomy|false|false||spinal canalnull|Spinal|Modifier|false|false||spinalnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Tooth Crowding|Finding|false|false||crowding
null|Crowding|Finding|false|false||crowdingnull|Malignant neoplasm of cauda equina|Disorder|false|false||cauda equinanull|Cauda Equina|Anatomy|false|false||cauda equinanull|Glanders|Disorder|false|false||equinanull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false||Varicose veinsnull|Varicose|Modifier|false|false||Varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false||A1Cnull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|false|false||colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|polyps|Disorder|false|false||polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false||CMC
null|Capillary malformation (disorder)|Disorder|false|false||CMCnull|MCC protocol|Procedure|false|false||CMCnull|Circulating Melanoma Cell|Anatomy|false|false||CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false||joint arthroplastynull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false||arthroplasty
null|Arthroplasty|Procedure|false|false||arthroplasty
null|Reconstruction of joint|Procedure|false|false||arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false||rotator cuff repairnull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Excision|Procedure|false|false||excision
null|removal technique|Procedure|false|false||excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false||digitnull|Digit structure|Anatomy|false|false||digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false||pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false||pancreatic duct
null|Pancreatic duct|Anatomy|false|false||pancreatic ductnull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false||pancreaticnull|Duct (organ) structure|Anatomy|false|false||duct
null|canal [body parts]|Anatomy|false|false||ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false||explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Malignant neoplasm of brain|Disorder|false|false||BRAIN CANCER
null|Brain Neoplasms|Disorder|false|false||BRAIN CANCERnull|Brain Diseases|Disorder|false|false||BRAINnull|Head>Brain|Anatomy|false|false||BRAIN
null|Brain|Anatomy|false|false||BRAINnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Platinum-Group Metal|Drug|false|false||PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false||PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false||PGMnull|phosphoglycerate mutase activity|Finding|false|false||PGMnull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Aunt|Subject|false|false||Auntnull|ovarian neoplasm|Disorder|false|true||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|true||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|Malignant Neoplasms|Disorder|false|true||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|true||CANCERnull|Paternal aunt|Subject|false|false||paternal auntnull|Paternal Relative|Subject|false|false||paternalnull|Paternal (qualifier value)|Modifier|false|false||paternalnull|Aunt|Subject|false|false||auntnull|Endometrial Carcinoma|Disorder|false|false||ENDOMETRIAL CANCER
null|Malignant neoplasm of endometrium|Disorder|false|false||ENDOMETRIAL CANCERnull|Endometrial|Modifier|false|false||ENDOMETRIALnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|STAT5A protein, human|Drug|false|false||MGF
null|IGF1 protein, human|Drug|false|false||MGF
null|IGF1 protein, human|Drug|false|false||MGF
null|STAT5A protein, human|Drug|false|false||MGF
null|Kit Ligand, human|Drug|false|false||MGF
null|Kit Ligand, human|Drug|false|false||MGFnull|STAT5A wt Allele|Finding|false|false||MGF
null|KITLG gene|Finding|false|false||MGF
null|STAT5A gene|Finding|false|false||MGF
null|KITLG wt Allele|Finding|false|false||MGFnull|Malignant neoplasm of prostate|Disorder|false|false||PROSTATE CANCER
null|Prostate carcinoma|Disorder|false|false||PROSTATE CANCERnull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false||PROSTATE
null|Prostatic Diseases|Disorder|false|false||PROSTATE
null|Carcinoma in situ of prostate|Disorder|false|false||PROSTATE
null|Benign neoplasm of prostate|Disorder|false|false||PROSTATEnull|Structure of prostate (body structure)|Anatomy|false|false||PROSTATE
null|Prostate|Anatomy|false|false||PROSTATEnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Malignant neoplasm of kidney|Disorder|false|false||KIDNEY CANCER
null|Renal carcinoma|Disorder|false|false||KIDNEY CANCERnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||KIDNEY
null|Benign neoplasm of kidney|Disorder|false|false||KIDNEYnull|Kidney problem|Finding|false|false||KIDNEYnull|examination of kidney|Procedure|false|false||KIDNEY
null|Procedures on Kidney|Procedure|false|false||KIDNEYnull|Kidney|Anatomy|false|false||KIDNEY
null|Both kidneys|Anatomy|false|false||KIDNEYnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Kidney Failure|Disorder|false|false||RENAL FAILUREnull|Urologic Diseases|Disorder|false|false||RENALnull|Kidney|Anatomy|false|false||RENALnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Congestive|Modifier|false|false||CONGESTIVEnull|Malignant neoplasm of heart|Disorder|false|false||HEART
null|benign neoplasm of heart|Disorder|false|false||HEARTnull|HEART PROBLEM|Finding|false|false||HEARTnull|Chest>Heart|Anatomy|false|false||HEART
null|Heart|Anatomy|false|false||HEARTnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Diabetes Mellitus|Disorder|false|false||DIABETES MELLITUSnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||DIABETES
null|Diabetes|Disorder|false|false||DIABETES
null|Diabetes Mellitus|Disorder|false|false||DIABETESnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Sister - courtesy title|Finding|false|false||Sister
null|Relationship - Sister|Finding|false|false||Sisternull|Sister|Subject|false|false||Sisternull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|true||age
null|Glycation End Products, Advanced|Drug|false|true||agenull|null|Attribute|false|true||agenull|Age|Subject|false|false||agenull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Throat cancer|Disorder|false|false||THROAT CANCERnull|Throat Homeopathic Medication|Drug|false|false||THROATnull|Specimen Type - Throat|Finding|false|false||THROAT
null|null|Finding|false|false||THROATnull|Throat|Anatomy|false|false||THROAT
null|Anterior portion of neck|Anatomy|false|false||THROAT
null|Pharyngeal structure|Anatomy|false|false||THROATnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Sister - courtesy title|Finding|false|false||Sister
null|Relationship - Sister|Finding|false|false||Sisternull|Sister|Subject|false|false||Sisternull|BRCA1 gene mutation|Disorder|false|false||BRCA1 MUTATIONnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||MUTATIONnull|Mutation|Finding|false|false||MUTATIONnull|Malignant neoplasm of breast|Disorder|false|true||BREAST CANCER
null|Breast Carcinoma|Disorder|false|true||BREAST CANCERnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||BREASTnull|Breast problem|Finding|false|false||BREASTnull|Procedures on breast|Procedure|false|false||BREASTnull|Breast|Anatomy|false|false||BREASTnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Daughter|Subject|false|false||Daughternull|Abnormal cervical smear|Finding|false|true||ABNORMAL PAP SMEARnull|Observation Interpretation - Abnormal|Finding|false|false||ABNORMAL
null|Abnormal|Finding|false|false||ABNORMALnull|Pap smear|Procedure|false|false||PAP SMEAR
null|Papanicolaou Test|Procedure|false|false||PAP SMEARnull|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false||PAP
null|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false||PAP
null|ACPP protein, human|Drug|false|false||PAP
null|ACPP protein, human|Drug|false|false||PAPnull|null|Finding|false|false||PAP
null|PAPOLA wt Allele|Finding|false|false||PAP
null|PDAP1 gene|Finding|false|false||PAP
null|TUSC2 wt Allele|Finding|false|false||PAP
null|ASAP1 wt Allele|Finding|false|false||PAP
null|ACP3 wt Allele|Finding|false|false||PAP
null|Pulmonary artery pressure|Finding|false|false||PAP
null|TUSC2 gene|Finding|false|false||PAP
null|ASAP2 gene|Finding|false|false||PAP
null|ASAP1 gene|Finding|false|false||PAP
null|REG3A gene|Finding|false|false||PAP
null|PITUITARY ADENOMA PREDISPOSITION|Finding|false|false||PAP
null|PAPOLA gene|Finding|false|false||PAP
null|ACP3 gene|Finding|false|false||PAP
null|REG3A wt Allele|Finding|false|false||PAP
null|MRPS30 gene|Finding|false|false||PAPnull|pars anterior of the paramedian lobule|Anatomy|false|false||PAPnull|Papiamento language|Entity|false|false||PAPnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|SON gene|Finding|false|false||Sonnull|Son (person)|Subject|false|false||Sonnull|Songhay Languages|Entity|false|false||Sonnull|Substance Abuse Problems|Disorder|false|false||SUBSTANCE ABUSE
null|Harmful pattern of substance use|Disorder|false|false||SUBSTANCE ABUSEnull|Substance|Drug|false|false||SUBSTANCEnull|administrative information regarding test substance|Finding|false|false||SUBSTANCEnull|null|Attribute|false|false||SUBSTANCEnull|Substance (attribute)|Modifier|false|false||SUBSTANCEnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Heroin overdose|Disorder|false|false||heroin overdosenull|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroinnull|Poisoning by heroin|Disorder|false|false||heroinnull|Drug Overdose|Disorder|false|false||overdosenull|Event Qualification - Overdose|Finding|false|false||overdose
null|Overdose|Finding|false|false||overdosenull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Weepiness|Finding|false|false||Tearfulnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Spasm|Finding|false|false||spasmsnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Surgical incisions|Procedure|false|false||incisionsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Healed|Finding|false|false||healednull|Axilla|Anatomy|false|false||axillanull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Movement|Finding|false|false||movementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||Swelling
null|Edema|Finding|false|false||Swellingnull|Palpable|Modifier|false|false||Palpablenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Medullary sponge kidney|Disorder|false|false||MSK
null|Medullary sponge kidney|Disorder|false|false||MSKnull|SIK1 gene|Finding|false|false||MSKnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|SI joint|Anatomy|false|false||SI Jointnull|Joint tenderness|Finding|false|false||Joint tendernessnull|Joint problem|Finding|false|false||Jointnull|null|Anatomy|false|false||Joint
null|Joints|Anatomy|false|false||Joint
null|Articular system|Anatomy|false|false||Jointnull|Joint Device|Device|false|false||Jointnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Radicular pain|Finding|false|false||Radicular painnull|Dermatomal|Modifier|false|false||Radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Hip flexion|Finding|false|false||hip flexionnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Knee flexion|Finding|false|false||knee flexionnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Plantar (qualifier value)|Anatomy|false|false||plantar
null|Sole of Foot|Anatomy|false|false||plantarnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Tact|Drug|false|false||tact
null|Tact|Drug|false|false||tact
null|Tact|Drug|false|false||tact
null|bis(tetraheptylammonium)tetraiodocyclopentane tellurate(IV)|Drug|false|false||tactnull|Ortho-|Finding|false|false||Orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||Orthonull|Spine Problem|Finding|false|false||Spinenull|Neuron spine|Anatomy|false|false||Spine
null|Vertebral column|Anatomy|false|false||Spinenull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|Telling untruths|Finding|false|false||Lyingnull|Supine Position|Modifier|false|false||Lyingnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|null|Attribute|false|false||resp effortnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||respnull|Respiratory rate|Attribute|false|false||respnull|Exertion|Finding|false|false||effortnull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|LAT protein, human|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|L-Type Amino Acid Transporter|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|ORC3 protein, human|Drug|false|false||lat
null|LAT protein, human|Drug|false|false||latnull|LAT gene|Finding|false|false||lat
null|ORC3 wt Allele|Finding|false|false||lat
null|ORC3 gene|Finding|false|false||lat
null|SPNS1 gene|Finding|false|false||latnull|Latin Language|Entity|false|false||latnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Thumb structure|Anatomy|false|false||thumbnull|Middle|Modifier|false|false||midnull|Upper extremity>Finger|Anatomy|false|false||finger
null|Fingers|Anatomy|false|false||finger
null|Fingers not including thumb|Anatomy|false|false||fingernull|Multiple Epiphyseal Dysplasia|Disorder|false|false||mednull|Master of Education|Finding|false|false||med
null|COMP wt Allele|Finding|false|false||med
null|COL9A3 gene|Finding|false|false||med
null|SCN8A wt Allele|Finding|false|false||med
null|COL9A2 gene|Finding|false|false||med
null|COMP gene|Finding|false|false||med
null|SCN8A gene|Finding|false|false||mednull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Trunk of elephant|Anatomy|false|false||Trunk
null|Trunk structure|Anatomy|false|false||Trunk
null|dendritic shaft|Anatomy|false|false||Trunknull|Pelvis>Groin|Anatomy|false|false||Groin
null|Inguinal region|Anatomy|false|false||Groin
null|Inguinal part of abdomen|Anatomy|false|false||Groinnull|Examination of knee joint|Procedure|false|false||Kneenull|Knee region structure|Anatomy|false|false||Knee
null|Knee|Anatomy|false|false||Knee
null|Lower extremity>Knee|Anatomy|false|false||Knee
null|Knee joint|Anatomy|false|false||Kneenull|Multiple Epiphyseal Dysplasia|Disorder|false|false||Mednull|Master of Education|Finding|false|false||Med
null|COMP wt Allele|Finding|false|false||Med
null|COL9A3 gene|Finding|false|false||Med
null|SCN8A wt Allele|Finding|false|false||Med
null|COL9A2 gene|Finding|false|false||Med
null|COMP gene|Finding|false|false||Med
null|SCN8A gene|Finding|false|false||Mednull|Structure of calf of leg|Anatomy|false|false||Calf
null|null|Anatomy|false|false||Calfnull|Cattle calf (organism)|Entity|false|false||Calfnull|Clava structure (body structure)|Anatomy|false|false||Grtnull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Toes|Anatomy|false|false||Toe
null|Toes|Anatomy|false|false||Toenull|Lower extremity>Thigh|Anatomy|false|false||Thigh
null|Thigh structure|Anatomy|false|false||Thighnull|motor movement|Finding|false|false||Motornull|Motor Device|Device|false|false||Motornull|CDAN1 wt Allele|Finding|false|false||Dlt
null|CDAN1 gene|Finding|false|false||Dltnull|imidazole mustard|Drug|false|false||Bic
null|imidazole mustard|Drug|false|false||Bicnull|MIR155HG gene|Finding|false|false||Bic
null|MIR155 gene|Finding|false|false||Bicnull|BIC Regimen|Procedure|false|false||Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false||Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false||Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Observation of reflex|Finding|false|false||Reflexes
null|Reflex action|Finding|false|false||Reflexesnull|Examination of reflexes|Procedure|false|false||Reflexesnull|imidazole mustard|Drug|false|false||Bic
null|imidazole mustard|Drug|false|false||Bicnull|MIR155HG gene|Finding|false|false||Bic
null|MIR155 gene|Finding|false|false||Bicnull|BIC Regimen|Procedure|false|false||Bicnull|Structure of inferior brachium of corpora quadrigemina|Anatomy|false|false||Bic
null|nucleus of the brachium of the inferior colliculus|Anatomy|false|false||Bicnull|TRI-AAT9-1 gene|Finding|false|false||Tri
null|Temptation and Restraint Inventory|Finding|false|false||Trinull|Fenamole|Drug|false|false||Pat
null|Fenamole|Drug|false|false||Patnull|Paroxysmal atrial tachycardia|Disorder|false|false||Patnull|glutamate-prephenate aminotransferase activity|Finding|false|false||Pat
null|aspartate-prephenate aminotransferase activity|Finding|false|false||Pat
null|protein acetyltransferase activity|Finding|false|false||Patnull|Thermoacoustic Computed Tomography|Procedure|false|false||Patnull|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Ach
null|acetylcholine|Drug|false|false||Achnull|Achondroplasia|Disorder|false|false||Achnull|FGFR3 wt Allele|Finding|false|false||Ach
null|FGFR3 gene|Finding|false|false||Ach
null|Ache|Finding|false|false||Achnull|Acoli Language|Entity|false|false||Achnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Babinski Reflex|Finding|false|false||Babinskinull|Clonus|Finding|false|false||Clonusnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|null|Attribute|false|false||MR THORACIC SPINEnull|Thoracic spine structure|Anatomy|false|false||THORACIC SPINEnull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false||THORACICnull|Chest|Anatomy|false|false||THORACICnull|Spine Problem|Finding|false|false||SPINEnull|Neuron spine|Anatomy|false|false||SPINE
null|Vertebral column|Anatomy|false|false||SPINEnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Spine Problem|Finding|false|false||SPINEnull|Neuron spine|Anatomy|false|false||SPINE
null|Vertebral column|Anatomy|false|false||SPINEnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|Central cord canal structure|Anatomy|false|false||central canalnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Level 5|Modifier|false|false||5 levelnull|Abnormal degeneration|Finding|false|false||degenerative changesnull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|LARGE1 wt Allele|Finding|false|false||Large
null|LARGE1 gene|Finding|false|false||Largenull|Large|LabModifier|false|false||Largenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Paramedian approach|Modifier|false|false||paramediannull|Upper|Modifier|false|false||superiornull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Extrusion|Finding|false|false||extrusionnull|Level 5|Modifier|false|false||5 levelnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lateral|Modifier|false|false||lateralnull|Mass Effect|Finding|false|false||mass effectnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Nerve|Anatomy|false|false||nervesnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Advanced phase|Modifier|false|false||Advancednull|Abnormal degeneration|Finding|false|false||degenerative changesnull|biologic degeneration|Finding|false|false||degenerative
null|Abnormal degeneration|Finding|false|false||degenerativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Lumbar spine structure|Anatomy|false|false||lumbar spine
null|Bone structure of lumbar vertebra|Anatomy|false|false||lumbar spinenull|Lumbar Region|Anatomy|false|false||lumbarnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Central cord canal structure|Anatomy|false|false||central canalnull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Moderate to severe|Modifier|false|false||moderate to severenull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Levels (qualifier value)|Modifier|false|false||levelsnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Lumbar spine structure|Anatomy|false|false||lumbar spine
null|Bone structure of lumbar vertebra|Anatomy|false|false||lumbar spinenull|Lumbar Region|Anatomy|false|false||lumbarnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Abnormal degeneration|Finding|false|false||Degenerative changesnull|biologic degeneration|Finding|false|false||Degenerative
null|Abnormal degeneration|Finding|false|false||Degenerativenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Thoracic spine structure|Anatomy|false|false||thoracic spinenull|Dissecting Thoracic Aortic Aneurysm|Disorder|false|false||thoracicnull|Chest|Anatomy|false|false||thoracicnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Mild to moderate|Modifier|false|false||mild-to-moderatenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Moderate - Severity of Illness Code|Finding|false|false||moderate
null|Moderate|Finding|false|false||moderatenull|Moderate (severity modifier)|Modifier|false|false||moderate
null|Moderate - Allergy Severity|Modifier|false|false||moderate
null|Moderation|Modifier|false|false||moderatenull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Foraminal|Modifier|false|false||foraminalnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|null|Attribute|false|false||CT ABDnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Malignant neoplasm of pelvis|Disorder|false|false||PELVISnull|Pelvis problem|Finding|false|false||PELVISnull|Pelvis+|Anatomy|false|false||PELVIS
null|Pelvic cavity structure|Anatomy|false|false||PELVIS
null|Pelvis|Anatomy|false|false||PELVISnull|Contrast Media|Drug|false|false||CONTRASTnull|Contrast|Modifier|false|false||CONTRASTnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Malignant neoplasm of abdomen|Disorder|true|false||abdomennull|Abdomen problem|Finding|true|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|true|false||pelvisnull|Pelvis problem|Finding|true|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Obstructed|Finding|true|false||obstructivenull|Nephrolithiasis|Disorder|false|false||renal stonenull|Renal stone (substance)|Finding|false|false||renal stone
null|Kidney Calculi|Finding|false|false||renal stonenull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Calculi|Finding|false|false||stonenull|Pyelonephritis|Disorder|false|false||pyelonephritisnull|Diverticulosis of sigmoid colon|Disorder|false|false||Sigmoid diverticulosisnull|Sigmoid colon|Anatomy|false|false||Sigmoidnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Diverticulitis|Disorder|false|false||diverticulitisnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||Labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Low Back Pain|Finding|false|false||Low Back painnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Back Pain|Finding|false|false||Back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in lower limb|Finding|false|false||Leg Painnull|Leg|Anatomy|false|false||Leg
null|Lower Extremity|Anatomy|false|false||Legnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Radiculopathy|Disorder|false|false||Radiculopathynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|right-sided low back pain|Finding|false|false||right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false||lower back painnull|Lower back (surface region)|Anatomy|false|false||lower back
null|Lower back structure|Anatomy|false|false||lower backnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Prominent|Modifier|false|false||prominentnull|Protein Component|Drug|false|false||component
null|Protein Component|Drug|false|false||componentnull|Specimen Child Role - Component|Finding|false|false||component
null|Component (part)|Finding|false|false||component
null|Component, LOINC Axis 1|Finding|false|false||componentnull|Component object|Device|false|false||componentnull|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT A
null|Choline-Phosphate Cytidylyltransferase A|Drug|false|false||CT Anull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Visceral|Modifier|false|false||visceralnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Nephrolithiasis|Disorder|false|false||nephrolithiasisnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Lumbar spine structure|Anatomy|false|false||L spinenull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Swelling|Finding|false|false||bulgenull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Narrow|Modifier|false|false||narrowing ofnull|Narrowing|Disorder|false|false||narrowingnull|Narrowed structure|Modifier|false|false||narrowing
null|Narrow|Modifier|false|false||narrowingnull|Spinal|Modifier|false|false||spinalnull|canal [body parts]|Anatomy|false|false||canal
null|Pulp Canals|Anatomy|false|false||canalnull|Geographic canal|Entity|false|false||canalnull|Extrusion|Finding|false|false||extrusionnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Fourth lumbar nerve|Anatomy|false|false||L4 nervenull|Nerve root structure|Anatomy|false|false||nerve rootnull|Nerve|Anatomy|false|false||nervenull|Tree Root (hierarchy)|Finding|false|false||rootnull|Tooth root structure|Anatomy|false|false||root
null|Root body part|Anatomy|false|false||rootnull|Plant Roots|Entity|false|false||rootnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Recent|Time|false|false||recentlynull|Pain in right leg|Finding|false|false||right leg painnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Bursitis|Disorder|false|false||bursitisnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Corticosteroid [EPC]|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroid
null|Adrenal Cortex Hormones|Drug|false|false||corticosteroidnull|Current (present time)|Time|false|false||Currentlynull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Compression of umbilical cord|Disorder|true|false||cord compression
null|Compression of spinal cord|Disorder|true|false||cord compressionnull|Cone-Rod Dystrophy 2|Disorder|false|false||cordnull|Cord - Body Parts|Anatomy|false|false||cordnull|Cord Device|Device|false|false||cordnull|null|Finding|true|false||compression
null|Compressed structure|Finding|true|false||compressionnull|Compression Therapy|Procedure|true|false||compression
null|Data Compression|Procedure|true|false||compressionnull|Compression|Phenomenon|true|false||compressionnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Ortho-|Finding|false|false||orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||orthonull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|Decompression - action (qualifier value)|Finding|false|false||DECOMPRESSIONnull|Decompression|Procedure|false|false||DECOMPRESSION
null|Decompressive incision|Procedure|false|false||DECOMPRESSIONnull|external decompression|Phenomenon|false|false||DECOMPRESSIONnull|Fused structure|Finding|false|false||FUSIONnull|Fusion procedure|Procedure|false|false||FUSIONnull|Duraplasty|Procedure|false|false||DURAPLASTYnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Dysuria|Finding|false|false||Dysurianull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Recent|Time|false|false||recentlynull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Specimen Type - Leukocytes|Finding|false|false||leukocytes
null|null|Finding|false|false||leukocytesnull|Leukocytes|Anatomy|false|false||leukocytesnull|Leukocytes|Anatomy|false|false||WBCnull|Urine culture|Procedure|false|false||urine culturenull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Bacterial|Modifier|false|false||bacterialnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Contamination|Finding|false|false||contaminationnull|adulteration|Phenomenon|false|false||contaminationnull|Specimen Reject Reason - Contamination|Modifier|false|false||contaminationnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Abdominal Pain|Finding|false|false||Abdominal painnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constipation|Finding|false|false||constipationnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|opioid use|Disorder|false|false||opioid usenull|Opioids|Drug|false|false||opioid
null|Opioids|Drug|false|false||opioid
null|Opioids|Drug|false|false||opioidnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Report (document)|Finding|false|false||Reportsnull|Reporting|Procedure|false|false||Reportsnull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Bactrim DS|Drug|false|false||bactrim DS
null|Bactrim DS|Drug|false|false||bactrim DSnull|Bactrim|Drug|false|false||bactrim
null|Bactrim|Drug|false|false||bactrimnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|Lupus anticoagulant positive|Lab|false|false||Lupus anticoagulant positivenull|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulant
null|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulantnull|Lupus anticoagulant disorder|Disorder|false|false||Lupus anticoagulantnull|null|Finding|false|false||Lupus anticoagulantnull|Lupus anticoagulant assay|Procedure|false|false||Lupus anticoagulantnull|Chronic discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus|Disorder|false|false||Lupus
null|Lupus Vulgaris|Disorder|false|false||Lupus
null|Discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus, Systemic|Disorder|false|false||Lupusnull|Anti-coagulant [EPC]|Drug|false|false||anticoagulant
null|Anticoagulants|Drug|false|false||anticoagulantnull|Bilateral|Modifier|false|false||bilateralnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|day|Time|false|false||daysnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin, porcine|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparin
null|heparin|Drug|false|false||heparinnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Charts (publication)|Finding|false|false||chartnull|chart [medical device]|Device|false|false||chartnull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|null|Attribute|false|false||CT abdnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||abdnull|ABD (body structure)|Anatomy|false|false||abd
null|Abdomen|Anatomy|false|false||abdnull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Aortic Aneurysm, Abdominal|Disorder|false|false||abdominal aortic aneurysmnull|null|Attribute|false|false||abdominal aortic aneurysmnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|null|Disorder|false|false||aortic aneurysm
null|Aortic Aneurysm|Disorder|false|false||aortic aneurysmnull|Aorta|Anatomy|false|false||aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Vitamin D Deficiency|Disorder|false|false||Vitamin D deficiencynull|Decreased circulating vitamin D concentration|Finding|false|false||Vitamin D deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Daily|Time|false|false||dailynull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPAPnull|Continuous Positive Airway Pressure|Procedure|false|false||CPAPnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||Medsnull|Medications|Finding|false|false||Medsnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|Daily|Time|false|false||dailynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|Opioids|Drug|false|false||opioids
null|Opioids|Drug|false|false||opioids
null|Opioids|Drug|false|false||opioids
null|Analgesics, Opioid|Drug|false|false||opioids
null|Analgesics, Opioid|Drug|false|false||opioidsnull|ARID1A protein, human|Drug|false|false||Held
null|ARID1A protein, human|Drug|false|false||Heldnull|Held - activity status|Finding|false|false||Held
null|ARID1A wt Allele|Finding|false|false||Heldnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Daily|Time|false|false||dailynull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Rare|Modifier|false|false||rarelynull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Ortho-|Finding|false|false||Orthonull|Ortho Pharmaceutical Ltd|Entity|false|false||Orthonull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aortic Aneurysm, Abdominal|Disorder|false|false||aneurysm, abdominal aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Aorta|Anatomy|false|false||aorticnull|Aneurysm|Finding|false|false||aneurysmnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Pallister W syndrome|Disorder|false|false||syndrome wnull|Syndrome|Disorder|false|false||syndromenull|Numerous|LabModifier|false|false||multiplenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Event|Event|false|false||eventnull|Bilateral|Modifier|false|false||bilateralnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|BRCA1 gene mutation|Disorder|false|false||BRCA1 mutationnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||mutationnull|Mutation|Finding|false|false||mutationnull|Malignant neoplasm of breast|Disorder|false|false||breast cancer
null|Breast Carcinoma|Disorder|false|false||breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|right-sided low back pain|Finding|false|false||right lower back painnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Low Back Pain|Finding|false|false||lower back painnull|Lower back (surface region)|Anatomy|false|false||lower back
null|Lower back structure|Anatomy|false|false||lower backnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Radicular pain|Finding|false|false||radicular painnull|Dermatomal|Modifier|false|false||radicularnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pain in right leg|Finding|false|false||right leg painnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Intervertebral Disk Displacement|Disorder|false|false||disc herniationsnull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Hernia|Disorder|false|false||herniationsnull|Diskectomy|Procedure|false|false||discectomynull|Fused structure|Finding|false|false||fusionnull|Fusion procedure|Procedure|false|false||fusionnull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Course|Time|false|false||coursenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Procedure on spinal cord (procedure)|Procedure|false|false||Spine Surgery
null|Operation on spinal cord (procedure)|Procedure|false|false||Spine Surgerynull|Spine Problem|Finding|false|false||Spinenull|Neuron spine|Anatomy|false|false||Spine
null|Vertebral column|Anatomy|false|false||Spinenull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Operating Room|Device|false|false||Operating Roomnull|Operating Room|Entity|false|false||Operating Roomnull|Patient location type - Operating Room|Modifier|false|false||Operating Roomnull|Operating|Finding|false|false||Operatingnull|Room - Patient location type|Modifier|false|false||Room
null|Room|Modifier|false|false||Roomnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|null|Attribute|false|false||operative notenull|Operative|Time|false|false||operativenull|Further|Modifier|false|false||furthernull|Details|Modifier|false|false||detailsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Complication (attribute)|Finding|false|false||complication
null|Complication|Finding|false|false||complicationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Postoperative deep vein thrombosis|Disorder|false|false||Postoperative DVTnull|Postoperative Period|Time|false|false||Postoperativenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Coumadin|Drug|false|false||coumadin
null|Coumadin|Drug|false|false||coumadinnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Bed rest|Procedure|false|false||bedrestnull|Dural tear|Disorder|false|false||dural tearnull|Laceration|Disorder|false|false||tear
null|Rupture|Disorder|false|false||tearnull|Tears (substance)|Finding|false|false||tearnull|Tear Shape|Modifier|false|false||tearnull|Precaution|Finding|false|false||precautionsnull|Hour|Time|false|false||hoursnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|Intravenous Route of Administration|Finding|false|false||Intravenousnull|Intravenous|Modifier|false|false||Intravenousnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Postoperative Period|Time|false|false||postopnull|Type of Agreement - Standard|Finding|false|false||standard
null|Standard (document)|Finding|false|false||standardnull|Standard base excess calculation technique|Procedure|false|false||standardnull|Standard (qualifier)|Modifier|false|false||standardnull|Clinical trial protocol document|Finding|false|false||protocol
null|Study Protocol|Finding|false|false||protocol
null|Protocols documentation|Finding|false|false||protocol
null|Protocol - answer to question|Finding|false|false||protocol
null|Library Protocol|Finding|false|false||protocolnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Pain, Postoperative|Finding|false|false||postop painnull|Postoperative Period|Time|false|false||postopnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical therapynull|Physical therapy|Procedure|false|false||Physical therapynull|Physical therapy (field)|Title|false|false||Physical therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Diagnostic Service Section ID - Occupational Therapy|Finding|false|false||Occupational therapynull|Occupational therapy (procedure)|Procedure|false|false||Occupational therapynull|Occupational|Finding|false|false||Occupationalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|physical therapy mobilization (treatment)|Procedure|false|false||mobilization
null|Mobilization (procedure)|Procedure|false|false||mobilizationnull|Ambulate|Finding|false|false||ambulatenull|VISCERAL LEIOMYOPATHY, AFRICAN DEGENERATIVE|Disorder|false|false||ADLnull|Activity of daily living (function)|Finding|false|false||ADL
null|SGCA gene|Finding|false|false||ADL
null|SGCA wt Allele|Finding|false|false||ADLnull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Course|Time|false|false||coursenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||acute blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||acute blood loss anemianull|Acute hemorrhage|Finding|false|false||acute blood lossnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||blood loss anemia
null|Anemia due to blood loss|Disorder|false|false||blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||blood loss anemianull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Constipation|Finding|false|false||constipationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Hypokalemia|Finding|false|false||hypokalemianull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||Acute blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||Acute blood loss anemianull|Acute hemorrhage|Finding|false|false||Acute blood lossnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Iron deficiency anemia secondary to chronic blood loss|Disorder|false|false||blood loss anemia
null|Anemia due to blood loss|Disorder|false|false||blood loss anemia
null|Acute posthaemorrhagic anaemia|Disorder|false|false||blood loss anemianull|Blood Loss|Finding|false|false||blood loss
null|Hemorrhage|Finding|false|false||blood lossnull|Actual blood loss|LabModifier|false|false||blood lossnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Intervention regimes|Procedure|true|false||intervention
null|Nursing interventions|Procedure|true|false||intervention
null|Interventional procedure|Procedure|true|false||interventionnull|Immediate Release Dosage Form|Drug|false|false||Immediate releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Valium|Drug|false|false||Valium
null|Valium|Drug|false|false||Valiumnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Drug|false|false||Oral Potassiumnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Hypokalemia|Finding|false|false||hypokalemianull|Laboratory test finding|Lab|false|false||labsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Hospital course|Finding|false|false||Hospital coursenull|null|Attribute|false|false||Hospital coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||coursenull|null|Modifier|false|false||unremarkablenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Feeling comfortable|Finding|false|false||comfortablenull|Oral pain|Finding|false|false||oral painnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false||PTCH
null|PTCH1 wt Allele|Finding|false|false||PTCH
null|PTCH1 gene|Finding|false|false||PTCH
null|PTCH1 protein, human|Finding|false|false||PTCHnull|Every morning|Time|false|false||QAMnull|Right hip region structure|Anatomy|false|false||right hipnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false||Leg swellingnull|Leg|Anatomy|false|false||Leg
null|Lower Extremity|Anatomy|false|false||Legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|diazepam|Drug|false|false||Diazepam
null|diazepam|Drug|false|false||Diazepamnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Spasm|Finding|false|false||spasm
null|KANTR gene|Finding|false|false||spasmnull|Somnolence|Disorder|false|false||drowsinessnull|Drowsiness|Finding|false|false||drowsinessnull|diazepam|Drug|false|false||diazepam
null|diazepam|Drug|false|false||diazepamnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid Syndromenull|Syndrome|Disorder|false|false||Syndromenull|Biomaterial Treatment|Finding|false|false||Treatment
null|Treating|Finding|false|false||Treatment
null|therapeutic aspects|Finding|false|false||Treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||Treatment
null|Administration (procedure)|Procedure|false|false||Treatment
null|Therapeutic procedure|Procedure|false|false||Treatmentnull|Fixation of dental bridge|Procedure|false|false||Bridgenull|Type of bridge device|Device|false|false||Bridgenull|morphine sulfate|Drug|false|false||Morphine Sulfate
null|morphine sulfate|Drug|false|false||Morphine Sulfatenull|morphine|Drug|false|false||Morphine
null|morphine|Drug|false|false||Morphinenull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfate
null|Sulfates, Inorganic|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|sulfate ion|Drug|false|false||Sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||Sulfatenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Intrinsic drive|Finding|false|false||drivenull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false||Leg swellingnull|Leg|Anatomy|false|false||Leg
null|Lower Extremity|Anatomy|false|false||Legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false||PTCH
null|PTCH1 wt Allele|Finding|false|false||PTCH
null|PTCH1 gene|Finding|false|false||PTCH
null|PTCH1 protein, human|Finding|false|false||PTCHnull|Every morning|Time|false|false||QAMnull|Right hip region structure|Anatomy|false|false||right hipnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Spinal stenosis of lumbar region|Disorder|false|false||Lumbar spinal stenosisnull|Lumbar Region|Anatomy|false|false||Lumbarnull|Spinal canal stenosis|Disorder|false|false||spinal stenosis
null|Spinal Stenosis|Disorder|false|false||spinal stenosisnull|Spinal|Modifier|false|false||spinalnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Spondylolisthesis, L4-L5|Finding|false|false||Spondylolisthesis, L4-L5null|Congenital spondylolisthesis|Disorder|false|false||Spondylolisthesis
null|Spondylolisthesis|Disorder|false|false||Spondylolisthesis
null|Acquired spondylolisthesis|Disorder|false|false||Spondylolisthesisnull|urinastatin|Drug|false|false||UTI
null|urinastatin|Drug|false|false||UTInull|Urinary tract infection|Disorder|false|false||UTInull|AMBP wt Allele|Finding|false|false||UTI
null|AMBP gene|Finding|false|false||UTInull|Constipation|Finding|false|false||Constipationnull|Neoplasm Metastasis|Disorder|false|false||Secondarynull|metastatic qualifier|Finding|false|false||Secondarynull|Secondary to|Modifier|false|false||Secondarynull|second (number)|LabModifier|false|false||Secondarynull|Diagnosis|Procedure|false|false||Diagnosesnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPAPnull|Continuous Positive Airway Pressure|Procedure|false|false||CPAPnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Back Pain|Finding|false|false||back painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Structure of right lower leg|Anatomy|false|false||right leg
null|Right lower extremity|Anatomy|false|false||right legnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Difficult (qualifier value)|Finding|false|false||difficultnull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Intervertebral Disk Displacement|Disorder|false|false||disc herniationnull|Disk Drug Form|Drug|false|false||discnull|Disc (List bullets)|Finding|false|false||disc
null|Discontinued|Finding|false|false||discnull|Disc - Body Part|Anatomy|false|false||disc
null|death-inducing signaling complex location|Anatomy|false|false||discnull|Disk Device|Device|false|false||discnull|Disk Shape|Modifier|false|false||discnull|Disk Dosing Unit|LabModifier|false|false||discnull|Hernia|Disorder|false|false||herniationnull|Lower back (surface region)|Anatomy|false|false||lower back
null|Lower back structure|Anatomy|false|false||lower backnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Science of Etiology|Finding|false|false||cause
null|Etiology aspects|Finding|false|false||causenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Surgeon|Subject|false|false||surgeonsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constant - dosing instruction fragment|Finding|false|false||constantnull|Constant (qualifier)|Modifier|false|false||constantnull|Past 30 days|Time|false|false||past monthnull|Transaction counts and value totals - month|Finding|false|false||month
null|Precision - month|Finding|false|false||monthnull|month|Time|false|false||month
null|Monthly (qualifier value)|Time|false|false||monthnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|SAFE-Biopharma Standard|Finding|false|false||safenull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Decompression of spinal cord|Procedure|false|false||spinal decompression
null|Laminectomy|Procedure|false|false||spinal decompressionnull|Spinal|Modifier|false|false||spinalnull|Decompression - action (qualifier value)|Finding|false|false||decompressionnull|Decompression|Procedure|false|false||decompression
null|Decompressive incision|Procedure|false|false||decompressionnull|external decompression|Phenomenon|false|false||decompressionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Pain, Burning|Finding|false|false||burning painnull|Burning sensation|Finding|false|false||burningnull|Burning sensation quality|Modifier|false|false||burningnull|Dysuria|Finding|false|false||pain with urinationnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Urination|Finding|false|false||urinationnull|Urinary tract infection|Disorder|false|false||urinary tract infectionnull|Urinary tract|Anatomy|false|false||urinary tract
null|Urinary system|Anatomy|false|false||urinary tractnull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Tract|Anatomy|false|false||tractnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Lumbar Region|Anatomy|false|false||Lumbarnull|Decompression - action (qualifier value)|Finding|false|false||Decompressionnull|Decompression|Procedure|false|false||Decompression
null|Decompressive incision|Procedure|false|false||Decompressionnull|external decompression|Phenomenon|false|false||Decompressionnull|Fused structure|Finding|false|false||Fusionnull|Fusion procedure|Procedure|false|false||Fusionnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Lumbar Region|Anatomy|false|false||Lumbarnull|Decompression - action (qualifier value)|Finding|false|false||Decompressionnull|Decompression|Procedure|false|false||Decompression
null|Decompressive incision|Procedure|false|false||Decompressionnull|external decompression|Phenomenon|false|false||Decompressionnull|Fused structure|Finding|false|false||Fusionnull|Fusion procedure|Procedure|false|false||Fusionnull|Stat (do immediately)|Time|false|false||Immediatelynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|Greater|LabModifier|false|false||greaternull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|More|LabModifier|false|false||morenull|Feeling comfortable|Finding|false|false||comfortablenull|Does sit|Finding|true|false||sit
null|Sitting position|Finding|true|false||sit
null|HHAT gene|Finding|true|false||sit
null|SIT1 gene|Finding|true|false||sitnull|Does stand|Finding|true|false||stand
null|standards characteristics|Finding|true|false||standnull|Stand (physical object)|Device|true|false||stand
null|Stand Device|Device|true|false||standnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|45 Minutes|Time|false|false||45 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Encounter due to care involving use of rehabilitation procedures|Finding|false|false||Rehabilitation
null|Rehabilitation aspects|Finding|false|false||Rehabilitationnull|Rehabilitation therapy|Procedure|false|false||Rehabilitationnull|null|Title|false|false||Rehabilitationnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Walking (function)|Finding|false|false||walknull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|part of|Modifier|false|false||part ofnull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Much|Finding|false|false||muchnull|Terminology Kind|Finding|false|false||kindnull|null|Modifier|false|false||kindnull|Lifting|Event|false|false||liftingnull|Diet (animal life circumstance)|Drug|false|false||Diet
null|Diet|Drug|false|false||Dietnull|diet - supply|Finding|false|false||Dietnull|Diet therapy|Procedure|false|false||Dietnull|MCL1 wt Allele|Finding|false|false||Eat
null|Eating|Finding|false|false||Eatnull|Diet, Healthy|Finding|false|false||healthy dietnull|Healthy|Modifier|false|false||healthynull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Constipation|Finding|false|false||constipationnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Issue (document)|Finding|false|false||issue
null|Problem|Finding|false|false||issuenull|Issue (action)|Event|false|false||issuenull|Application of brace (procedure)|Procedure|false|false||Bracenull|Braces - Orthopedic appliances|Device|false|false||Brace
null|Braces - garment|Device|false|false||Bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|Application of brace (procedure)|Procedure|false|false||bracenull|Braces - Orthopedic appliances|Device|false|false||brace
null|Braces - garment|Device|false|false||bracenull|history of recreational walking|Finding|false|false||walking
null|walking - neurological symptom|Finding|false|false||walking
null|Walking (function)|Finding|false|false||walkingnull|Chairs|Device|false|false||chairnull|Chairperson|Subject|false|false||chairnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Wound care management|Procedure|false|false||Wound Care
null|wound care|Procedure|false|false||Wound Carenull|Wound Care kit|Device|false|false||Wound Carenull|Traumatic Wound|Disorder|false|false||Wound
null|Wounds and Injuries|Disorder|false|false||Wound
null|Traumatic injury|Disorder|false|false||Woundnull|Route of Administration - Wound|Finding|false|false||Wound
null|null|Finding|false|false||Wound
null|Specimen Type - Wound|Finding|false|false||Woundnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|null|Device|false|false||dry dressingnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Appointments|Event|false|false||appointmentnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Bathing|Procedure|false|false||bathnull|Pool (action)|Finding|false|false||poolnull|Sample pool|Attribute|false|false||poolnull|Pool (environment)|Entity|false|false||poolnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Moist|Modifier|false|false||wetnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Additional|Finding|false|false||Additionalnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|72 Hours|Time|false|false||72 hoursnull|Hour|Time|false|false||hoursnull|refill|Finding|false|false||refillnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Authorization Mode - Fax|Finding|false|false||fax
null|Fax Number|Finding|false|false||faxnull|Facsimile Machine|Device|false|false||fax
null|Telefacsimile|Device|false|false||faxnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Prescription (procedure)|Procedure|false|false||prescriptionsnull|null|Attribute|false|false||prescriptionsnull|Oxycontin|Drug|false|false||oxycontin
null|Oxycontin|Drug|false|false||oxycontinnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Percocet|Drug|false|false||percocet
null|Percocet|Drug|false|false||percocetnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|90 days|Time|false|false||90 daysnull|day|Time|false|false||daysnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Follow-up status|Finding|false|false||Follow upnull|follow-up|Procedure|false|false||Follow upnull|Follow - dosing instruction imperative|Finding|false|false||Follow
null|Follow|Finding|false|false||Follownull|Followed by|Time|false|false||Follownull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Appointments|Event|false|false||appointmentnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Visit|Finding|false|false||visitnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|X-rays, Homeopathic Preparations|Drug|false|false||X-raysnull|Plain x-ray|Procedure|false|false||X-rays
null|Diagnostic radiologic examination|Procedure|false|false||X-raysnull|Roentgen Rays|Phenomenon|false|false||X-raysnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|Full|Modifier|false|false||fullnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Academic degree|Finding|false|false||degreesnull|Degree or extent|LabModifier|false|false||degreesnull|Degrees fahrenheit|LabModifier|false|false||Fahrenheitnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|Weight-Bearing state|Subject|false|false||Weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|Bearing Device|Device|false|false||bearingnull|Gait|Finding|false|false||Gaitnull|Balance training|Procedure|false|false||balance trainingnull|Balance (substance)|Drug|false|false||balance
null|Balance (substance)|Drug|false|false||balancenull|Ability to balance|Finding|false|false||balance
null|Equilibrium|Finding|false|false||balancenull|examination of balance|Procedure|false|false||balancenull|balance device|Device|false|false||balancenull|Balanced (qualifier value)|Modifier|false|false||balancenull|Processing ID - Training|Finding|false|false||trainingnull|Training Programs|Procedure|false|false||training
null|Training|Procedure|false|false||trainingnull|training aspects|Modifier|false|false||trainingnull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|Significant|Finding|true|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Decompression Sickness|Disorder|true|false||bendingnull|Bending - Changing basic body position|Finding|true|false||bending
null|Does bend|Finding|true|false||bendingnull|Bent|Modifier|false|false||bendingnull|Musculoskeletal torsion (function)|Finding|true|false||twisting
null|Torsion (malposition)|Finding|true|false||twistingnull|Therapeutic procedure|Procedure|false|false||Treatmentsnull|Frequency|Finding|false|false||Frequency
null|How Often|Finding|false|false||Frequencynull|With frequency|Time|false|false||Frequency
null|Frequencies (time pattern)|Time|false|false||Frequencynull|Kind of quantity - Frequency|LabModifier|false|false||Frequency
null|Statistical Frequency|LabModifier|false|false||Frequency
null|Spatial Frequency|LabModifier|false|false||Frequencynull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|null|Device|false|false||dry dressingnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Bathing|Procedure|false|false||bathnull|Pool (action)|Finding|false|false||poolnull|Sample pool|Attribute|false|false||poolnull|Pool (environment)|Entity|false|false||poolnull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Surgical wound|Disorder|false|false||incisionnull|Surgical incisions|Procedure|false|false||incisionnull|Cranial incision point|Anatomy|false|false||incisionnull|Moist|Modifier|false|false||wetnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions