 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
Allergies|160,169
:|169,170
<EOL>|171,172
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
Chief|236,241
Complaint|242,251
:|251,252
<EOL>|252,253
DVT|253,256
<EOL>|256,257
<EOL>|258,259
Major|259,264
Surgical|265,273
or|274,276
Invasive|277,285
Procedure|286,295
:|295,296
<EOL>|296,297
EGD|297,300
<EOL>|300,301
<EOL>|301,302
<EOL>|303,304
History|304,311
of|312,314
Present|315,322
Illness|323,330
:|330,331
<EOL>|331,332
This|332,336
is|337,339
a|340,341
_|342,343
_|343,344
_|344,345
y|346,347
/|347,348
o|348,349
female|350,356
with|357,361
PMHx|362,366
significant|367,378
for|379,382
CAD|383,386
,|386,387
HTN|388,391
,|391,392
HLD|393,396
,|396,397
<EOL>|398,399
T2DM|399,403
,|403,404
CKD|405,408
stage|409,414
IV|415,417
,|417,418
PVD|419,422
(|423,424
s|424,425
/|425,426
p|426,427
in|428,430
_|431,432
_|432,433
_|433,434
,|434,435
left|436,440
superficial|441,452
femoral|453,460
<EOL>|461,462
artery|462,468
)|468,469
,|469,470
presents|471,479
with|480,484
lower|485,490
Left|491,495
leg|496,499
numbness|500,508
and|509,512
pain|513,517
since|518,523
<EOL>|524,525
yesterday|525,534
evening|535,542
.|542,543
The|544,547
numbness|548,556
started|557,564
last|565,569
night|570,575
in|576,578
bed|579,582
.|582,583
The|584,587
<EOL>|588,589
onset|589,594
was|595,598
gradual|599,606
,|606,607
and|608,611
it|612,614
was|615,618
associated|619,629
with|630,634
pain|635,639
/|639,640
cramping|640,648
over|649,653
<EOL>|654,655
her|655,658
lateral|659,666
calf|667,671
,|671,672
radiating|673,682
down|683,687
into|688,692
her|693,696
foot|697,701
.|701,702
She|703,706
has|707,710
had|711,714
sx|715,717
<EOL>|718,719
like|719,723
this|724,728
before|729,735
,|735,736
usually|737,744
when|745,749
resting|750,757
or|758,760
lying|761,766
in|767,769
bed|770,773
,|773,774
not|775,778
with|779,783
<EOL>|784,785
exertion|785,793
.|793,794
She|795,798
denies|799,805
leg|806,809
weakness|810,818
at|819,821
this|822,826
time|827,831
,|831,832
and|833,836
is|837,839
able|840,844
to|845,847
<EOL>|848,849
walk|849,853
without|854,861
assistance|862,872
.|872,873
Today|874,879
the|880,883
pain|884,888
and|889,892
numbness|893,901
is|902,904
<EOL>|905,906
improved|906,914
;|914,915
residual|916,924
numbness|925,933
in|934,936
her|937,940
lateral|941,948
calf|949,953
.|953,954
Denies|955,961
hx|962,964
DVT|965,968
.|968,969
<EOL>|970,971
Denies|971,977
spine|978,983
sx|984,986
:|986,987
no|988,990
trauma|991,997
,|997,998
no|999,1001
back|1002,1006
pain|1007,1011
,|1011,1012
no|1013,1015
incontinence|1016,1028
,|1028,1029
no|1030,1032
<EOL>|1033,1034
fevers|1034,1040
/|1040,1041
chills|1041,1047
.|1047,1048
No|1049,1051
numbness|1052,1060
elsewhere|1061,1070
.|1070,1071
Additionally|1072,1084
,|1084,1085
she|1086,1089
denies|1090,1096
<EOL>|1097,1098
headache|1098,1106
,|1106,1107
visual|1108,1114
changes|1115,1122
,|1122,1123
chest|1124,1129
pain|1130,1134
,|1134,1135
chest|1136,1141
pressure|1142,1150
,|1150,1151
chest|1152,1157
<EOL>|1158,1159
palpitations|1159,1171
,|1171,1172
shortness|1173,1182
of|1183,1185
breath|1186,1192
abdominal|1193,1202
pain|1203,1207
,|1207,1208
dysuria|1209,1216
,|1216,1217
or|1218,1220
<EOL>|1221,1222
diarrhea|1222,1230
.|1230,1231
<EOL>|1232,1233
<EOL>|1234,1235
Past|1235,1239
Medical|1240,1247
History|1248,1255
:|1255,1256
<EOL>|1256,1257
-|1257,1258
hypertension|1259,1271
<EOL>|1273,1274
-|1274,1275
diabetes|1276,1284
<EOL>|1286,1287
-|1287,1288
hx|1289,1291
CVA|1292,1295
(|1296,1297
cerebellar|1297,1307
-|1307,1308
medullary|1308,1317
stroke|1318,1324
in|1325,1327
_|1328,1329
_|1329,1330
_|1330,1331
<EOL>|1333,1334
-|1334,1335
CAD|1336,1339
(|1340,1341
hx|1341,1343
of|1344,1346
MI|1347,1349
in|1350,1352
_|1353,1354
_|1354,1355
_|1355,1356
BMS|1357,1360
to|1361,1363
circumflex|1364,1374
and|1375,1378
POBA|1379,1383
_|1384,1385
_|1385,1386
_|1386,1387
<EOL>|1389,1390
-|1390,1391
peripheral|1392,1402
arterial|1403,1411
disease|1412,1419
-|1419,1420
claudication|1421,1433
,|1433,1434
followed|1435,1443
by|1444,1446
<EOL>|1447,1448
vascular|1448,1456
,|1456,1457
managed|1458,1465
conservatively|1466,1480
<EOL>|1480,1481
-|1481,1482
stage|1483,1488
IV|1489,1491
CKD|1492,1495
(|1496,1497
baseline|1497,1505
2.1|1506,1509
-|1509,1510
2.6|1510,1513
)|1513,1514
<EOL>|1516,1517
-|1517,1518
GERD|1519,1523
/|1523,1524
esophageal|1524,1534
rings|1535,1540
<EOL>|1540,1541
<EOL>|1542,1543
Social|1543,1549
History|1550,1557
:|1557,1558
<EOL>|1558,1559
_|1559,1560
_|1560,1561
_|1561,1562
<EOL>|1562,1563
Family|1563,1569
History|1570,1577
:|1577,1578
<EOL>|1578,1579
Niece|1579,1584
had|1585,1588
some|1589,1593
sort|1594,1598
of|1599,1601
cancer|1602,1608
.|1608,1609
Father|1610,1616
died|1617,1621
in|1622,1624
his|1625,1628
_|1629,1630
_|1630,1631
_|1631,1632
due|1633,1636
to|1637,1639
<EOL>|1640,1641
lung|1641,1645
disease|1646,1653
.|1653,1654
Mother|1656,1662
died|1663,1667
in|1668,1670
her|1671,1674
_|1675,1676
_|1676,1677
_|1677,1678
due|1679,1682
to|1683,1685
an|1686,1688
unknown|1689,1696
cause|1697,1702
.|1702,1703
<EOL>|1705,1706
No|1706,1708
early|1709,1714
CAD|1715,1718
or|1719,1721
sudden|1722,1728
cardiac|1729,1736
death|1737,1742
.|1742,1743
No|1744,1746
other|1747,1752
known|1753,1758
history|1759,1766
of|1767,1769
<EOL>|1770,1771
cancer|1771,1777
.|1777,1778
<EOL>|1778,1779
<EOL>|1780,1781
Physical|1781,1789
Exam|1790,1794
:|1794,1795
<EOL>|1795,1796
ADMISSION|1796,1805
PHYSICAL|1806,1814
EXAM|1815,1819
:|1819,1820
<EOL>|1820,1821
<EOL>|1821,1822
Vitals|1822,1828
:|1828,1829
97.7|1830,1834
,|1834,1835
166|1836,1839
/|1839,1840
85|1840,1842
,|1842,1843
59|1844,1846
,|1846,1847
16|1848,1850
,|1850,1851
100|1852,1855
%|1855,1856
on|1857,1859
RA|1860,1862
.|1862,1863
<EOL>|1865,1866
General|1866,1873
:|1873,1874
Pleasant|1875,1883
affect|1884,1890
,|1890,1891
laying|1892,1898
in|1899,1901
bed|1902,1905
,|1905,1906
resting|1907,1914
comfortably|1915,1926
in|1927,1929
<EOL>|1930,1931
NAD|1931,1934
.|1934,1935
<EOL>|1937,1938
HEENT|1938,1943
:|1943,1944
Sclera|1945,1951
anicteric|1952,1961
,|1961,1962
MMM|1963,1966
,|1966,1967
oropharynx|1968,1978
clear|1979,1984
,|1984,1985
EOMI|1986,1990
,|1990,1991
PERRL|1992,1997
<EOL>|1999,2000
Neck|2000,2004
:|2004,2005
Supple|2006,2012
,|2012,2013
JVP|2014,2017
not|2018,2021
elevated|2022,2030
.|2030,2031
<EOL>|2033,2034
CV|2034,2036
:|2036,2037
Regular|2038,2045
rate|2046,2050
and|2051,2054
rhythm|2055,2061
,|2061,2062
normal|2063,2069
S1|2070,2072
+|2073,2074
S2|2075,2077
,|2077,2078
no|2079,2081
murmurs|2082,2089
,|2089,2090
rubs|2091,2095
,|2095,2096
<EOL>|2097,2098
gallops|2098,2105
<EOL>|2107,2108
Lungs|2108,2113
:|2113,2114
Minimal|2115,2122
bibasilar|2123,2132
crackles|2133,2141
improved|2142,2150
with|2151,2155
cough|2156,2161
.|2161,2162
<EOL>|2164,2165
Abdomen|2165,2172
:|2172,2173
obese|2174,2179
abdomen|2180,2187
,|2187,2188
soft|2189,2193
,|2193,2194
non-tender|2195,2205
,|2205,2206
non-distended|2207,2220
,|2220,2221
no|2222,2224
<EOL>|2225,2226
rebound|2226,2233
or|2234,2236
guarding|2237,2245
.|2245,2246
<EOL>|2248,2249
Ext|2249,2252
:|2252,2253
Warm|2254,2258
,|2258,2259
well|2260,2264
perfused|2265,2273
,|2273,2274
1|2275,2276
+|2276,2277
pulses|2278,2284
,|2284,2285
right|2286,2291
calf|2292,2296
swelling|2297,2305
greater|2306,2313
<EOL>|2314,2315
than|2315,2319
left|2320,2324
calf|2325,2329
swelling|2330,2338
.|2338,2339
No|2340,2342
calf|2343,2347
tenderness|2348,2358
to|2359,2361
palpation|2362,2371
.|2371,2372
Thick|2373,2378
<EOL>|2379,2380
toenails|2380,2388
,|2388,2389
dry|2390,2393
skin|2394,2398
along|2399,2404
toes|2405,2409
.|2409,2410
Hallux|2411,2417
valgus|2418,2424
.|2424,2425
<EOL>|2427,2428
Neuro|2428,2433
:|2433,2434
CNII|2435,2439
-|2439,2440
XII|2440,2443
intact|2444,2450
,|2450,2451
_|2452,2453
_|2453,2454
_|2454,2455
strength|2456,2464
upper|2465,2470
/|2470,2471
lower|2471,2476
extremities|2477,2488
,|2488,2489
<EOL>|2490,2491
grossly|2491,2498
normal|2499,2505
sensation|2506,2515
.|2515,2516
<EOL>|2517,2518
<EOL>|2518,2519
DISCHARGE|2519,2528
PHYSICAL|2529,2537
EXAM|2538,2542
<EOL>|2542,2543
Vitals|2543,2549
:|2549,2550
Tmax|2552,2556
99.1|2557,2561
HR|2562,2564
_|2565,2566
_|2566,2567
_|2567,2568
BP|2569,2571
97|2572,2574
-|2574,2575
168|2575,2578
/|2578,2579
50s|2579,2582
-|2582,2583
70s|2583,2586
RR|2587,2589
18|2590,2592
SpO2|2593,2597
<EOL>|2598,2599
97|2599,2601
-|2601,2602
100|2602,2605
%|2605,2606
RA|2606,2608
<EOL>|2608,2609
FSG|2609,2612
90|2613,2615
-|2615,2616
307|2616,2619
<EOL>|2619,2620
General|2620,2627
:|2627,2628
Pleasant|2629,2637
affect|2638,2644
,|2644,2645
laying|2646,2652
in|2653,2655
bed|2656,2659
,|2659,2660
resting|2661,2668
comfortably|2669,2680
in|2681,2683
<EOL>|2684,2685
NAD|2685,2688
.|2688,2689
<EOL>|2691,2692
HEENT|2692,2697
:|2697,2698
Sclera|2699,2705
anicteric|2706,2715
,|2715,2716
MMM|2717,2720
,|2720,2721
oropharynx|2722,2732
clear|2733,2738
,|2738,2739
EOMI|2740,2744
,|2744,2745
PERRL|2746,2751
<EOL>|2753,2754
Neck|2754,2758
:|2758,2759
Supple|2760,2766
,|2766,2767
JVP|2768,2771
not|2772,2775
elevated|2776,2784
.|2784,2785
<EOL>|2787,2788
CV|2788,2790
:|2790,2791
Regular|2792,2799
rate|2800,2804
and|2805,2808
rhythm|2809,2815
,|2815,2816
normal|2817,2823
S1|2824,2826
+|2827,2828
S2|2829,2831
,|2831,2832
no|2833,2835
murmurs|2836,2843
,|2843,2844
rubs|2845,2849
,|2849,2850
<EOL>|2851,2852
gallops|2852,2859
<EOL>|2861,2862
Lungs|2862,2867
:|2867,2868
clear|2869,2874
to|2875,2877
auscultation|2878,2890
in|2891,2893
all|2894,2897
fields|2898,2904
without|2905,2912
wheezes|2913,2920
or|2921,2923
<EOL>|2924,2925
ronchi|2925,2931
<EOL>|2931,2932
Abdomen|2932,2939
:|2939,2940
obese|2941,2946
abdomen|2947,2954
,|2954,2955
soft|2956,2960
,|2960,2961
non-tender|2962,2972
,|2972,2973
non-distended|2974,2987
,|2987,2988
no|2989,2991
<EOL>|2992,2993
rebound|2993,3000
or|3001,3003
guarding|3004,3012
.|3012,3013
<EOL>|3015,3016
Ext|3016,3019
:|3019,3020
Warm|3021,3025
,|3025,3026
well|3027,3031
perfused|3032,3040
,|3040,3041
dopplerable|3042,3053
pulses|3054,3060
_|3061,3062
_|3062,3063
_|3063,3064
on|3065,3067
RLE|3068,3071
,|3071,3072
<EOL>|3073,3074
dopplerable|3074,3085
_|3086,3087
_|3087,3088
_|3088,3089
pulse|3090,3095
on|3096,3098
LLE|3099,3102
,|3102,3103
dopplerable|3104,3115
DP|3116,3118
pulse|3119,3124
on|3125,3127
LLE|3128,3131
,|3131,3132
R|3133,3134
<EOL>|3135,3136
radial|3136,3142
pulse|3143,3148
2|3149,3150
+|3150,3151
,|3151,3152
L|3153,3154
radial|3155,3161
pulse|3162,3167
1|3168,3169
+|3169,3170
,|3170,3171
mild|3172,3176
right|3177,3182
calf|3183,3187
swelling|3188,3196
<EOL>|3197,3198
greater|3198,3205
than|3206,3210
left|3211,3215
calf|3216,3220
swelling|3221,3229
.|3229,3230
No|3231,3233
calf|3234,3238
tenderness|3239,3249
to|3250,3252
<EOL>|3253,3254
palpation|3254,3263
.|3263,3264
No|3265,3267
pain|3268,3272
to|3273,3275
palpation|3276,3285
on|3286,3288
left|3289,3293
dorsal|3294,3300
and|3301,3304
lateral|3305,3312
foot|3313,3317
<EOL>|3318,3319
-|3319,3320
callous|3321,3328
present|3329,3336
on|3337,3339
left|3340,3344
lateral|3345,3352
foot|3353,3357
.|3357,3358
Thick|3359,3364
toenails|3365,3373
,|3373,3374
dry|3375,3378
skin|3379,3383
<EOL>|3384,3385
along|3385,3390
toes|3391,3395
.|3395,3396
Non-tender|3397,3407
indurated|3408,3417
cord|3418,3422
in|3423,3425
left|3426,3430
antecubital|3431,3442
fossa|3443,3448
.|3448,3449
<EOL>|3449,3450
Neuro|3450,3455
:|3455,3456
alert|3457,3462
and|3463,3466
oriented|3467,3475
x|3476,3477
3|3478,3479
,|3479,3480
CNII|3481,3485
-|3485,3486
XII|3486,3489
intact|3490,3496
,|3496,3497
_|3498,3499
_|3499,3500
_|3500,3501
RUE|3502,3505
,|3505,3506
_|3507,3508
_|3508,3509
_|3509,3510
<EOL>|3511,3512
strength|3512,3520
LUE|3521,3524
,|3524,3525
_|3526,3527
_|3527,3528
_|3528,3529
hip|3530,3533
flexor|3534,3540
strength|3541,3549
,|3549,3550
_|3551,3552
_|3552,3553
_|3553,3554
dorsi|3555,3560
and|3561,3564
plantar|3565,3572
<EOL>|3573,3574
flexion|3574,3581
of|3582,3584
bilateral|3585,3594
lower|3595,3600
extremities|3601,3612
(|3613,3614
4|3614,3615
+|3615,3616
/|3616,3617
5|3617,3618
on|3619,3621
right|3622,3627
lower|3628,3633
<EOL>|3634,3635
extremity|3635,3644
,|3644,3645
4|3646,3647
-|3647,3648
on|3649,3651
LLE|3652,3655
)|3655,3656
,|3656,3657
fine|3658,3662
touch|3663,3668
sensation|3669,3678
on|3679,3681
extremities|3682,3693
<EOL>|3694,3695
bilaterally|3695,3706
<EOL>|3707,3708
<EOL>|3708,3709
<EOL>|3710,3711
Pertinent|3711,3720
Results|3721,3728
:|3728,3729
<EOL>|3729,3730
ADMISSION|3730,3739
LABS|3740,3744
:|3744,3745
<EOL>|3745,3746
<EOL>|3746,3747
_|3747,3748
_|3748,3749
_|3749,3750
02|3751,3753
:|3753,3754
45PM|3754,3758
BLOOD|3759,3764
WBC|3765,3768
-|3768,3769
5.1|3769,3772
RBC|3773,3776
-|3776,3777
2|3777,3778
.|3778,3779
50|3779,3781
*|3781,3782
Hgb|3783,3786
-|3786,3787
7|3787,3788
.|3788,3789
7|3789,3790
*|3790,3791
Hct|3792,3795
-|3795,3796
23|3796,3798
.|3798,3799
4|3799,3800
*|3800,3801
<EOL>|3802,3803
MCV|3803,3806
-|3806,3807
94|3807,3809
MCH|3810,3813
-|3813,3814
30.8|3814,3818
MCHC|3819,3823
-|3823,3824
32.9|3824,3828
RDW|3829,3832
-|3832,3833
14.7|3833,3837
RDWSD|3838,3843
-|3843,3844
50|3844,3846
.|3846,3847
0|3847,3848
*|3848,3849
Plt|3850,3853
_|3854,3855
_|3855,3856
_|3856,3857
<EOL>|3857,3858
_|3858,3859
_|3859,3860
_|3860,3861
02|3862,3864
:|3864,3865
45PM|3865,3869
BLOOD|3870,3875
Neuts|3876,3881
-|3881,3882
74|3882,3884
.|3884,3885
4|3885,3886
*|3886,3887
Lymphs|3888,3894
-|3894,3895
15|3895,3897
.|3897,3898
1|3898,3899
*|3899,3900
Monos|3901,3906
-|3906,3907
7.7|3907,3910
<EOL>|3911,3912
Eos|3912,3915
-|3915,3916
2.4|3916,3919
Baso|3920,3924
-|3924,3925
0.2|3925,3928
Im|3929,3931
_|3932,3933
_|3933,3934
_|3934,3935
AbsNeut|3936,3943
-|3943,3944
3|3944,3945
.|3945,3946
79|3946,3948
AbsLymp|3949,3956
-|3956,3957
0|3957,3958
.|3958,3959
77|3959,3961
*|3961,3962
<EOL>|3963,3964
AbsMono|3964,3971
-|3971,3972
0|3972,3973
.|3973,3974
39|3974,3976
AbsEos|3977,3983
-|3983,3984
0|3984,3985
.|3985,3986
12|3986,3988
AbsBaso|3989,3996
-|3996,3997
0.01|3997,4001
<EOL>|4001,4002
_|4002,4003
_|4003,4004
_|4004,4005
02|4006,4008
:|4008,4009
45PM|4009,4013
BLOOD|4014,4019
_|4020,4021
_|4021,4022
_|4022,4023
PTT|4024,4027
-|4027,4028
26.1|4028,4032
_|4033,4034
_|4034,4035
_|4035,4036
<EOL>|4036,4037
_|4037,4038
_|4038,4039
_|4039,4040
02|4041,4043
:|4043,4044
45PM|4044,4048
BLOOD|4049,4054
Glucose|4055,4062
-|4062,4063
107|4063,4066
*|4066,4067
UreaN|4068,4073
-|4073,4074
72|4074,4076
*|4076,4077
Creat|4078,4083
-|4083,4084
2|4084,4085
.|4085,4086
9|4086,4087
*|4087,4088
Na|4089,4091
-|4091,4092
141|4092,4095
<EOL>|4096,4097
K|4097,4098
-|4098,4099
4.3|4099,4102
Cl|4103,4105
-|4105,4106
108|4106,4109
HCO3|4110,4114
-|4114,4115
21|4115,4117
*|4117,4118
AnGap|4119,4124
-|4124,4125
16|4125,4127
<EOL>|4127,4128
_|4128,4129
_|4129,4130
_|4130,4131
02|4132,4134
:|4134,4135
45PM|4135,4139
BLOOD|4140,4145
calTIBC|4146,4153
-|4153,4154
303|4154,4157
Ferritn|4158,4165
-|4165,4166
153|4166,4169
*|4169,4170
TRF|4171,4174
-|4174,4175
233|4175,4178
<EOL>|4178,4179
<EOL>|4179,4180
PERTINENT|4180,4189
LABS|4190,4194
/|4194,4195
IMAGING|4195,4202
:|4202,4203
<EOL>|4203,4204
<EOL>|4204,4205
-|4205,4206
She|4206,4209
received|4210,4218
1U|4219,4221
pRBCs|4222,4227
on|4228,4230
admission|4231,4240
on|4241,4243
_|4244,4245
_|4245,4246
_|4246,4247
07|4248,4250
:|4250,4251
00AM|4251,4255
BLOOD|4256,4261
WBC|4262,4265
-|4265,4266
6.0|4266,4269
RBC|4270,4273
-|4273,4274
2|4274,4275
.|4275,4276
83|4276,4278
*|4278,4279
Hgb|4280,4283
-|4283,4284
8|4284,4285
.|4285,4286
7|4286,4287
*|4287,4288
Hct|4289,4292
-|4292,4293
26|4293,4295
.|4295,4296
3|4296,4297
*|4297,4298
<EOL>|4299,4300
MCV|4300,4303
-|4303,4304
93|4304,4306
MCH|4307,4310
-|4310,4311
30.7|4311,4315
MCHC|4316,4320
-|4320,4321
33.1|4321,4325
RDW|4326,4329
-|4329,4330
14.7|4330,4334
RDWSD|4335,4340
-|4340,4341
50|4341,4343
.|4343,4344
2|4344,4345
*|4345,4346
Plt|4347,4350
_|4351,4352
_|4352,4353
_|4353,4354
<EOL>|4354,4355
-|4355,4356
She|4356,4359
had|4360,4363
one|4364,4367
large|4368,4373
episode|4374,4381
of|4382,4384
coffee|4385,4391
ground|4392,4398
emesis|4399,4405
-|4405,4406
<EOL>|4406,4407
_|4407,4408
_|4408,4409
_|4409,4410
05|4411,4413
:|4413,4414
10PM|4414,4418
BLOOD|4419,4424
WBC|4425,4428
-|4428,4429
5.6|4429,4432
RBC|4433,4436
-|4436,4437
2|4437,4438
.|4438,4439
44|4439,4441
*|4441,4442
Hgb|4443,4446
-|4446,4447
7|4447,4448
.|4448,4449
4|4449,4450
*|4450,4451
Hct|4452,4455
-|4455,4456
22|4456,4458
.|4458,4459
7|4459,4460
*|4460,4461
<EOL>|4462,4463
MCV|4463,4466
-|4466,4467
93|4467,4469
MCH|4470,4473
-|4473,4474
30.3|4474,4478
MCHC|4479,4483
-|4483,4484
32.6|4484,4488
RDW|4489,4492
-|4492,4493
14.7|4493,4497
RDWSD|4498,4503
-|4503,4504
49|4504,4506
.|4506,4507
8|4507,4508
*|4508,4509
Plt|4510,4513
_|4514,4515
_|4515,4516
_|4516,4517
<EOL>|4517,4518
-|4518,4519
She|4519,4522
received|4523,4531
500cc|4532,4537
NS|4538,4540
and|4541,4544
2UpRBCs|4545,4552
-|4552,4553
<EOL>|4553,4554
_|4554,4555
_|4555,4556
_|4556,4557
07|4558,4560
:|4560,4561
45AM|4561,4565
BLOOD|4566,4571
WBC|4572,4575
-|4575,4576
5.7|4576,4579
RBC|4580,4583
-|4583,4584
3|4584,4585
.|4585,4586
49|4586,4588
*|4588,4589
#|4589,4590
Hgb|4591,4594
-|4594,4595
10|4595,4597
.|4597,4598
7|4598,4599
*|4599,4600
#|4600,4601
Hct|4602,4605
-|4605,4606
32|4606,4608
.|4608,4609
3|4609,4610
*|4610,4611
<EOL>|4612,4613
MCV|4613,4616
-|4616,4617
93|4617,4619
MCH|4620,4623
-|4623,4624
30.7|4624,4628
MCHC|4629,4633
-|4633,4634
33.1|4634,4638
RDW|4639,4642
-|4642,4643
14.9|4643,4647
RDWSD|4648,4653
-|4653,4654
49|4654,4656
.|4656,4657
1|4657,4658
*|4658,4659
Plt|4660,4663
_|4664,4665
_|4665,4666
_|4666,4667
<EOL>|4667,4668
<EOL>|4668,4669
_|4669,4670
_|4670,4671
_|4671,4672
bilateral|4673,4682
lower|4683,4688
extremity|4689,4698
doppler|4699,4706
U|4707,4708
/|4708,4709
S|4709,4710
<EOL>|4710,4711
IMPRESSION|4711,4721
:|4721,4722
<EOL>|4724,4725
1.|4725,4727
Deep|4729,4733
venous|4734,4740
thrombosis|4741,4751
in|4752,4754
the|4755,4758
bilateral|4759,4768
posterior|4769,4778
tibial|4779,4785
<EOL>|4786,4787
veins|4787,4792
.|4792,4793
<EOL>|4794,4795
2.|4795,4797
2.0|4799,4802
x|4803,4804
1.3|4805,4808
x|4809,4810
1.8|4811,4814
cm|4815,4817
right|4818,4823
-|4823,4824
sided|4824,4829
_|4830,4831
_|4831,4832
_|4832,4833
cyst|4834,4838
.|4838,4839
<EOL>|4840,4841
<EOL>|4841,4842
EGD|4842,4845
_|4846,4847
_|4847,4848
_|4848,4849
<EOL>|4849,4850
Small|4850,4855
amount|4856,4862
of|4863,4865
hematin|4866,4873
without|4874,4881
evidence|4882,4890
of|4891,4893
ulceration|4894,4904
or|4905,4907
active|4908,4914
<EOL>|4915,4916
bleeding|4916,4924
seen|4925,4929
at|4930,4932
the|4933,4936
GE|4937,4939
junction|4940,4948
.|4948,4949
<EOL>|4949,4950
The|4950,4953
stomach|4954,4961
is|4962,4964
significantly|4965,4978
deformed|4979,4987
.|4987,4988
Diffuse|4989,4996
erythema|4997,5005
and|5006,5009
<EOL>|5010,5011
superficial|5011,5022
ulcerations|5023,5034
in|5035,5037
the|5038,5041
stomach|5042,5049
consistent|5050,5060
with|5061,5065
severe|5066,5072
<EOL>|5073,5074
gastritis|5074,5083
.|5083,5084
No|5085,5087
active|5088,5094
bleeding|5095,5103
identified|5104,5114
.|5114,5115
<EOL>|5115,5116
Medium|5116,5122
hiatal|5123,5129
hernia|5130,5136
<EOL>|5136,5137
Erythema|5137,5145
and|5146,5149
superficial|5150,5161
ulcerations|5162,5173
in|5174,5176
the|5177,5180
duodenal|5181,5189
bulb|5190,5194
<EOL>|5195,5196
consistent|5196,5206
with|5207,5211
duodenitis|5212,5222
.|5222,5223
<EOL>|5223,5224
Otherwise|5224,5233
normal|5234,5240
EGD|5241,5244
to|5245,5247
third|5248,5253
part|5254,5258
of|5259,5261
the|5262,5265
duodenum|5266,5274
<EOL>|5274,5275
<EOL>|5275,5276
_|5276,5277
_|5277,5278
_|5278,5279
Left|5280,5284
upper|5285,5290
extremity|5291,5300
ultrasound|5301,5311
<EOL>|5311,5312
IMPRESSION|5312,5322
:|5322,5323
<EOL>|5325,5326
1|5326,5327
.|5327,5328
No|5330,5332
evidence|5333,5341
of|5342,5344
deep|5345,5349
vein|5350,5354
thrombosis|5355,5365
in|5366,5368
the|5369,5372
left|5373,5377
upper|5378,5383
<EOL>|5384,5385
extremity|5385,5394
.|5394,5395
<EOL>|5396,5397
2.|5397,5399
Likely|5401,5407
evolving|5408,5416
hematoma|5417,5425
in|5426,5428
the|5429,5432
left|5433,5437
antecubital|5438,5449
fossa|5450,5455
.|5455,5456
<EOL>|5457,5458
<EOL>|5458,5459
_|5459,5460
_|5460,5461
_|5461,5462
CT|5463,5465
head|5466,5470
non|5471,5474
contrast|5475,5483
<EOL>|5483,5484
IMPRESSION|5484,5494
:|5494,5495
1|5496,5497
.|5497,5498
No|5499,5501
evidence|5502,5510
of|5511,5513
acute|5514,5519
infarction|5520,5530
,|5530,5531
hemorrhage|5532,5542
,|5542,5543
<EOL>|5544,5545
fractures|5545,5554
.|5554,5555
<EOL>|5556,5557
<EOL>|5557,5558
DISCHARGE|5558,5567
LABS|5568,5572
:|5572,5573
<EOL>|5573,5574
_|5574,5575
_|5575,5576
_|5576,5577
07|5578,5580
:|5580,5581
30AM|5581,5585
BLOOD|5586,5591
WBC|5592,5595
-|5595,5596
5.8|5596,5599
RBC|5600,5603
-|5603,5604
2|5604,5605
.|5605,5606
44|5606,5608
*|5608,5609
Hgb|5610,5613
-|5613,5614
7|5614,5615
.|5615,5616
4|5616,5617
*|5617,5618
Hct|5619,5622
-|5622,5623
22|5623,5625
.|5625,5626
9|5626,5627
*|5627,5628
<EOL>|5629,5630
MCV|5630,5633
-|5633,5634
94|5634,5636
MCH|5637,5640
-|5640,5641
30.3|5641,5645
MCHC|5646,5650
-|5650,5651
32.3|5651,5655
RDW|5656,5659
-|5659,5660
14.6|5660,5664
RDWSD|5665,5670
-|5670,5671
50|5671,5673
.|5673,5674
2|5674,5675
*|5675,5676
Plt|5677,5680
_|5681,5682
_|5682,5683
_|5683,5684
<EOL>|5684,5685
_|5685,5686
_|5686,5687
_|5687,5688
07|5689,5691
:|5691,5692
30AM|5692,5696
BLOOD|5697,5702
Plt|5703,5706
_|5707,5708
_|5708,5709
_|5709,5710
<EOL>|5710,5711
_|5711,5712
_|5712,5713
_|5713,5714
07|5715,5717
:|5717,5718
30AM|5718,5722
BLOOD|5723,5728
Glucose|5729,5736
-|5736,5737
78|5737,5739
UreaN|5740,5745
-|5745,5746
45|5746,5748
*|5748,5749
Creat|5750,5755
-|5755,5756
1|5756,5757
.|5757,5758
7|5758,5759
*|5759,5760
Na|5761,5763
-|5763,5764
142|5764,5767
<EOL>|5768,5769
K|5769,5770
-|5770,5771
4.7|5771,5774
Cl|5775,5777
-|5777,5778
109|5778,5781
*|5781,5782
HCO3|5783,5787
-|5787,5788
20|5788,5790
*|5790,5791
AnGap|5792,5797
-|5797,5798
18|5798,5800
<EOL>|5800,5801
_|5801,5802
_|5802,5803
_|5803,5804
:|5804,5805
30AM|5805,5809
BLOOD|5810,5815
Calcium|5816,5823
-|5823,5824
9.4|5824,5827
Phos|5828,5832
-|5832,5833
4.5|5833,5836
Mg|5837,5839
-|5839,5840
2.0|5840,5843
<EOL>|5843,5844
_|5844,5845
_|5845,5846
_|5846,5847
07|5848,5850
:|5850,5851
30AM|5851,5855
BLOOD|5856,5861
EDTA|5862,5866
_|5867,5868
_|5868,5869
_|5869,5870
<EOL>|5870,5871
<EOL>|5872,5873
Brief|5873,5878
Hospital|5879,5887
Course|5888,5894
:|5894,5895
<EOL>|5895,5896
Outpatient|5896,5906
Providers|5907,5916
:|5916,5917
_|5918,5919
_|5919,5920
_|5920,5921
with|5922,5926
PMHx|5927,5931
significant|5932,5943
for|5944,5947
CAD|5948,5951
,|5951,5952
HTN|5953,5956
,|5956,5957
<EOL>|5958,5959
HLD|5959,5962
,|5962,5963
T2DM|5964,5968
,|5968,5969
CKD|5970,5973
stage|5974,5979
IV|5980,5982
,|5982,5983
PVD|5984,5987
(|5988,5989
s|5989,5990
/|5990,5991
p|5991,5992
in|5993,5995
_|5996,5997
_|5997,5998
_|5998,5999
,|5999,6000
left|6001,6005
superficial|6006,6017
<EOL>|6018,6019
femoral|6019,6026
artery|6027,6033
)|6033,6034
,|6034,6035
presents|6036,6044
with|6045,6049
lower|6050,6055
left|6056,6060
leg|6061,6064
numbness|6065,6073
and|6074,6077
pain|6078,6082
,|6082,6083
<EOL>|6084,6085
found|6085,6090
to|6091,6093
have|6094,6098
bilateral|6099,6108
unprovoked|6109,6119
DVT|6120,6123
.|6123,6124
She|6125,6128
was|6129,6132
treated|6133,6140
with|6141,6145
a|6146,6147
<EOL>|6148,6149
heparin|6149,6156
drip|6157,6161
and|6162,6165
had|6166,6169
many|6170,6174
bleeding|6175,6183
events|6184,6190
during|6191,6197
her|6198,6201
stay|6202,6206
:|6206,6207
she|6208,6211
<EOL>|6212,6213
developed|6213,6222
an|6223,6225
upper|6226,6231
GIB|6232,6235
,|6235,6236
had|6237,6240
an|6241,6243
EGD|6244,6247
,|6247,6248
and|6249,6252
was|6253,6256
followed|6257,6265
by|6266,6268
GI|6269,6271
<EOL>|6272,6273
during|6273,6279
her|6280,6283
admission|6284,6293
.|6293,6294
The|6295,6298
heparin|6299,6306
drip|6307,6311
was|6312,6315
stopped|6316,6323
and|6324,6327
then|6328,6332
<EOL>|6333,6334
re-started|6334,6344
once|6345,6349
her|6350,6353
coffee|6354,6360
-|6360,6361
ground|6361,6367
emesis|6368,6374
resolved|6375,6383
.|6383,6384
Her|6385,6388
stools|6389,6395
<EOL>|6396,6397
were|6397,6401
guiac|6402,6407
positive|6408,6416
,|6416,6417
however|6418,6425
no|6426,6428
active|6429,6435
blood|6436,6441
was|6442,6445
found|6446,6451
on|6452,6454
rectal|6455,6461
<EOL>|6462,6463
exam|6463,6467
.|6467,6468
GI|6469,6471
felt|6472,6476
that|6477,6481
colonoscopy|6482,6493
could|6494,6499
be|6500,6502
deferred|6503,6511
to|6512,6514
out|6515,6518
patient|6519,6526
.|6526,6527
<EOL>|6528,6529
Additionally|6529,6541
she|6542,6545
developed|6546,6555
a|6556,6557
left|6558,6562
arm|6563,6566
hematoma|6567,6575
.|6575,6576
The|6577,6580
heparin|6581,6588
drip|6589,6593
<EOL>|6594,6595
was|6595,6598
stopped|6599,6606
and|6607,6610
then|6611,6615
re-started|6616,6626
once|6627,6631
her|6632,6635
hematoma|6636,6644
was|6645,6648
felt|6649,6653
to|6654,6656
be|6657,6659
<EOL>|6660,6661
stable|6661,6667
.|6667,6668
She|6669,6672
had|6673,6676
left|6677,6681
radial|6682,6688
as|6689,6691
well|6692,6696
as|6697,6699
bilateral|6700,6709
lower|6710,6715
extremity|6716,6725
<EOL>|6726,6727
_|6727,6728
_|6728,6729
_|6729,6730
dopplerable|6731,6742
pulses|6743,6749
throughout|6750,6760
admission|6761,6770
.|6770,6771
Hematology|6772,6782
was|6783,6786
<EOL>|6787,6788
consulted|6788,6797
after|6798,6803
the|6804,6807
patient|6808,6815
developed|6816,6825
a|6826,6827
left|6828,6832
arm|6833,6836
hematoma|6837,6845
and|6846,6849
<EOL>|6850,6851
the|6851,6854
drip|6855,6859
was|6860,6863
slowly|6864,6870
uptitrated|6871,6881
as|6882,6884
per|6885,6888
their|6889,6894
recommendations|6895,6910
.|6910,6911
She|6912,6915
<EOL>|6916,6917
was|6917,6920
successfully|6921,6933
bridged|6934,6941
to|6942,6944
coumadin|6945,6953
with|6954,6958
an|6959,6961
INR|6962,6965
on|6966,6968
discharge|6969,6978
of|6979,6981
<EOL>|6982,6983
2.0|6983,6986
.|6986,6987
She|6988,6991
was|6992,6995
discharged|6996,7006
to|7007,7009
rehab|7010,7015
as|7016,7018
per|7019,7022
_|7023,7024
_|7024,7025
_|7025,7026
recs|7027,7031
.|7031,7032
<EOL>|7033,7034
<EOL>|7034,7035
Please|7035,7041
see|7042,7045
below|7046,7051
for|7052,7055
a|7056,7057
more|7058,7062
problem|7063,7070
based|7071,7076
/|7076,7077
detailed|7077,7085
summary|7086,7093
and|7094,7097
<EOL>|7098,7099
transitional|7099,7111
issues|7112,7118
.|7118,7119
<EOL>|7119,7120
<EOL>|7120,7121
=|7121,7122
<EOL>|7122,7123
=|7123,7124
<EOL>|7124,7125
=|7125,7126
<EOL>|7126,7127
=|7127,7128
<EOL>|7128,7129
=|7129,7130
<EOL>|7130,7131
=|7131,7132
<EOL>|7132,7133
=|7133,7134
<EOL>|7134,7135
=|7135,7136
<EOL>|7136,7137
=|7137,7138
<EOL>|7138,7139
=|7139,7140
<EOL>|7140,7141
=|7141,7142
<EOL>|7142,7143
=|7143,7144
<EOL>|7144,7145
=|7145,7146
<EOL>|7146,7147
=|7147,7148
<EOL>|7148,7149
=|7149,7150
<EOL>|7150,7151
=|7151,7152
<EOL>|7152,7153
=|7153,7154
<EOL>|7154,7155
=|7155,7156
<EOL>|7156,7157
=|7157,7158
=|7158,7159
=|7159,7160
=|7160,7161
=|7161,7162
=|7162,7163
=|7163,7164
=|7164,7165
=|7165,7166
=|7166,7167
=|7167,7168
=|7168,7169
=|7169,7170
=|7170,7171
=|7171,7172
=|7172,7173
=|7173,7174
=|7174,7175
=|7175,7176
=|7176,7177
=|7177,7178
=|7178,7179
=|7179,7180
=|7180,7181
=|7181,7182
=|7182,7183
=|7183,7184
=|7184,7185
=|7185,7186
=|7186,7187
=|7187,7188
=|7188,7189
=|7189,7190
=|7190,7191
=|7191,7192
=|7192,7193
=|7193,7194
=|7194,7195
=|7195,7196
=|7196,7197
=|7197,7198
=|7198,7199
=|7199,7200
=|7200,7201
=|7201,7202
=|7202,7203
=|7203,7204
=|7204,7205
=|7205,7206
=|7206,7207
=|7207,7208
=|7208,7209
=|7209,7210
=|7210,7211
=|7211,7212
=|7212,7213
=|7213,7214
=|7214,7215
=|7215,7216
=|7216,7217
=|7217,7218
=|7218,7219
=|7219,7220
=|7220,7221
<EOL>|7221,7222
<EOL>|7222,7223
_|7223,7224
_|7224,7225
_|7225,7226
y|7227,7228
/|7228,7229
o|7229,7230
female|7231,7237
with|7238,7242
PMHx|7243,7247
significant|7248,7259
for|7260,7263
CAD|7264,7267
,|7267,7268
HTN|7269,7272
,|7272,7273
HLD|7274,7277
,|7277,7278
T2DM|7279,7283
,|7283,7284
CKD|7285,7288
<EOL>|7289,7290
stage|7290,7295
IV|7296,7298
,|7298,7299
PVD|7300,7303
(|7304,7305
s|7305,7306
/|7306,7307
p|7307,7308
in|7309,7311
_|7312,7313
_|7313,7314
_|7314,7315
,|7315,7316
left|7317,7321
superficial|7322,7333
femoral|7334,7341
artery|7342,7348
)|7348,7349
,|7349,7350
<EOL>|7351,7352
presented|7352,7361
with|7362,7366
lower|7367,7372
Left|7373,7377
leg|7378,7381
numbness|7382,7390
and|7391,7394
pain|7395,7399
since|7400,7405
yesterday|7406,7415
<EOL>|7416,7417
evening|7417,7424
,|7424,7425
with|7426,7430
ultrasound|7431,7441
bilateral|7442,7451
lower|7452,7457
extremities|7458,7469
showing|7470,7477
<EOL>|7478,7479
bilateral|7479,7488
posterior|7489,7498
tibial|7499,7505
veins|7506,7511
DVT|7512,7515
's|7515,7517
.|7517,7518
<EOL>|7518,7519
<EOL>|7519,7520
#|7520,7521
Unprovoked|7522,7532
Bilateral|7533,7542
DVTs|7543,7547
:|7547,7548
No|7549,7551
clinical|7552,7560
signs|7561,7566
of|7567,7569
PE|7570,7572
on|7573,7575
<EOL>|7576,7577
admission|7577,7586
or|7587,7589
during|7590,7596
stay|7597,7601
,|7601,7602
positive|7603,7611
bilateral|7612,7621
DVTs|7622,7626
on|7627,7629
LENIs|7630,7635
.|7635,7636
Pain|7637,7641
<EOL>|7642,7643
and|7643,7646
swelling|7647,7655
improved|7656,7664
on|7665,7667
anticoagulation|7668,7683
.|7683,7684
Patient|7685,7692
was|7693,7696
bridged|7697,7704
<EOL>|7705,7706
with|7706,7710
heparin|7711,7718
drip|7719,7723
to|7724,7726
therapeutic|7727,7738
warfarin|7739,7747
with|7748,7752
INR|7753,7756
goal|7757,7761
_|7762,7763
_|7763,7764
_|7764,7765
.|7765,7766
Due|7767,7770
<EOL>|7771,7772
to|7772,7774
continually|7775,7786
supratherapeutic|7787,7803
PTT|7804,7807
>|7808,7809
150|7810,7813
on|7814,7816
heparin|7817,7824
drip|7825,7829
,|7829,7830
<EOL>|7831,7832
hematology|7832,7842
was|7843,7846
consulted|7847,7856
and|7857,7860
no|7861,7863
further|7864,7871
workup|7872,7878
was|7879,7882
deemed|7883,7889
<EOL>|7890,7891
necessary|7891,7900
.|7900,7901
Heparin|7902,7909
drip|7910,7914
was|7915,7918
carefully|7919,7928
uptitrated|7929,7939
as|7940,7942
needed|7943,7949
.|7949,7950
<EOL>|7951,7952
Clopidogrel|7952,7963
was|7964,7967
stopped|7968,7975
per|7976,7979
outpatient|7980,7990
cardiologist|7991,8003
.|8003,8004
Patient|8005,8012
<EOL>|8013,8014
will|8014,8018
need|8019,8023
age|8024,8027
-|8027,8028
appropriate|8028,8039
cancer|8040,8046
screening|8047,8056
including|8057,8066
colonoscopy|8067,8078
<EOL>|8079,8080
and|8080,8083
mammogram|8084,8093
.|8093,8094
Patient|8095,8102
will|8103,8107
follow|8108,8114
-|8114,8115
up|8115,8117
in|8118,8120
_|8121,8122
_|8122,8123
_|8123,8124
clinic|8125,8131
for|8132,8135
<EOL>|8136,8137
anticoagulation|8137,8152
management|8153,8163
and|8164,8167
should|8168,8174
continue|8175,8183
on|8184,8186
warfarin|8187,8195
for|8196,8199
<EOL>|8200,8201
at|8201,8203
least|8204,8209
3|8210,8211
months|8212,8218
.|8218,8219
<EOL>|8220,8221
<EOL>|8221,8222
#|8222,8223
Upper|8224,8229
GI|8230,8232
bleed|8233,8238
:|8238,8239
Patient|8240,8247
developed|8248,8257
1|8258,8259
episode|8260,8267
large|8268,8273
coffee|8274,8280
<EOL>|8281,8282
ground|8282,8288
emesis|8289,8295
while|8296,8301
on|8302,8304
heparin|8305,8312
drip|8313,8317
with|8318,8322
PTT|8323,8326
>|8327,8328
150|8329,8332
.|8332,8333
Received|8334,8342
2U|8343,8345
<EOL>|8346,8347
pRBCs|8347,8352
.|8352,8353
GI|8354,8356
consulted|8357,8366
and|8367,8370
EGD|8371,8374
showed|8375,8381
gastritis|8382,8391
and|8392,8395
superficial|8396,8407
<EOL>|8408,8409
erosions|8409,8417
but|8418,8421
no|8422,8424
active|8425,8431
bleeding|8432,8440
.|8440,8441
Incidental|8442,8452
finding|8453,8460
of|8461,8463
medium|8464,8470
<EOL>|8471,8472
sized|8472,8477
hiatal|8478,8484
hernia|8485,8491
.|8491,8492
Stool|8493,8498
h.|8499,8501
pylori|8502,8508
antigen|8509,8516
was|8517,8520
negative|8521,8529
.|8529,8530
GI|8531,8533
<EOL>|8534,8535
recommended|8535,8546
8|8547,8548
weeks|8549,8554
of|8555,8557
high|8558,8562
dose|8563,8567
PPI|8568,8571
.|8571,8572
<EOL>|8572,8573
<EOL>|8573,8574
#|8574,8575
Left|8576,8580
antecubital|8581,8592
hematoma|8593,8601
:|8601,8602
Patient|8603,8610
developed|8611,8620
large|8621,8626
left|8627,8631
<EOL>|8632,8633
antecubital|8633,8644
hematoma|8645,8653
in|8654,8656
setting|8657,8664
of|8665,8667
phlebotomy|8668,8678
and|8679,8682
PTT|8683,8686
>|8687,8688
150|8689,8692
on|8693,8695
<EOL>|8696,8697
heparin|8697,8704
gtt|8705,8708
.|8708,8709
Heparin|8710,8717
gtt|8718,8721
held|8722,8726
while|8727,8732
hematoma|8733,8741
improved|8742,8750
.|8750,8751
Repeat|8752,8758
<EOL>|8759,8760
h|8760,8761
/|8761,8762
h|8762,8763
were|8764,8768
stable|8769,8775
.|8775,8776
<EOL>|8777,8778
<EOL>|8778,8779
#|8779,8780
Acute|8781,8786
on|8787,8789
CKD|8790,8793
Stage|8794,8799
IV|8800,8802
:|8802,8803
Patient|8804,8811
with|8812,8816
creatinine|8817,8827
of|8828,8830
2.9|8831,8834
on|8835,8837
<EOL>|8838,8839
admission|8839,8848
with|8849,8853
baseline|8854,8862
2.0|8863,8866
-|8866,8867
2.5|8867,8870
.|8870,8871
Improved|8872,8880
with|8881,8885
hydration|8886,8895
.|8895,8896
Home|8897,8901
<EOL>|8902,8903
lasix|8903,8908
and|8909,8912
lisinopril|8913,8923
were|8924,8928
initially|8929,8938
held|8939,8943
.|8943,8944
Home|8945,8949
lasix|8950,8955
restarted|8956,8965
<EOL>|8966,8967
on|8967,8969
discharge|8970,8979
at|8980,8982
20mg|8983,8987
daily|8988,8993
.|8993,8994
<EOL>|8995,8996
<EOL>|8996,8997
#|8997,8998
Normocytic|8999,9009
Anemia|9010,9016
:|9016,9017
Patient|9018,9025
has|9026,9029
normocytic|9030,9040
anemia|9041,9047
.|9047,9048
Rectal|9049,9055
exam|9056,9060
<EOL>|9061,9062
in|9062,9064
ED|9065,9067
was|9068,9071
guaiac|9072,9078
negative|9079,9087
.|9087,9088
In|9089,9091
past|9092,9096
treated|9097,9104
with|9105,9109
aransep|9110,9117
as|9118,9120
well|9121,9125
<EOL>|9126,9127
as|9127,9129
EPO|9130,9133
.|9133,9134
Etiology|9135,9143
likely|9144,9150
related|9151,9158
to|9159,9161
underlying|9162,9172
CKD|9173,9176
,|9176,9177
however|9178,9185
also|9186,9190
<EOL>|9191,9192
must|9192,9196
consider|9197,9205
slow|9206,9210
GI|9211,9213
bleed|9214,9219
(|9220,9221
patient|9221,9228
has|9229,9232
gastritis|9233,9242
/|9242,9243
duodenitis|9243,9253
on|9254,9256
<EOL>|9257,9258
EGD|9258,9261
but|9262,9265
no|9266,9268
evidence|9269,9277
of|9278,9280
active|9281,9287
bleeding|9288,9296
.|9296,9297
Iron|9298,9302
studies|9303,9310
were|9311,9315
<EOL>|9316,9317
normal|9317,9323
.|9323,9324
<EOL>|9325,9326
<EOL>|9326,9327
#|9327,9328
HFpEF|9329,9334
:|9334,9335
Home|9336,9340
furosemide|9341,9351
and|9352,9355
Lisinopril|9356,9366
were|9367,9371
held|9372,9376
on|9377,9379
admission|9380,9389
<EOL>|9390,9391
for|9391,9394
_|9395,9396
_|9396,9397
_|9397,9398
followed|9399,9407
by|9408,9410
GI|9411,9413
bleed|9414,9419
.|9419,9420
Carvedilol|9421,9431
and|9432,9435
nifedine|9436,9444
were|9445,9449
held|9450,9454
<EOL>|9455,9456
in|9456,9458
setting|9459,9466
of|9467,9469
GIB|9470,9473
(|9474,9475
see|9475,9478
above|9479,9484
)|9484,9485
.|9485,9486
Nifedipine|9487,9497
was|9498,9501
restarted|9502,9511
at|9512,9514
30mg|9515,9519
<EOL>|9520,9521
bid|9521,9524
and|9525,9528
lasix|9529,9534
was|9535,9538
decreased|9539,9548
from|9549,9553
40mg|9554,9558
to|9559,9561
20mg|9562,9566
daily|9567,9572
.|9572,9573
<EOL>|9573,9574
<EOL>|9574,9575
#|9575,9576
CAD|9577,9580
:|9580,9581
hx|9582,9584
of|9585,9587
MI|9588,9590
in|9591,9593
_|9594,9595
_|9595,9596
_|9596,9597
BMS|9598,9601
to|9602,9604
circumflex|9605,9615
and|9616,9619
POBA|9620,9624
_|9625,9626
_|9626,9627
_|9627,9628
.|9628,9629
Per|9630,9633
<EOL>|9634,9635
discussions|9635,9646
with|9647,9651
Dr.|9652,9655
_|9656,9657
_|9657,9658
_|9658,9659
,|9659,9660
patient|9661,9668
's|9668,9670
cardiologist|9671,9683
,|9683,9684
<EOL>|9685,9686
clopidogrel|9686,9697
was|9698,9701
held|9702,9706
given|9707,9712
GI|9713,9715
bleed|9716,9721
and|9722,9725
initiation|9726,9736
of|9737,9739
warfarin|9740,9748
.|9748,9749
<EOL>|9750,9751
Lasix|9751,9756
initially|9757,9766
held|9767,9771
as|9772,9774
above|9775,9780
,|9780,9781
but|9782,9785
restarted|9786,9795
on|9796,9798
discharge|9799,9808
at|9809,9811
<EOL>|9812,9813
20mg|9813,9817
daily|9818,9823
.|9823,9824
Home|9825,9829
ASA|9830,9833
,|9833,9834
statin|9835,9841
,|9841,9842
and|9843,9846
carvedilol|9847,9857
were|9858,9862
continued|9863,9872
.|9872,9873
<EOL>|9874,9875
<EOL>|9875,9876
#|9876,9877
HTN|9878,9881
:|9881,9882
Nifedipine|9883,9893
was|9894,9897
decreased|9898,9907
to|9908,9910
30mg|9911,9915
BID|9916,9919
from|9920,9924
60mg|9925,9929
BID|9930,9933
given|9934,9939
<EOL>|9940,9941
multiple|9941,9949
bleeding|9950,9958
episodes|9959,9967
and|9968,9971
normal|9972,9978
blood|9979,9984
pressures|9985,9994
.|9994,9995
Home|9996,10000
<EOL>|10001,10002
carvedilol|10002,10012
continued|10013,10022
.|10022,10023
Patient|10024,10031
's|10031,10033
nifedipine|10034,10044
was|10045,10048
decreased|10049,10058
to|10059,10061
30mg|10062,10066
<EOL>|10067,10068
daily|10068,10073
given|10074,10079
acute|10080,10085
bleed|10086,10091
and|10092,10095
SBPs|10096,10100
in|10101,10103
the|10104,10107
_|10108,10109
_|10109,10110
_|10110,10111
<EOL>|10111,10112
Lasix|10112,10117
was|10118,10121
decreased|10122,10131
from|10132,10136
40|10137,10139
daily|10140,10145
to|10146,10148
20|10149,10151
daily|10152,10157
.|10157,10158
<EOL>|10158,10159
<EOL>|10160,10161
#|10161,10162
Diabetes|10163,10171
Mellitus|10172,10180
:|10180,10181
Stable|10182,10188
on|10189,10191
home|10192,10196
30|10197,10199
units|10200,10205
70|10206,10208
/|10208,10209
30|10209,10211
insulin|10212,10219
at|10220,10222
<EOL>|10223,10224
bedtime|10224,10231
.|10231,10232
<EOL>|10234,10235
<EOL>|10235,10236
TRANSITIONAL|10236,10248
ISSUES|10249,10255
:|10255,10256
<EOL>|10256,10257
-|10257,10258
Out|10259,10262
patient|10263,10270
hypercoaguability|10271,10288
work|10289,10293
up|10294,10296
including|10297,10306
screening|10307,10316
<EOL>|10317,10318
colonoscopy|10318,10329
(|10330,10331
last|10331,10335
in|10336,10338
_|10339,10340
_|10340,10341
_|10341,10342
and|10343,10346
mammogram|10347,10356
<EOL>|10356,10357
-|10357,10358
Patient|10359,10366
will|10367,10371
need|10372,10376
to|10377,10379
complete|10380,10388
an|10389,10391
8|10392,10393
week|10394,10398
course|10399,10405
of|10406,10408
high|10409,10413
dose|10414,10418
<EOL>|10419,10420
PPI|10420,10423
(|10424,10425
started|10425,10432
40mg|10433,10437
pantoprazole|10438,10450
PO|10451,10453
twice|10454,10459
daily|10460,10465
on|10466,10468
_|10469,10470
_|10470,10471
_|10471,10472
with|10473,10477
<EOL>|10478,10479
projected|10479,10488
end|10489,10492
date|10493,10497
_|10498,10499
_|10499,10500
_|10500,10501
for|10502,10505
upper|10506,10511
GI|10512,10514
bleed|10515,10520
likely|10521,10527
from|10528,10532
<EOL>|10533,10534
gastritis|10534,10543
.|10543,10544
<EOL>|10544,10545
-|10545,10546
Patient|10547,10554
's|10554,10556
hypertension|10557,10569
medications|10570,10581
(|10582,10583
Lisinopril|10583,10593
and|10594,10597
nifedipine|10598,10608
)|10608,10609
<EOL>|10610,10611
were|10611,10615
held|10616,10620
due|10621,10624
to|10625,10627
upper|10628,10633
GI|10634,10636
bleed|10637,10642
.|10642,10643
<EOL>|10643,10644
-|10644,10645
Patient|10646,10653
's|10653,10655
furosemide|10656,10666
was|10667,10670
decreased|10671,10680
to|10681,10683
20mg|10684,10688
daily|10689,10694
<EOL>|10694,10695
-|10695,10696
Patient|10697,10704
's|10704,10706
nifedipine|10707,10717
was|10718,10721
decreased|10722,10731
to|10732,10734
30mg|10735,10739
daily|10740,10745
given|10746,10751
acute|10752,10757
<EOL>|10758,10759
bleed|10759,10764
and|10765,10768
SBPs|10769,10773
in|10774,10776
the|10777,10780
_|10781,10782
_|10782,10783
_|10783,10784
<EOL>|10784,10785
-|10785,10786
Patient|10787,10794
was|10795,10798
started|10799,10806
on|10807,10809
Coumadin|10810,10818
.|10818,10819
Clopidogrel|10820,10831
was|10832,10835
stopped|10836,10843
per|10844,10847
<EOL>|10848,10849
cardiology|10849,10859
.|10859,10860
ASA|10861,10864
81mg|10865,10869
was|10870,10873
continued|10874,10883
.|10883,10884
<EOL>|10884,10885
-|10885,10886
Please|10887,10893
address|10894,10901
patient|10902,10909
's|10909,10911
home|10912,10916
environment|10917,10928
for|10929,10932
fall|10933,10937
risk|10938,10942
given|10943,10948
<EOL>|10949,10950
recent|10950,10956
"|10957,10958
trip|10958,10962
"|10962,10963
at|10964,10966
home|10967,10971
and|10972,10975
new|10976,10979
anticoagulation|10980,10995
.|10995,10996
<EOL>|10996,10997
-|10997,10998
please|10999,11005
ensure|11006,11012
patient|11013,11020
has|11021,11024
outpatient|11025,11035
anticoagulation|11036,11051
follow|11052,11058
-|11058,11059
up|11059,11061
<EOL>|11062,11063
and|11063,11066
management|11067,11077
upon|11078,11082
discharge|11083,11092
from|11093,11097
rehab|11098,11103
<EOL>|11103,11104
<EOL>|11105,11106
<EOL>|11106,11107
<EOL>|11108,11109
Medications|11109,11120
on|11121,11123
Admission|11124,11133
:|11133,11134
<EOL>|11134,11135
The|11135,11138
Preadmission|11139,11151
Medication|11152,11162
list|11163,11167
is|11168,11170
accurate|11171,11179
and|11180,11183
complete|11184,11192
.|11192,11193
<EOL>|11193,11194
1.|11194,11196
Lisinopril|11197,11207
40|11208,11210
mg|11211,11213
PO|11214,11216
DAILY|11217,11222
<EOL>|11223,11224
2.|11224,11226
Allopurinol|11227,11238
_|11239,11240
_|11240,11241
_|11241,11242
mg|11243,11245
PO|11246,11248
DAILY|11249,11254
<EOL>|11255,11256
3.|11256,11258
Atorvastatin|11259,11271
80|11272,11274
mg|11275,11277
PO|11278,11280
QPM|11281,11284
<EOL>|11285,11286
4.|11286,11288
Carvedilol|11289,11299
12.5|11300,11304
mg|11305,11307
PO|11308,11310
BID|11311,11314
<EOL>|11315,11316
5.|11316,11318
Clopidogrel|11319,11330
75|11331,11333
mg|11334,11336
PO|11337,11339
DAILY|11340,11345
<EOL>|11346,11347
6.|11347,11349
Furosemide|11350,11360
40|11361,11363
mg|11364,11366
PO|11367,11369
DAILY|11370,11375
<EOL>|11376,11377
7.|11377,11379
Ranitidine|11380,11390
150|11391,11394
mg|11395,11397
PO|11398,11400
DAILY|11401,11406
:|11406,11407
PRN|11407,11410
reflux|11411,11417
<EOL>|11418,11419
8.|11419,11421
Aspirin|11422,11429
81|11430,11432
mg|11433,11435
PO|11436,11438
DAILY|11439,11444
<EOL>|11445,11446
9.|11446,11448
Multivitamins|11449,11462
1|11463,11464
TAB|11465,11468
PO|11469,11471
DAILY|11472,11477
<EOL>|11478,11479
10|11479,11481
.|11481,11482
Vitamin|11483,11490
D|11491,11492
_|11493,11494
_|11494,11495
_|11495,11496
UNIT|11497,11501
PO|11502,11504
DAILY|11505,11510
<EOL>|11511,11512
11.|11512,11515
NIFEdipine|11516,11526
CR|11527,11529
60|11530,11532
mg|11533,11535
PO|11536,11538
BID|11539,11542
<EOL>|11543,11544
12.|11544,11547
Nitroglycerin|11548,11561
SL|11562,11564
0.3|11565,11568
mg|11569,11571
SL|11572,11574
Q5MIN|11575,11580
:|11580,11581
PRN|11581,11584
chest|11585,11590
pain|11591,11595
<EOL>|11596,11597
13.|11597,11600
70|11601,11603
/|11603,11604
30|11604,11606
30|11607,11609
Units|11610,11615
Dinner|11616,11622
<EOL>|11622,11623
<EOL>|11623,11624
<EOL>|11625,11626
Discharge|11626,11635
Medications|11636,11647
:|11647,11648
<EOL>|11648,11649
1.|11649,11651
Allopurinol|11652,11663
_|11664,11665
_|11665,11666
_|11666,11667
mg|11668,11670
PO|11671,11673
EVERY|11674,11679
OTHER|11680,11685
DAY|11686,11689
<EOL>|11690,11691
2.|11691,11693
Aspirin|11694,11701
81|11702,11704
mg|11705,11707
PO|11708,11710
DAILY|11711,11716
<EOL>|11717,11718
3.|11718,11720
Atorvastatin|11721,11733
80|11734,11736
mg|11737,11739
PO|11740,11742
QPM|11743,11746
<EOL>|11747,11748
4.|11748,11750
Carvedilol|11751,11761
12.5|11762,11766
mg|11767,11769
PO|11770,11772
BID|11773,11776
<EOL>|11777,11778
5.|11778,11780
70|11781,11783
/|11783,11784
30|11784,11786
30|11787,11789
Units|11790,11795
Dinner|11796,11802
<EOL>|11802,11803
6.|11803,11805
Lisinopril|11806,11816
40|11817,11819
mg|11820,11822
PO|11823,11825
DAILY|11826,11831
<EOL>|11832,11833
7.|11833,11835
Multivitamins|11836,11849
1|11850,11851
TAB|11852,11855
PO|11856,11858
DAILY|11859,11864
<EOL>|11865,11866
8.|11866,11868
NIFEdipine|11869,11879
CR|11880,11882
30|11883,11885
mg|11886,11888
PO|11889,11891
BID|11892,11895
<EOL>|11896,11897
9.|11897,11899
Vitamin|11900,11907
D|11908,11909
_|11910,11911
_|11911,11912
_|11912,11913
UNIT|11914,11918
PO|11919,11921
DAILY|11922,11927
<EOL>|11928,11929
10.|11929,11932
Docusate|11933,11941
Sodium|11942,11948
100|11949,11952
mg|11953,11955
PO|11956,11958
BID|11959,11962
<EOL>|11963,11964
11.|11964,11967
Gabapentin|11968,11978
100|11979,11982
mg|11983,11985
PO|11986,11988
QHS|11989,11992
neuropathic|11993,12004
pain|12005,12009
<EOL>|12010,12011
12.|12011,12014
Pantoprazole|12015,12027
40|12028,12030
mg|12031,12033
PO|12034,12036
Q12H|12037,12041
<EOL>|12042,12043
13.|12043,12046
Senna|12047,12052
8.6|12053,12056
mg|12057,12059
PO|12060,12062
BID|12063,12066
constipation|12067,12079
<EOL>|12080,12081
14.|12081,12084
Warfarin|12085,12093
5|12094,12095
mg|12096,12098
PO|12099,12101
DAILY16|12102,12109
<EOL>|12110,12111
please|12111,12117
dose|12118,12122
and|12123,12126
adjust|12127,12133
for|12134,12137
INR|12138,12141
<EOL>|12142,12143
15|12143,12145
.|12145,12146
Nitroglycerin|12147,12160
SL|12161,12163
0.3|12164,12167
mg|12168,12170
SL|12171,12173
Q5MIN|12174,12179
:|12179,12180
PRN|12180,12183
chest|12184,12189
pain|12190,12194
<EOL>|12195,12196
16|12196,12198
.|12198,12199
Furosemide|12200,12210
20|12211,12213
mg|12214,12216
PO|12217,12219
DAILY|12220,12225
<EOL>|12226,12227
17.|12227,12230
Polyethylene|12231,12243
Glycol|12244,12250
17|12251,12253
g|12254,12255
PO|12256,12258
DAILY|12259,12264
<EOL>|12265,12266
18.|12266,12269
Acetaminophen|12270,12283
325|12284,12287
-|12287,12288
650|12288,12291
mg|12292,12294
PO|12295,12297
Q6H|12298,12301
:|12301,12302
PRN|12302,12305
pain|12306,12310
or|12311,12313
fever|12314,12319
<EOL>|12320,12321
<EOL>|12321,12322
<EOL>|12323,12324
Discharge|12324,12333
Disposition|12334,12345
:|12345,12346
<EOL>|12346,12347
Extended|12347,12355
Care|12356,12360
<EOL>|12360,12361
<EOL>|12362,12363
Facility|12363,12371
:|12371,12372
<EOL>|12372,12373
_|12373,12374
_|12374,12375
_|12375,12376
<EOL>|12376,12377
<EOL>|12378,12379
Discharge|12379,12388
Diagnosis|12389,12398
:|12398,12399
<EOL>|12399,12400
Primary|12400,12407
:|12407,12408
<EOL>|12408,12409
Deep|12409,12413
vein|12414,12418
thrombosis|12419,12429
(|12430,12431
DVT|12431,12434
)|12434,12435
<EOL>|12435,12436
<EOL>|12436,12437
Secondary|12437,12446
:|12446,12447
<EOL>|12447,12448
Upper|12448,12453
GI|12454,12456
bleed|12457,12462
<EOL>|12462,12463
L|12463,12464
arm|12465,12468
hematoma|12469,12477
<EOL>|12477,12478
Superficial|12478,12489
thrombophlebitis|12490,12506
,|12506,12507
L|12508,12509
antecubital|12510,12521
fossa|12522,12527
<EOL>|12527,12528
Chronic|12528,12535
kidney|12536,12542
disease|12543,12550
(|12551,12552
Stage|12552,12557
IV|12558,12560
)|12560,12561
<EOL>|12561,12562
Peripheral|12562,12572
vascular|12573,12581
disease|12582,12589
<EOL>|12589,12590
Diabetes|12590,12598
mellitus|12599,12607
type|12608,12612
II|12613,12615
<EOL>|12615,12616
Coronary|12616,12624
artery|12625,12631
disease|12632,12639
<EOL>|12639,12640
<EOL>|12640,12641
<EOL>|12642,12643
Discharge|12643,12652
Condition|12653,12662
:|12662,12663
<EOL>|12663,12664
Mental|12664,12670
Status|12671,12677
:|12677,12678
Clear|12679,12684
and|12685,12688
coherent|12689,12697
.|12697,12698
<EOL>|12698,12699
Level|12699,12704
of|12705,12707
Consciousness|12708,12721
:|12721,12722
Alert|12723,12728
and|12729,12732
interactive|12733,12744
.|12744,12745
<EOL>|12745,12746
<EOL>|12746,12747
<EOL>|12748,12749
Discharge|12749,12758
Instructions|12759,12771
:|12771,12772
<EOL>|12772,12773
Dear|12773,12777
_|12778,12779
_|12779,12780
_|12780,12781
,|12781,12782
<EOL>|12782,12783
<EOL>|12783,12784
It|12784,12786
was|12787,12790
a|12791,12792
pleasure|12793,12801
caring|12802,12808
for|12809,12812
you|12813,12816
at|12817,12819
_|12820,12821
_|12821,12822
_|12822,12823
.|12823,12824
You|12825,12828
were|12829,12833
admitted|12834,12842
for|12843,12846
<EOL>|12847,12848
leg|12848,12851
swelling|12852,12860
and|12861,12864
pain|12865,12869
.|12869,12870
Diagnostic|12871,12881
tests|12882,12887
were|12888,12892
performed|12893,12902
and|12903,12906
you|12907,12910
<EOL>|12911,12912
were|12912,12916
diagnosed|12917,12926
with|12927,12931
deep|12932,12936
vein|12937,12941
thrombosis|12942,12952
,|12952,12953
blood|12954,12959
clots|12960,12965
in|12966,12968
your|12969,12973
<EOL>|12974,12975
legs|12975,12979
.|12979,12980
You|12981,12984
were|12985,12989
treated|12990,12997
with|12998,13002
blood|13003,13008
thinning|13009,13017
medications|13018,13029
that|13030,13034
you|13035,13038
<EOL>|13039,13040
will|13040,13044
continue|13045,13053
at|13054,13056
home|13057,13061
.|13061,13062
You|13063,13066
had|13067,13070
an|13071,13073
episode|13074,13081
of|13082,13084
upper|13085,13090
GI|13091,13093
bleeding|13094,13102
<EOL>|13103,13104
during|13104,13110
your|13111,13115
stay|13116,13120
for|13121,13124
which|13125,13130
you|13131,13134
are|13135,13138
being|13139,13144
treated|13145,13152
with|13153,13157
medication|13158,13168
<EOL>|13169,13170
and|13170,13173
you|13174,13177
underwent|13178,13187
an|13188,13190
EGD|13191,13194
.|13194,13195
You|13196,13199
developed|13200,13209
a|13210,13211
left|13212,13216
arm|13217,13220
hematoma|13221,13229
as|13230,13232
<EOL>|13233,13234
well|13234,13238
during|13239,13245
your|13246,13250
stay|13251,13255
which|13256,13261
will|13262,13266
resolve|13267,13274
on|13275,13277
its|13278,13281
own|13282,13285
over|13286,13290
time|13291,13295
.|13295,13296
<EOL>|13296,13297
<EOL>|13297,13298
For|13298,13301
your|13302,13306
blood|13307,13312
clots|13313,13318
,|13318,13319
you|13320,13323
were|13324,13328
started|13329,13336
on|13337,13339
a|13340,13341
new|13342,13345
drug|13346,13350
called|13351,13357
<EOL>|13358,13359
warfarin|13359,13367
.|13367,13368
You|13369,13372
will|13373,13377
need|13378,13382
to|13383,13385
have|13386,13390
your|13391,13395
blood|13396,13401
checked|13402,13409
to|13410,13412
adjust|13413,13419
the|13420,13423
<EOL>|13424,13425
dosing|13425,13431
.|13431,13432
For|13433,13436
your|13437,13441
upper|13442,13447
GI|13448,13450
bleed|13451,13456
,|13456,13457
you|13458,13461
were|13462,13466
started|13467,13474
on|13475,13477
<EOL>|13478,13479
Pantoprazole|13479,13491
40mg|13492,13496
twice|13497,13502
daily|13503,13508
.|13508,13509
You|13510,13513
will|13514,13518
continue|13519,13527
this|13528,13532
drug|13533,13537
as|13538,13540
an|13541,13543
<EOL>|13544,13545
outpatient|13545,13555
for|13556,13559
at|13560,13562
least|13563,13568
8|13569,13570
weeks|13571,13576
.|13576,13577
Additionally|13578,13590
,|13590,13591
you|13592,13595
will|13596,13600
no|13601,13603
<EOL>|13604,13605
longer|13605,13611
be|13612,13614
taking|13615,13621
Clopidogrel|13622,13633
(|13634,13635
Plavix|13635,13641
)|13641,13642
,|13642,13643
until|13644,13649
you|13650,13653
speak|13654,13659
with|13660,13664
your|13665,13669
<EOL>|13670,13671
cardiologist|13671,13683
.|13683,13684
<EOL>|13684,13685
<EOL>|13685,13686
It|13686,13688
was|13689,13692
a|13693,13694
pleasure|13695,13703
taking|13704,13710
care|13711,13715
you|13716,13719
during|13720,13726
your|13727,13731
hospital|13732,13740
stay|13741,13745
.|13745,13746
<EOL>|13746,13747
<EOL>|13747,13748
Best|13748,13752
wishes|13753,13759
,|13759,13760
<EOL>|13760,13761
<EOL>|13761,13762
Your|13762,13766
_|13767,13768
_|13768,13769
_|13769,13770
Care|13771,13775
Team|13776,13780
<EOL>|13780,13781
<EOL>|13782,13783
Followup|13783,13791
Instructions|13792,13804
:|13804,13805
<EOL>|13805,13806
_|13806,13807
_|13807,13808
_|13808,13809
<EOL>|13809,13810

