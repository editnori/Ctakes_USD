 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
_|28,29
_|29,30
_|30,31
No|32,34
:|34,35
_|38,39
_|39,40
_|40,41
<EOL>|41,42
<EOL>|43,44
Admission|44,53
Date|54,58
:|58,59
_|61,62
_|62,63
_|63,64
Discharge|78,87
Date|88,92
:|92,93
_|96,97
_|97,98
_|98,99
<EOL>|99,100
<EOL>|101,102
Date|102,106
of|107,109
Birth|110,115
:|115,116
_|118,119
_|119,120
_|120,121
Sex|134,137
:|137,138
M|141,142
<EOL>|142,143
<EOL>|144,145
Service|145,152
:|152,153
NEUROSURGERY|154,166
<EOL>|166,167
<EOL>|168,169
Patient|181,188
recorded|189,197
as|198,200
having|201,207
No|208,210
Known|211,216
Allergies|217,226
to|227,229
Drugs|230,235
<EOL>|235,236
<EOL>|237,238
Attending|238,247
:|247,248
_|249,250
_|250,251
_|251,252
.|252,253
<EOL>|253,254
<EOL>|255,256
Gait|273,277
instability|278,289
,|289,290
multiple|291,299
falls|300,305
<EOL>|305,306
<EOL>|307,308
Major|308,313
Surgical|314,322
or|323,325
Invasive|326,334
Procedure|335,344
:|344,345
<EOL>|345,346
None|346,350
<EOL>|350,351
<EOL>|351,352
<EOL>|353,354
Mr|382,384
_|385,386
_|386,387
_|387,388
is|389,391
a|392,393
pleasant|394,402
right|403,408
handed|409,415
_|416,417
_|417,418
_|418,419
year|420,424
old|425,428
male|429,433
with|434,438
Afib|439,443
,|443,444
<EOL>|445,446
on|446,448
coumadin|449,457
,|457,458
who|459,462
is|463,465
quite|466,471
independent|472,483
,|483,484
living|485,491
with|492,496
his|497,500
wife|501,505
and|506,509
<EOL>|510,511
was|511,514
in|515,517
a|518,519
good|520,524
state|525,530
of|531,533
health|534,540
until|541,546
mid|547,550
last|551,555
year|556,560
.|560,561
At|562,564
that|565,569
time|570,574
<EOL>|575,576
his|576,579
wife|580,584
reports|585,592
that|593,597
he|598,600
began|601,606
having|607,613
periods|614,621
of|622,624
disorganized|625,637
<EOL>|638,639
speech|639,645
and|646,649
gait|650,654
instability|655,666
.|666,667
He|668,670
did|671,674
not|675,678
have|679,683
a|684,685
fall|686,690
until|691,696
3|697,698
<EOL>|699,700
months|700,706
ago|707,710
when|711,715
he|716,718
broke|719,724
several|725,732
ribs|733,737
on|738,740
his|741,744
coffee|745,751
table|752,757
.|757,758
He|759,761
<EOL>|762,763
did|763,766
not|767,770
have|771,775
any|776,779
head|780,784
trauma|785,791
and|792,795
was|796,799
not|800,803
scanned|804,811
at|812,814
an|815,817
OSH|818,821
.|821,822
His|823,826
<EOL>|827,828
garbled|828,835
speech|836,842
and|843,846
unsteadiness|847,859
have|860,864
waxed|865,870
and|871,874
waned|875,880
over|881,885
the|886,889
<EOL>|890,891
past|891,895
6|896,897
months|898,904
and|905,908
his|909,912
wife|913,917
reports|918,925
that|926,930
they|931,935
are|936,939
much|940,944
improved|945,953
<EOL>|954,955
when|955,959
he|960,962
takes|963,968
his|969,972
diuretics|973,982
.|982,983
Over|984,988
this|989,993
period|994,1000
he|1001,1003
has|1004,1007
lost|1008,1012
~|1013,1014
20|1014,1016
<EOL>|1017,1018
lbs|1018,1021
.|1021,1022
<EOL>|1023,1024
Last|1024,1028
night|1029,1034
he|1035,1037
was|1038,1041
sorting|1042,1049
papers|1050,1056
at|1057,1059
the|1060,1063
dining|1064,1070
room|1071,1075
table|1076,1081
when|1082,1086
<EOL>|1087,1088
he|1088,1090
fell|1091,1095
from|1096,1100
standing|1101,1109
because|1110,1117
of|1118,1120
the|1121,1124
dizziness|1125,1134
.|1134,1135
He|1136,1138
reports|1139,1146
no|1147,1149
<EOL>|1150,1151
LOC|1151,1154
,|1154,1155
no|1156,1158
head|1159,1163
trauma|1164,1170
and|1171,1174
was|1175,1178
able|1179,1183
to|1184,1186
stand|1187,1192
back|1193,1197
up|1198,1200
and|1201,1204
continue|1205,1213
<EOL>|1214,1215
his|1215,1218
work|1219,1223
.|1223,1224
His|1225,1228
wife|1229,1233
placed|1234,1240
him|1241,1244
on|1245,1247
the|1248,1251
couch|1252,1257
,|1257,1258
but|1259,1262
he|1263,1265
got|1266,1269
back|1270,1274
up|1275,1277
<EOL>|1278,1279
and|1279,1282
fell|1283,1287
in|1288,1290
the|1291,1294
bathroom|1295,1303
-|1304,1305
again|1306,1311
he|1312,1314
denies|1315,1321
any|1322,1325
LOC|1326,1329
or|1330,1332
head|1333,1337
<EOL>|1338,1339
trauma|1339,1345
,|1345,1346
blaming|1347,1354
his|1355,1358
instability|1359,1370
and|1371,1374
_|1375,1376
_|1376,1377
_|1377,1378
weakness|1379,1387
.|1387,1388
He|1389,1391
had|1392,1395
no|1396,1398
<EOL>|1399,1400
tongue|1400,1406
biting|1407,1413
or|1414,1416
loss|1417,1421
of|1422,1424
bowel|1425,1430
/|1430,1431
bladder|1431,1438
continence|1439,1449
.|1449,1450
He|1451,1453
went|1454,1458
to|1459,1461
<EOL>|1462,1463
bed|1463,1466
last|1467,1471
night|1472,1477
,|1477,1478
but|1479,1482
the|1483,1486
morning|1487,1494
of|1495,1497
presentation|1498,1510
his|1511,1514
wife|1515,1519
was|1520,1523
<EOL>|1524,1525
concerned|1525,1534
about|1535,1540
his|1541,1544
falls|1545,1550
and|1551,1554
brought|1555,1562
him|1563,1566
to|1567,1569
the|1570,1573
ED|1574,1576
.|1576,1577
He|1578,1580
does|1581,1585
<EOL>|1586,1587
have|1587,1591
a|1592,1593
diagnosis|1594,1603
of|1604,1606
DM|1607,1609
II|1610,1612
from|1613,1617
just|1618,1622
over|1623,1627
a|1628,1629
month|1630,1635
ago|1636,1639
and|1640,1643
has|1644,1647
<EOL>|1648,1649
started|1649,1656
oral|1657,1661
hypoglycemics|1662,1675
for|1676,1679
which|1680,1685
he|1686,1688
reports|1689,1696
having|1697,1703
low|1704,1707
_|1708,1709
_|1709,1710
_|1710,1711
at|1712,1714
<EOL>|1715,1716
home|1716,1720
.|1720,1721
He|1722,1724
was|1725,1728
seen|1729,1733
by|1734,1736
an|1737,1739
outside|1740,1747
neurologist|1748,1759
the|1760,1763
week|1764,1768
prior|1769,1774
who|1775,1778
<EOL>|1779,1780
had|1780,1783
ordered|1784,1791
a|1792,1793
CT|1794,1796
head|1797,1801
to|1802,1804
be|1805,1807
completed|1808,1817
the|1818,1821
following|1822,1831
week|1832,1836
.|1836,1837
In|1838,1840
the|1841,1844
<EOL>|1845,1846
ED|1846,1848
his|1849,1852
head|1853,1857
was|1858,1861
scanned|1862,1869
which|1870,1875
revealed|1876,1884
no|1885,1887
bleed|1888,1893
but|1894,1897
a|1898,1899
3x3|1900,1903
L|1904,1905
<EOL>|1906,1907
frontal|1907,1914
lobe|1915,1919
extra-axial|1920,1931
mass|1932,1936
with|1937,1941
compressive|1942,1953
effect|1954,1960
but|1961,1964
<EOL>|1964,1965
no|1965,1967
midline|1968,1975
shift|1976,1981
.|1981,1982
Neurosurgery|1983,1995
was|1996,1999
contacted|2000,2009
for|2010,2013
evaluation|2014,2024
of|2025,2027
<EOL>|2028,2029
the|2029,2032
mass|2033,2037
and|2038,2041
its|2042,2045
possible|2046,2054
role|2055,2059
in|2060,2062
the|2063,2066
patient|2067,2074
's|2074,2076
recent|2077,2083
symptoms|2084,2092
.|2092,2093
<EOL>|2094,2095
<EOL>|2095,2096
<EOL>|2097,2098
DM|2120,2122
II|2123,2125
,|2125,2126
HTN|2127,2130
,|2130,2131
HL|2132,2134
,|2134,2135
MI|2136,2138
(|2139,2140
in|2140,2142
past|2143,2147
)|2147,2148
,|2148,2149
AF|2150,2152
on|2153,2155
coumadin|2156,2164
,|2164,2165
prostate|2166,2174
CA|2175,2177
<EOL>|2178,2179
treated|2179,2186
non-operatively|2187,2202
<EOL>|2202,2203
<EOL>|2203,2204
<EOL>|2205,2206
:|2220,2221
<EOL>|2221,2222
_|2222,2223
_|2223,2224
_|2224,2225
<EOL>|2225,2226
:|2240,2241
<EOL>|2241,2242
Non-contributory|2242,2258
<EOL>|2259,2260
<EOL>|2261,2262
At|2277,2279
Admission|2280,2289
:|2289,2290
<EOL>|2291,2292
<EOL>|2292,2293
Gen|2293,2296
:|2296,2297
WD|2298,2300
/|2300,2301
WN|2301,2303
,|2303,2304
comfortable|2305,2316
,|2316,2317
NAD|2318,2321
.|2321,2322
<EOL>|2322,2323
HEENT|2323,2328
:|2328,2329
Pupils|2330,2336
:|2336,2337
4|2338,2339
-|2339,2340
>|2340,2341
3|2341,2342
EOMs|2346,2350
intact|2351,2357
b|2358,2359
/|2359,2360
l|2360,2361
<EOL>|2361,2362
Lungs|2362,2367
:|2367,2368
CTA|2369,2372
bilaterally|2373,2384
.|2384,2385
<EOL>|2385,2386
Cardiac|2386,2393
:|2393,2394
irreg|2395,2400
irreg|2401,2406
with|2407,2411
_|2412,2413
_|2413,2414
_|2414,2415
holosystolic|2416,2428
murmur|2429,2435
.|2435,2436
<EOL>|2436,2437
Abd|2437,2440
:|2440,2441
Soft|2442,2446
,|2446,2447
NT|2448,2450
,|2450,2451
BS|2452,2454
+|2454,2455
<EOL>|2455,2456
Extrem|2456,2462
:|2462,2463
Warm|2464,2468
and|2469,2472
well|2473,2477
-|2477,2478
perfused|2478,2486
.|2486,2487
<EOL>|2487,2488
Neuro|2488,2493
:|2493,2494
<EOL>|2494,2495
Mental|2495,2501
status|2502,2508
:|2508,2509
Awake|2510,2515
and|2516,2519
cooperative|2520,2531
with|2532,2536
exam|2537,2541
,|2541,2542
normal|2543,2549
affect|2550,2556
.|2556,2557
<EOL>|2557,2558
Orientation|2558,2569
:|2569,2570
Oriented|2571,2579
to|2580,2582
person|2583,2589
,|2589,2590
place|2591,2596
,|2596,2597
and|2598,2601
date|2602,2606
.|2606,2607
<EOL>|2607,2608
Recall|2608,2614
:|2614,2615
_|2616,2617
_|2617,2618
_|2618,2619
objects|2620,2627
at|2628,2630
5|2631,2632
minutes|2633,2640
.|2640,2641
<EOL>|2641,2642
Language|2642,2650
:|2650,2651
Speech|2652,2658
is|2659,2661
fluent|2662,2668
,|2668,2669
good|2670,2674
comprehension|2675,2688
.|2688,2689
Difficulty|2690,2700
with|2701,2705
<EOL>|2705,2706
repitition|2706,2716
.|2716,2717
Naming|2718,2724
intact|2725,2731
.|2731,2732
No|2733,2735
dysarthria|2736,2746
or|2747,2749
paraphasic|2750,2760
errors|2761,2767
.|2767,2768
<EOL>|2768,2769
<EOL>|2769,2770
Cranial|2770,2777
Nerves|2778,2784
:|2784,2785
<EOL>|2785,2786
I|2786,2787
:|2787,2788
Not|2789,2792
tested|2793,2799
<EOL>|2799,2800
II|2800,2802
:|2802,2803
Pupils|2804,2810
equally|2811,2818
round|2819,2824
and|2825,2828
reactive|2829,2837
to|2838,2840
light|2841,2846
,|2846,2847
to|2848,2850
<EOL>|2850,2851
mm|2851,2853
bilaterally|2854,2865
.|2865,2866
Visual|2867,2873
fields|2874,2880
are|2881,2884
full|2885,2889
to|2890,2892
confrontation|2893,2906
.|2906,2907
<EOL>|2907,2908
III|2908,2911
,|2911,2912
IV|2913,2915
,|2915,2916
VI|2917,2919
:|2919,2920
Extraocular|2921,2932
movements|2933,2942
intact|2943,2949
bilaterally|2950,2961
without|2962,2969
<EOL>|2969,2970
nystagmus|2970,2979
.|2979,2980
<EOL>|2980,2981
V|2981,2982
,|2982,2983
VII|2984,2987
:|2987,2988
Facial|2989,2995
strength|2996,3004
and|3005,3008
sensation|3009,3018
intact|3019,3025
and|3026,3029
symmetric|3030,3039
.|3039,3040
<EOL>|3040,3041
VIII|3041,3045
:|3045,3046
Hearing|3047,3054
intact|3055,3061
to|3062,3064
voice|3065,3070
.|3070,3071
<EOL>|3071,3072
IX|3072,3074
,|3074,3075
X|3076,3077
:|3077,3078
Palatal|3079,3086
elevation|3087,3096
symmetrical|3097,3108
.|3108,3109
<EOL>|3109,3110
XI|3110,3112
:|3112,3113
Sternocleidomastoid|3114,3133
and|3134,3137
trapezius|3138,3147
normal|3148,3154
bilaterally|3155,3166
.|3166,3167
<EOL>|3167,3168
XII|3168,3171
:|3171,3172
Tongue|3173,3179
midline|3180,3187
without|3188,3195
fasciculations|3196,3210
.|3210,3211
<EOL>|3211,3212
<EOL>|3212,3213
Motor|3213,3218
:|3218,3219
Normal|3220,3226
bulk|3227,3231
and|3232,3235
tone|3236,3240
bilaterally|3241,3252
.|3252,3253
No|3254,3256
abnormal|3257,3265
movements|3266,3275
,|3275,3276
<EOL>|3276,3277
tremors|3277,3284
.|3284,3285
Strength|3286,3294
full|3295,3299
power|3300,3305
_|3306,3307
_|3307,3308
_|3308,3309
throughout|3310,3320
.|3320,3321
Mild|3322,3326
R|3327,3328
sided|3329,3334
<EOL>|3334,3335
pronator|3335,3343
drift|3344,3349
.|3349,3350
Gait|3351,3355
unsteady|3356,3364
,|3364,3365
rhomberg|3366,3374
test|3375,3379
with|3380,3384
unsteadiness|3385,3397
.|3397,3398
<EOL>|3398,3399
<EOL>|3399,3400
Sensation|3400,3409
:|3409,3410
Intact|3411,3417
to|3418,3420
light|3421,3426
touch|3427,3432
,|3432,3433
propioception|3434,3447
,|3447,3448
pinprick|3449,3457
and|3458,3461
<EOL>|3461,3462
vibration|3462,3471
bilaterally|3472,3483
.|3483,3484
<EOL>|3484,3485
<EOL>|3485,3486
Reflexes|3486,3494
:|3494,3495
B|3496,3497
T|3498,3499
Br|3500,3502
Pa|3503,3505
Ac|3506,3508
<EOL>|3508,3509
Right|3509,3514
_|3519,3520
_|3520,3521
_|3521,3522
1|3523,3524
1|3526,3527
<EOL>|3527,3528
Left|3528,3532
_|3538,3539
_|3539,3540
_|3540,3541
1|3542,3543
1|3545,3546
<EOL>|3546,3547
<EOL>|3547,3548
Toes|3548,3552
downgoing|3553,3562
bilaterally|3563,3574
<EOL>|3574,3575
<EOL>|3575,3576
Coordination|3576,3588
:|3588,3589
heel|3590,3594
to|3595,3597
shin|3598,3602
intact|3603,3609
,|3609,3610
finger|3611,3617
nose|3618,3622
-|3622,3623
finger|3623,3629
slowed|3630,3636
and|3637,3640
<EOL>|3640,3641
overshooting|3641,3653
with|3654,3658
R|3659,3660
hand|3661,3665
.|3665,3666
Difficulty|3667,3677
with|3678,3682
rapid|3683,3688
alternating|3689,3700
<EOL>|3700,3701
movements|3701,3710
with|3711,3715
R|3716,3717
hand|3718,3722
.|3722,3723
<EOL>|3723,3724
<EOL>|3724,3725
AT|3725,3727
DISCHARGE|3728,3737
:|3737,3738
<EOL>|3739,3740
Afeb|3740,3744
,|3744,3745
VSS|3746,3749
<EOL>|3749,3750
Gen|3750,3753
:|3753,3754
NAD|3755,3758
.|3758,3759
<EOL>|3759,3760
HEENT|3760,3765
:|3765,3766
Pupils|3767,3773
:|3773,3774
3|3775,3776
-|3776,3777
>|3777,3778
2|3778,3779
EOMs|3781,3785
intact|3786,3792
b|3793,3794
/|3794,3795
l|3795,3796
<EOL>|3796,3797
Lungs|3797,3802
:|3802,3803
clear|3804,3809
b|3810,3811
/|3811,3812
l|3812,3813
<EOL>|3813,3814
Cardiac|3814,3821
:|3821,3822
irreg|3823,3828
irreg|3829,3834
with|3835,3839
_|3840,3841
_|3841,3842
_|3842,3843
holosystolic|3844,3856
murmur|3857,3863
.|3863,3864
<EOL>|3864,3865
Abd|3865,3868
:|3868,3869
non-tender|3870,3880
/|3880,3881
non-distended|3881,3894
<EOL>|3894,3895
Extrem|3895,3901
:|3901,3902
no|3903,3905
edema|3906,3911
or|3912,3914
erythema|3915,3923
,|3923,3924
warm|3925,3929
well|3930,3934
perfused|3935,3943
.|3943,3944
<EOL>|3944,3945
<EOL>|3945,3946
Neuro|3946,3951
:|3951,3952
<EOL>|3952,3953
Mental|3953,3959
status|3960,3966
:|3966,3967
Awake|3968,3973
and|3974,3977
cooperative|3978,3989
with|3990,3994
exam|3995,3999
,|3999,4000
normal|4001,4007
affect|4008,4014
.|4014,4015
<EOL>|4015,4016
Orientation|4016,4027
:|4027,4028
Oriented|4029,4037
to|4038,4040
person|4041,4047
,|4047,4048
place|4049,4054
,|4054,4055
and|4056,4059
date|4060,4064
.|4064,4065
<EOL>|4065,4066
Language|4066,4074
:|4074,4075
Speech|4076,4082
is|4083,4085
fluent|4086,4092
,|4092,4093
good|4094,4098
comprehension|4099,4112
.|4112,4113
<EOL>|4113,4114
<EOL>|4114,4115
Cranial|4115,4122
Nerves|4123,4129
:|4129,4130
<EOL>|4130,4131
II|4131,4133
-|4133,4134
XII|4134,4137
tested|4138,4144
and|4145,4148
intact|4149,4155
b|4156,4157
/|4157,4158
l|4158,4159
<EOL>|4159,4160
<EOL>|4160,4161
Motor|4161,4166
:|4166,4167
_|4168,4169
_|4169,4170
_|4170,4171
strength|4172,4180
b|4181,4182
/|4182,4183
l|4183,4184
in|4185,4187
UE|4188,4190
and|4191,4194
_|4195,4196
_|4196,4197
_|4197,4198
.|4198,4199
No|4200,4202
pronator|4203,4211
drift|4212,4217
.|4217,4218
Gait|4219,4223
<EOL>|4224,4225
steady|4225,4231
,|4231,4232
walking|4233,4240
without|4241,4248
assistance|4249,4259
.|4259,4260
<EOL>|4260,4261
<EOL>|4261,4262
Sensation|4262,4271
:|4271,4272
Grossly|4273,4280
intact|4281,4287
b|4288,4289
/|4289,4290
l|4290,4291
.|4291,4292
<EOL>|4292,4293
<EOL>|4293,4294
Reflexes|4294,4302
:|4302,4303
B|4304,4305
T|4306,4307
Br|4308,4310
Pa|4311,4313
Ac|4314,4316
<EOL>|4316,4317
Right|4317,4322
_|4327,4328
_|4328,4329
_|4329,4330
1|4331,4332
1|4334,4335
<EOL>|4335,4336
Left|4336,4340
_|4346,4347
_|4347,4348
_|4348,4349
1|4350,4351
1|4353,4354
<EOL>|4354,4355
<EOL>|4355,4356
Toes|4356,4360
downgoing|4361,4370
bilaterally|4371,4382
<EOL>|4382,4383
<EOL>|4384,4385
Pertinent|4385,4394
Results|4395,4402
:|4402,4403
<EOL>|4403,4404
_|4404,4405
_|4405,4406
_|4406,4407
04|4408,4410
:|4410,4411
55AM|4411,4415
BLOOD|4416,4421
WBC|4422,4425
-|4425,4426
3|4426,4427
.|4427,4428
9|4428,4429
*|4429,4430
RBC|4431,4434
-|4434,4435
4|4435,4436
.|4436,4437
39|4437,4439
*|4439,4440
Hgb|4441,4444
-|4444,4445
13|4445,4447
.|4447,4448
5|4448,4449
*|4449,4450
Hct|4451,4454
-|4454,4455
40.7|4455,4459
<EOL>|4460,4461
MCV|4461,4464
-|4464,4465
93|4465,4467
MCH|4468,4471
-|4471,4472
30.7|4472,4476
MCHC|4477,4481
-|4481,4482
33.1|4482,4486
RDW|4487,4490
-|4490,4491
15.5|4491,4495
Plt|4496,4499
_|4500,4501
_|4501,4502
_|4502,4503
<EOL>|4503,4504
_|4504,4505
_|4505,4506
_|4506,4507
04|4508,4510
:|4510,4511
55AM|4511,4515
BLOOD|4516,4521
_|4522,4523
_|4523,4524
_|4524,4525
<EOL>|4525,4526
_|4526,4527
_|4527,4528
_|4528,4529
04|4530,4532
:|4532,4533
55AM|4533,4537
BLOOD|4538,4543
Glucose|4544,4551
-|4551,4552
115|4552,4555
*|4555,4556
UreaN|4557,4562
-|4562,4563
33|4563,4565
*|4565,4566
Creat|4567,4572
-|4572,4573
1.2|4573,4576
Na|4577,4579
-|4579,4580
142|4580,4583
<EOL>|4584,4585
K|4585,4586
-|4586,4587
3.7|4587,4590
Cl|4591,4593
-|4593,4594
104|4594,4597
HCO3|4598,4602
-|4602,4603
33|4603,4605
*|4605,4606
AnGap|4607,4612
-|4612,4613
9|4613,4614
<EOL>|4614,4615
_|4615,4616
_|4616,4617
_|4617,4618
06|4619,4621
:|4621,4622
25AM|4622,4626
BLOOD|4627,4632
Albumin|4633,4640
-|4640,4641
3|4641,4642
.|4642,4643
2|4643,4644
*|4644,4645
<EOL>|4645,4646
_|4646,4647
_|4647,4648
_|4648,4649
02|4650,4652
:|4652,4653
39PM|4653,4657
BLOOD|4658,4663
%|4664,4665
HbA1c|4665,4670
-|4670,4671
7|4671,4672
.|4672,4673
7|4673,4674
*|4674,4675
eAG|4676,4679
-|4679,4680
174|4680,4683
*|4683,4684
<EOL>|4684,4685
_|4685,4686
_|4686,4687
_|4687,4688
06|4689,4691
:|4691,4692
25AM|4692,4696
BLOOD|4697,4702
Phenyto|4703,4710
-|4710,4711
4|4711,4712
.|4712,4713
6|4713,4714
*|4714,4715
<EOL>|4715,4716
<EOL>|4716,4717
CT|4717,4719
Head|4720,4724
_|4725,4726
_|4726,4727
_|4727,4728
:|4728,4729
<EOL>|4730,4731
1.|4744,4746
Extra-axial|4747,4758
lesion|4759,4765
,|4765,4766
containing|4767,4777
foci|4778,4782
of|4783,4785
calcifications|4786,4800
<EOL>|4801,4802
measuring|4802,4811
up|4812,4814
to|4815,4817
3|4818,4819
cm|4820,4822
,|4822,4823
which|4824,4829
likely|4830,4836
reflects|4837,4845
an|4846,4848
extra-axial|4849,4860
mass|4861,4865
<EOL>|4866,4867
such|4867,4871
as|4872,4874
a|4875,4876
meningioma|4877,4887
.|4887,4888
An|4889,4891
<EOL>|4892,4893
extra-axial|4893,4904
hematoma|4905,4913
,|4913,4914
which|4915,4920
would|4921,4926
be|4927,4929
subacute|4930,4938
to|4939,4941
chronic|4942,4949
,|4949,4950
is|4951,4953
<EOL>|4954,4955
considered|4955,4965
less|4966,4970
likely|4971,4977
.|4977,4978
<EOL>|4979,4980
2.|4980,4982
Loss|4983,4987
of|4988,4990
gray|4991,4995
-|4995,4996
white|4996,5001
differentiation|5002,5017
in|5018,5020
the|5021,5024
high|5025,5029
left|5030,5034
<EOL>|5035,5036
frontoparietal|5036,5050
lobe|5051,5055
,|5055,5056
could|5057,5062
reflect|5063,5070
an|5071,5073
acute|5074,5079
infarct|5080,5087
.|5087,5088
<EOL>|5089,5090
<EOL>|5090,5091
MRI|5091,5094
Head|5095,5099
_|5100,5101
_|5101,5102
_|5102,5103
:|5103,5104
<EOL>|5104,5105
Acute|5105,5110
to|5111,5113
subacute|5114,5122
bilateral|5123,5132
infarctions|5133,5144
with|5145,5149
the|5150,5153
largest|5154,5161
focus|5162,5167
<EOL>|5168,5169
in|5169,5171
the|5172,5175
left|5176,5180
post-central|5181,5193
gyrus|5194,5199
.|5199,5200
Appearance|5201,5211
of|5212,5214
the|5215,5218
post-gyrus|5219,5229
<EOL>|5230,5231
lesion|5231,5237
is|5238,5240
somewhat|5241,5249
<EOL>|5250,5251
heterogeneous|5251,5264
however|5265,5272
and|5273,5276
recommend|5277,5286
attention|5287,5296
on|5297,5299
followup|5300,5308
<EOL>|5309,5310
imaging|5310,5317
for|5318,5321
further|5322,5329
evaluation|5330,5340
to|5341,5343
exclude|5344,5351
the|5352,5355
presence|5356,5364
of|5365,5367
an|5368,5370
<EOL>|5371,5372
underlying|5372,5382
mass|5383,5387
.|5387,5388
Two|5389,5392
meningiomas|5393,5404
in|5405,5407
the|5408,5411
left|5412,5416
frontal|5417,5424
region|5425,5431
<EOL>|5432,5433
without|5433,5440
significant|5441,5452
mass|5453,5457
effect|5458,5464
.|5464,5465
<EOL>|5465,5466
<EOL>|5466,5467
ECHO|5467,5471
_|5472,5473
_|5473,5474
_|5474,5475
:|5475,5476
<EOL>|5476,5477
Marked|5477,5483
symmetric|5484,5493
left|5494,5498
ventricular|5499,5510
hypertrophy|5511,5522
with|5523,5527
normal|5528,5534
cavity|5535,5541
<EOL>|5542,5543
size|5543,5547
and|5548,5551
regional|5552,5560
/|5560,5561
global|5561,5567
systolic|5568,5576
function|5577,5585
.|5585,5586
Mild|5587,5591
aortic|5592,5598
valve|5599,5604
<EOL>|5605,5606
stenosis|5606,5614
.|5614,5615
Mild|5616,5620
aortic|5621,5627
regurgitation|5628,5641
.|5641,5642
Right|5643,5648
ventricular|5649,5660
free|5661,5665
wall|5666,5670
<EOL>|5671,5672
hypertrophy|5672,5683
.|5683,5684
Pulmonary|5685,5694
artery|5695,5701
systolic|5702,5710
hypertension|5711,5723
.|5723,5724
Dilated|5725,5732
<EOL>|5733,5734
ascending|5734,5743
aorta|5744,5749
.|5749,5750
<EOL>|5751,5752
CLINICAL|5752,5760
IMPLICATIONS|5761,5773
:|5773,5774
<EOL>|5775,5776
The|5776,5779
patient|5780,5787
has|5788,5791
mild|5792,5796
aortic|5797,5803
stenosis|5804,5812
.|5812,5813
Based|5814,5819
on|5820,5822
_|5823,5824
_|5824,5825
_|5825,5826
ACC|5827,5830
/|5830,5831
AHA|5831,5834
<EOL>|5835,5836
Valvular|5836,5844
Heart|5845,5850
Disease|5851,5858
Guidelines|5859,5869
,|5869,5870
a|5871,5872
follow|5873,5879
-|5879,5880
up|5880,5882
echocardiogram|5883,5897
is|5898,5900
<EOL>|5901,5902
suggested|5902,5911
in|5912,5914
_|5915,5916
_|5916,5917
_|5917,5918
years|5919,5924
.|5924,5925
<EOL>|5926,5927
Based|5927,5932
on|5933,5935
_|5936,5937
_|5937,5938
_|5938,5939
AHA|5940,5943
endocarditis|5944,5956
prophylaxis|5957,5968
recommendations|5969,5984
,|5984,5985
the|5986,5989
<EOL>|5990,5991
echo|5991,5995
findings|5996,6004
indicate|6005,6013
prophylaxis|6014,6025
is|6026,6028
NOT|6029,6032
recommended|6033,6044
.|6044,6045
Clinical|6046,6054
<EOL>|6055,6056
decisions|6056,6065
regarding|6066,6075
the|6076,6079
need|6080,6084
for|6085,6088
prophylaxis|6089,6100
should|6101,6107
be|6108,6110
based|6111,6116
on|6117,6119
<EOL>|6120,6121
clinical|6121,6129
and|6130,6133
echocardiographic|6134,6151
data|6152,6156
.|6156,6157
<EOL>|6158,6159
<EOL>|6159,6160
MRA|6160,6163
Head|6164,6168
/|6168,6169
Neck|6169,6173
_|6174,6175
_|6175,6176
_|6176,6177
:|6177,6178
<EOL>|6178,6179
Mild|6179,6183
atherosclerotic|6184,6199
disease|6200,6207
of|6208,6210
the|6211,6214
basilar|6215,6222
artery|6223,6229
.|6229,6230
There|6231,6236
is|6237,6239
no|6240,6242
<EOL>|6243,6244
evidence|6244,6252
of|6253,6255
acute|6256,6261
vascular|6262,6270
abnormalities|6271,6284
involving|6285,6294
the|6295,6298
<EOL>|6299,6300
intracranial|6300,6312
arteries|6313,6321
<EOL>|6322,6323
<EOL>|6323,6324
<EOL>|6325,6326
<EOL>|6326,6327
<EOL>|6328,6329
Mr.|6352,6355
_|6356,6357
_|6357,6358
_|6358,6359
was|6360,6363
admitted|6364,6372
to|6373,6375
the|6376,6379
neurosurgical|6380,6393
service|6394,6401
on|6402,6404
_|6405,6406
_|6406,6407
_|6407,6408
<EOL>|6409,6410
from|6410,6414
the|6415,6418
emergency|6419,6428
room|6429,6433
after|6434,6439
having|6440,6446
a|6447,6448
series|6449,6455
of|6456,6458
falls|6459,6464
on|6465,6467
<EOL>|6468,6469
_|6469,6470
_|6470,6471
_|6471,6472
.|6472,6473
A|6474,6475
CT|6476,6478
of|6479,6481
the|6482,6485
head|6486,6490
demonstrated|6491,6503
a|6504,6505
left|6506,6510
frontal|6511,6518
<EOL>|6519,6520
extra-axial|6520,6531
mass|6532,6536
as|6537,6539
well|6540,6544
as|6545,6547
a|6548,6549
more|6550,6554
acute|6555,6560
lesion|6561,6567
in|6568,6570
the|6571,6574
parietal|6575,6583
<EOL>|6584,6585
lobe|6585,6589
on|6590,6592
the|6593,6596
left|6597,6601
.|6601,6602
Because|6603,6610
of|6611,6613
his|6614,6617
recent|6618,6624
falls|6625,6630
,|6630,6631
his|6632,6635
coumadin|6636,6644
was|6645,6648
<EOL>|6649,6650
held|6650,6654
and|6655,6658
he|6659,6661
was|6662,6665
placed|6666,6672
on|6673,6675
an|6676,6678
insulin|6679,6686
sliding|6687,6694
scale|6695,6700
as|6701,6703
there|6704,6709
was|6710,6713
<EOL>|6714,6715
some|6715,6719
concern|6720,6727
for|6728,6731
hypoglycemia|6732,6744
contributing|6745,6757
to|6758,6760
the|6761,6764
unsteadiness|6765,6777
.|6777,6778
<EOL>|6779,6780
<EOL>|6780,6781
An|6781,6783
MRI|6784,6787
of|6788,6790
this|6791,6795
head|6796,6800
was|6801,6804
obtained|6805,6813
which|6814,6819
confirmed|6820,6829
a|6830,6831
meningioma|6832,6842
<EOL>|6843,6844
overlying|6844,6853
the|6854,6857
L|6858,6859
frontal|6860,6867
lobe|6868,6872
and|6873,6876
a|6877,6878
sub-acute|6879,6888
infarct|6889,6896
in|6897,6899
the|6900,6903
<EOL>|6904,6905
post-central|6905,6917
gyrus|6918,6923
on|6924,6926
the|6927,6930
left|6931,6935
.|6935,6936
While|6937,6942
he|6943,6945
did|6946,6949
have|6950,6954
distinct|6955,6963
right|6964,6969
<EOL>|6970,6971
sided|6971,6976
weakness|6977,6985
in|6986,6988
the|6989,6992
emergency|6993,7002
room|7003,7007
,|7007,7008
on|7009,7011
hospital|7012,7020
day|7021,7024
#|7025,7026
2|7026,7027
this|7028,7032
<EOL>|7033,7034
weakness|7034,7042
had|7043,7046
nearly|7047,7053
completely|7054,7064
resolved|7065,7073
and|7074,7077
his|7078,7081
confusion|7082,7091
was|7092,7095
<EOL>|7096,7097
also|7097,7101
better|7102,7108
.|7108,7109
A|7110,7111
neurology|7112,7121
consult|7122,7129
was|7130,7133
obtained|7134,7142
given|7143,7148
what|7149,7153
<EOL>|7154,7155
appeared|7155,7163
to|7164,7166
be|7167,7169
a|7170,7171
sub-acute|7172,7181
stroke|7182,7188
on|7189,7191
his|7192,7195
MRI|7196,7199
-|7200,7201
they|7202,7206
recommended|7207,7218
<EOL>|7219,7220
restarting|7220,7230
the|7231,7234
pt|7235,7237
's|7237,7239
coumadin|7240,7248
,|7248,7249
holding|7250,7257
the|7258,7261
dilantin|7262,7270
and|7271,7274
checking|7275,7283
<EOL>|7284,7285
an|7285,7287
EEG|7288,7291
,|7291,7292
these|7293,7298
were|7299,7303
done|7304,7308
while|7309,7314
he|7315,7317
was|7318,7321
an|7322,7324
inpatient|7325,7334
.|7334,7335
He|7336,7338
also|7339,7343
<EOL>|7344,7345
underwent|7345,7354
a|7355,7356
surface|7357,7364
echo|7365,7369
and|7370,7373
an|7374,7376
MRA|7377,7380
of|7381,7383
the|7384,7387
brain|7388,7393
and|7394,7397
neck|7398,7402
given|7403,7408
<EOL>|7409,7410
the|7410,7413
likely|7414,7420
embolic|7421,7428
nature|7429,7435
of|7436,7438
his|7439,7442
strokes|7443,7450
.|7450,7451
<EOL>|7452,7453
<EOL>|7453,7454
Neurology|7454,7463
will|7464,7468
see|7469,7472
him|7473,7476
in|7477,7479
3|7480,7481
months|7482,7488
with|7489,7493
a|7494,7495
repeat|7496,7502
head|7503,7507
MRI|7508,7511
.|7511,7512
<EOL>|7513,7514
_|7514,7515
_|7515,7516
_|7516,7517
also|7518,7522
saw|7523,7526
him|7527,7530
for|7531,7534
his|7535,7538
diabetes|7539,7547
managment|7548,7557
<EOL>|7558,7559
and|7559,7562
recommended|7563,7574
changing|7575,7583
his|7584,7587
glipizide|7588,7597
to|7598,7600
10|7601,7603
BID|7604,7607
,|7607,7608
and|7609,7612
not|7613,7616
<EOL>|7617,7618
starting|7618,7626
insulin|7627,7634
.|7634,7635
His|7636,7639
sugars|7640,7646
were|7647,7651
well|7652,7656
controlled|7657,7667
while|7668,7673
in|7674,7676
house|7677,7682
<EOL>|7683,7684
and|7684,7687
he|7688,7690
did|7691,7694
not|7695,7698
have|7699,7703
any|7704,7707
episodes|7708,7716
of|7717,7719
hypoglycemia|7720,7732
.|7732,7733
From|7734,7738
a|7739,7740
<EOL>|7741,7742
neurologic|7742,7752
standpoing|7753,7763
,|7763,7764
in|7765,7767
-|7767,7768
house|7768,7773
he|7774,7776
did|7777,7780
quite|7781,7786
well|7787,7791
with|7792,7796
resultion|7797,7806
<EOL>|7807,7808
of|7808,7810
his|7811,7814
right|7815,7820
sided|7821,7826
weakness|7827,7835
although|7836,7844
his|7845,7848
unsteadiness|7849,7861
continued|7862,7871
<EOL>|7872,7873
and|7873,7876
he|7877,7879
needed|7880,7886
support|7887,7894
while|7895,7900
ambulating|7901,7911
.|7911,7912
<EOL>|7913,7914
<EOL>|7914,7915
_|7915,7916
_|7916,7917
_|7917,7918
recommended|7919,7930
he|7931,7933
go|7934,7936
to|7937,7939
a|7940,7941
short|7942,7947
term|7948,7952
rehab|7953,7958
until|7959,7964
he|7965,7967
was|7968,7971
better|7972,7978
<EOL>|7979,7980
able|7980,7984
to|7985,7987
compete|7988,7995
transfers|7996,8005
and|8006,8009
ambulate|8010,8018
with|8019,8023
a|8024,8025
walker|8026,8032
.|8032,8033
He|8034,8036
will|8037,8041
<EOL>|8042,8043
follow|8043,8049
up|8050,8052
with|8053,8057
neurology|8058,8067
and|8068,8071
neurosurgery|8072,8084
to|8085,8087
discuss|8088,8095
how|8096,8099
to|8100,8102
best|8103,8107
<EOL>|8108,8109
manage|8109,8115
his|8116,8119
ischemic|8120,8128
strokes|8129,8136
and|8137,8140
address|8141,8148
the|8149,8152
meningioma|8153,8163
,|8163,8164
<EOL>|8165,8166
respectively|8166,8178
.|8178,8179
<EOL>|8179,8180
<EOL>|8181,8182
Medications|8182,8193
on|8194,8196
Admission|8197,8206
:|8206,8207
<EOL>|8207,8208
Coumadin|8208,8216
2.5|8217,8220
'|8220,8221
,|8221,8222
prandin|8223,8230
0.5|8231,8234
'|8234,8235
'|8235,8236
'|8236,8237
,|8237,8238
glipizide|8239,8248
5|8249,8250
'|8250,8251
'|8251,8252
,|8252,8253
isosorbide|8254,8264
<EOL>|8265,8266
dinitrate|8266,8275
10|8276,8278
'|8278,8279
'|8279,8280
,|8280,8281
lisinopril|8282,8292
20|8293,8295
,|8295,8296
allopurinol|8297,8308
_|8309,8310
_|8310,8311
_|8311,8312
,|8312,8313
torsemide|8314,8323
5|8324,8325
,|8325,8326
<EOL>|8327,8328
metoprolol|8328,8338
50|8339,8341
'|8341,8342
'|8342,8343
'|8343,8344
,|8344,8345
lipitor|8346,8353
10|8354,8356
'|8356,8357
<EOL>|8357,8358
<EOL>|8358,8359
<EOL>|8360,8361
Discharge|8361,8370
Medications|8371,8382
:|8382,8383
<EOL>|8383,8384
1.|8384,8386
Isosorbide|8387,8397
Dinitrate|8398,8407
10|8408,8410
mg|8411,8413
Tablet|8414,8420
Sig|8421,8424
:|8424,8425
One|8426,8429
(|8430,8431
1|8431,8432
)|8432,8433
Tablet|8434,8440
PO|8441,8443
BID|8444,8447
<EOL>|8448,8449
(|8449,8450
2|8450,8451
times|8452,8457
a|8458,8459
day|8460,8463
)|8463,8464
.|8464,8465
<EOL>|8467,8468
2.|8468,8470
Lisinopril|8471,8481
20|8482,8484
mg|8485,8487
Tablet|8488,8494
Sig|8495,8498
:|8498,8499
One|8500,8503
(|8504,8505
1|8505,8506
)|8506,8507
Tablet|8508,8514
PO|8515,8517
DAILY|8518,8523
(|8524,8525
Daily|8525,8530
)|8530,8531
.|8531,8532
<EOL>|8533,8534
<EOL>|8535,8536
3.|8536,8538
Metoprolol|8539,8549
Tartrate|8550,8558
50|8559,8561
mg|8562,8564
Tablet|8565,8571
Sig|8572,8575
:|8575,8576
One|8577,8580
(|8581,8582
1|8582,8583
)|8583,8584
Tablet|8585,8591
PO|8592,8594
TID|8595,8598
<EOL>|8599,8600
(|8600,8601
3|8601,8602
times|8603,8608
a|8609,8610
day|8611,8614
)|8614,8615
.|8615,8616
<EOL>|8618,8619
4.|8619,8621
Simvastatin|8622,8633
10|8634,8636
mg|8637,8639
Tablet|8640,8646
Sig|8647,8650
:|8650,8651
Two|8652,8655
(|8656,8657
2|8657,8658
)|8658,8659
Tablet|8660,8666
PO|8667,8669
DAILY|8670,8675
<EOL>|8676,8677
(|8677,8678
Daily|8678,8683
)|8683,8684
.|8684,8685
<EOL>|8687,8688
5.|8688,8690
Allopurinol|8691,8702
_|8703,8704
_|8704,8705
_|8705,8706
mg|8707,8709
Tablet|8710,8716
Sig|8717,8720
:|8720,8721
One|8722,8725
(|8726,8727
1|8727,8728
)|8728,8729
Tablet|8730,8736
PO|8737,8739
DAILY|8740,8745
<EOL>|8746,8747
(|8747,8748
Daily|8748,8753
)|8753,8754
.|8754,8755
<EOL>|8757,8758
6.|8758,8760
Warfarin|8761,8769
2.5|8770,8773
mg|8774,8776
Tablet|8777,8783
Sig|8784,8787
:|8787,8788
One|8789,8792
(|8793,8794
1|8794,8795
)|8795,8796
Tablet|8797,8803
PO|8804,8806
Once|8807,8811
Daily|8812,8817
at|8818,8820
4|8821,8822
<EOL>|8823,8824
_|8824,8825
_|8825,8826
_|8826,8827
.|8827,8828
<EOL>|8830,8831
7.|8831,8833
Torsemide|8834,8843
5|8844,8845
mg|8846,8848
Tablet|8849,8855
Sig|8856,8859
:|8859,8860
One|8861,8864
(|8865,8866
1|8866,8867
)|8867,8868
Tablet|8869,8875
PO|8876,8878
DAILY|8879,8884
(|8885,8886
Daily|8886,8891
)|8891,8892
.|8892,8893
<EOL>|8895,8896
8.|8896,8898
Glipizide|8899,8908
10|8909,8911
mg|8912,8914
Tablet|8915,8921
Sig|8922,8925
:|8925,8926
One|8927,8930
(|8931,8932
1|8932,8933
)|8933,8934
Tablet|8935,8941
PO|8942,8944
BID|8945,8948
(|8949,8950
2|8950,8951
times|8952,8957
a|8958,8959
<EOL>|8960,8961
day|8961,8964
)|8964,8965
.|8965,8966
<EOL>|8968,8969
<EOL>|8969,8970
<EOL>|8971,8972
Discharge|8972,8981
Disposition|8982,8993
:|8993,8994
<EOL>|8994,8995
Extended|8995,9003
Care|9004,9008
<EOL>|9008,9009
<EOL>|9010,9011
Facility|9011,9019
:|9019,9020
<EOL>|9020,9021
-|9021,9022
<EOL>|9022,9023
<EOL>|9024,9025
Discharge|9025,9034
Diagnosis|9035,9044
:|9044,9045
<EOL>|9045,9046
Left|9046,9050
frontal|9051,9058
meningioma|9059,9069
,|9069,9070
left|9071,9075
parietal|9076,9084
sub-acute|9085,9094
infarct|9095,9102
,|9102,9103
<EOL>|9104,9105
Diabetes|9105,9113
<EOL>|9113,9114
<EOL>|9114,9115
<EOL>|9116,9117
Mental|9138,9144
Status|9145,9151
:|9151,9152
Confused|9153,9161
-|9162,9163
sometimes|9164,9173
.|9173,9174
<EOL>|9174,9175
Level|9175,9180
of|9181,9183
Consciousness|9184,9197
:|9197,9198
Alert|9199,9204
and|9205,9208
interactive|9209,9220
.|9220,9221
<EOL>|9221,9222
Activity|9222,9230
Status|9231,9237
:|9237,9238
Ambulatory|9239,9249
-|9250,9251
requires|9252,9260
assistance|9261,9271
or|9272,9274
aid|9275,9278
(|9279,9280
walker|9280,9286
<EOL>|9287,9288
or|9288,9290
cane|9291,9295
)|9295,9296
.|9296,9297
<EOL>|9297,9298
<EOL>|9298,9299
<EOL>|9300,9301
You|9325,9328
should|9329,9335
take|9336,9340
your|9341,9345
coumadin|9346,9354
as|9355,9357
prescribed|9358,9368
.|9368,9369
<EOL>|9369,9370
You|9370,9373
do|9374,9376
not|9377,9380
need|9381,9385
anti-seizure|9386,9398
medications|9399,9410
any|9411,9414
longer|9415,9421
.|9421,9422
<EOL>|9422,9423
You|9423,9426
should|9427,9433
follow|9434,9440
up|9441,9443
with|9444,9448
Dr.|9449,9452
_|9453,9454
_|9454,9455
_|9455,9456
Dr.|9457,9460
_|9461,9462
_|9462,9463
_|9463,9464
as|9465,9467
<EOL>|9468,9469
listed|9469,9475
below|9476,9481
.|9481,9482
You|9483,9486
will|9487,9491
need|9492,9496
a|9497,9498
follow|9499,9505
up|9506,9508
MRI|9509,9512
to|9513,9515
evaluate|9516,9524
the|9525,9528
<EOL>|9529,9530
small|9530,9535
stroke|9536,9542
you|9543,9546
had|9547,9550
on|9551,9553
the|9554,9557
left|9558,9562
side|9563,9567
of|9568,9570
your|9571,9575
brain|9576,9581
.|9581,9582
Take|9583,9587
all|9588,9591
<EOL>|9592,9593
medications|9593,9604
as|9605,9607
prescribed|9608,9618
and|9619,9622
follow|9623,9629
up|9630,9632
with|9633,9637
Dr.|9638,9641
_|9642,9643
_|9643,9644
_|9644,9645
<EOL>|9646,9647
this|9647,9651
week|9652,9656
to|9657,9659
check|9660,9665
in|9666,9668
.|9668,9669
<EOL>|9669,9670
<EOL>|9670,9671
General|9671,9678
Instructions|9679,9691
/|9691,9692
Information|9692,9703
<EOL>|9703,9704
|9704,9705
Take|9705,9709
your|9710,9714
pain|9715,9719
medicine|9720,9728
as|9729,9731
prescribed|9732,9742
.|9742,9743
<EOL>|9743,9744
|9744,9745
Exercise|9745,9753
should|9754,9760
be|9761,9763
limited|9764,9771
to|9772,9774
walking|9775,9782
;|9782,9783
no|9784,9786
lifting|9787,9794
,|9794,9795
straining|9796,9805
,|9805,9806
<EOL>|9807,9808
or|9808,9810
excessive|9811,9820
bending|9821,9828
.|9828,9829
<EOL>|9829,9830
|9830,9831
Increase|9831,9839
your|9840,9844
intake|9845,9851
of|9852,9854
fluids|9855,9861
and|9862,9865
fiber|9866,9871
,|9871,9872
as|9873,9875
narcotic|9876,9884
pain|9885,9889
<EOL>|9890,9891
medicine|9891,9899
can|9900,9903
cause|9904,9909
constipation|9910,9922
.|9922,9923
We|9924,9926
generally|9927,9936
recommend|9937,9946
taking|9947,9953
<EOL>|9954,9955
an|9955,9957
over|9958,9962
the|9963,9966
counter|9967,9974
stool|9975,9980
softener|9981,9989
,|9989,9990
such|9991,9995
as|9996,9998
Docusate|9999,10007
(|10008,10009
Colace|10009,10015
)|10015,10016
<EOL>|10017,10018
while|10018,10023
taking|10024,10030
narcotic|10031,10039
pain|10040,10044
medication|10045,10055
.|10055,10056
<EOL>|10056,10057
|10057,10058
Unless|10058,10064
directed|10065,10073
by|10074,10076
your|10077,10081
doctor|10082,10088
,|10088,10089
do|10090,10092
not|10093,10096
take|10097,10101
any|10102,10105
<EOL>|10106,10107
anti-inflammatory|10107,10124
medicines|10125,10134
such|10135,10139
as|10140,10142
Motrin|10143,10149
,|10149,10150
Aspirin|10151,10158
,|10158,10159
Advil|10160,10165
,|10165,10166
and|10167,10170
<EOL>|10171,10172
Ibuprofen|10172,10181
etc|10182,10185
.|10185,10186
<EOL>|10188,10189
|10189,10190
If|10191,10193
you|10194,10197
are|10198,10201
being|10202,10207
sent|10208,10212
home|10213,10217
on|10218,10220
steroid|10221,10228
medication|10229,10239
,|10239,10240
make|10241,10245
sure|10246,10250
<EOL>|10251,10252
you|10252,10255
are|10256,10259
taking|10260,10266
a|10267,10268
medication|10269,10279
to|10280,10282
protect|10283,10290
your|10291,10295
stomach|10296,10303
(|10304,10305
Prilosec|10305,10313
,|10313,10314
<EOL>|10315,10316
Protonix|10316,10324
,|10324,10325
or|10326,10328
Pepcid|10329,10335
)|10335,10336
,|10336,10337
as|10338,10340
these|10341,10346
medications|10347,10358
can|10359,10362
cause|10363,10368
stomach|10369,10376
<EOL>|10377,10378
irritation|10378,10388
.|10388,10389
Make|10391,10395
sure|10396,10400
to|10401,10403
take|10404,10408
your|10409,10413
steroid|10414,10421
medication|10422,10432
with|10433,10437
<EOL>|10438,10439
meals|10439,10444
,|10444,10445
or|10446,10448
a|10449,10450
glass|10451,10456
of|10457,10459
milk|10460,10464
.|10464,10465
<EOL>|10466,10467
|10467,10468
Clearance|10468,10477
to|10478,10480
drive|10481,10486
and|10487,10490
return|10491,10497
to|10498,10500
work|10501,10505
will|10506,10510
be|10511,10513
addressed|10514,10523
at|10524,10526
your|10527,10531
<EOL>|10532,10533
post-operative|10533,10547
office|10548,10554
visit|10555,10560
.|10560,10561
<EOL>|10561,10562
|10562,10563
Make|10563,10567
sure|10568,10572
to|10573,10575
continue|10576,10584
to|10585,10587
use|10588,10591
your|10592,10596
incentive|10597,10606
spirometer|10607,10617
while|10618,10623
<EOL>|10624,10625
at|10625,10627
home|10628,10632
.|10632,10633
<EOL>|10633,10634
CALL|10634,10638
YOUR|10639,10643
SURGEON|10644,10651
IMMEDIATELY|10652,10663
IF|10664,10666
YOU|10667,10670
EXPERIENCE|10671,10681
ANY|10682,10685
OF|10686,10688
THE|10689,10692
<EOL>|10693,10694
FOLLOWING|10694,10703
<EOL>|10703,10704
<EOL>|10704,10705
|10705,10706
New|10706,10709
onset|10710,10715
of|10716,10718
tremors|10719,10726
or|10727,10729
seizures|10730,10738
.|10738,10739
<EOL>|10739,10740
|10740,10741
Any|10741,10744
confusion|10745,10754
or|10755,10757
change|10758,10764
in|10765,10767
mental|10768,10774
status|10775,10781
.|10781,10782
<EOL>|10783,10784
|10784,10785
Any|10785,10788
numbness|10789,10797
,|10797,10798
tingling|10799,10807
,|10807,10808
weakness|10809,10817
in|10818,10820
your|10821,10825
extremities|10826,10837
.|10837,10838
<EOL>|10838,10839
|10839,10840
Pain|10840,10844
or|10845,10847
headache|10848,10856
that|10857,10861
is|10862,10864
continually|10865,10876
increasing|10877,10887
,|10887,10888
or|10889,10891
not|10892,10895
<EOL>|10896,10897
relieved|10897,10905
by|10906,10908
pain|10909,10913
medication|10914,10924
.|10924,10925
<EOL>|10925,10926
|10926,10927
Fever|10927,10932
greater|10933,10940
than|10941,10945
or|10946,10948
equal|10949,10954
to|10955,10957
101|10958,10961
°|10961,10962
F|10963,10964
.|10964,10965
<EOL>|10965,10966
<EOL>|10966,10967
<EOL>|10968,10969
Followup|10969,10977
Instructions|10978,10990
:|10990,10991
<EOL>|10991,10992
_|10992,10993
_|10993,10994
_|10994,10995
<EOL>|10995,10996

