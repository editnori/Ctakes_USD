 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|185,194|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|210,219|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|222,231|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|246,255|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|257,266|false|false|false|C0018965|Hematuria|Hematuria
Event|Event|SIMPLE_SEGMENT|257,266|false|false|false|||Hematuria
Event|Event|SIMPLE_SEGMENT|268,276|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|268,276|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Classification|SIMPLE_SEGMENT|279,284|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|285,293|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|285,293|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|297,315|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|306,315|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|306,315|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|306,315|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|306,315|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|306,315|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|325,332|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|325,332|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|325,332|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|325,332|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|325,335|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|325,351|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|325,351|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|336,343|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|336,343|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|336,351|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|344,351|true|false|false|C0221423|Illness (finding)|Illness
Drug|Organic Chemical|SIMPLE_SEGMENT|384,391|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|384,391|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|384,391|false|false|false|||lovenox
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|394,401|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|394,401|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|394,401|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|394,401|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|394,408|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|402,408|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|402,408|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|423,426|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|423,426|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|427,430|false|false|false|||BSO
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|432,435|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|432,435|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|432,435|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|432,435|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|432,435|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|432,435|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|432,435|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|436,443|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|436,454|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|444,454|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|444,454|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|460,465|false|false|false|C0020885|ileum|ileal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|460,470|false|false|false|C1550266|Ileal Loop|ileal loop
Event|Event|SIMPLE_SEGMENT|472,481|false|false|false|||diversion
Finding|Finding|SIMPLE_SEGMENT|472,481|false|false|false|C0439843;C3840275|Diversion|diversion
Finding|Functional Concept|SIMPLE_SEGMENT|472,481|false|false|false|C0439843;C3840275|Diversion|diversion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|472,481|false|false|false|C0185033|Diversion procedure|diversion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|486,494|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|495,506|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|495,506|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Location or Region|SIMPLE_SEGMENT|518,527|false|false|false|C0000726|Abdomen|abdominal
Drug|Substance|SIMPLE_SEGMENT|529,534|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|529,534|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|529,534|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|535,544|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|545,554|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|545,554|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|545,554|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|558,566|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|558,566|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|558,566|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|558,566|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|567,576|false|false|false|||catheters
Anatomy|Body Location or Region|SIMPLE_SEGMENT|586,595|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|586,603|false|false|false|C4481095|abdominal imaging|abdominal imaging
Event|Event|SIMPLE_SEGMENT|596,603|false|false|false|||imaging
Finding|Finding|SIMPLE_SEGMENT|596,603|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|596,603|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|SIMPLE_SEGMENT|604,609|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|610,619|false|false|false|||worsening
Finding|Idea or Concept|SIMPLE_SEGMENT|610,619|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|SIMPLE_SEGMENT|637,643|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|637,643|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|637,643|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|645,659|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|645,659|false|false|false|||hydronephrosis
Event|Event|SIMPLE_SEGMENT|675,680|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|689,694|false|false|false|||risen
Finding|Intellectual Product|SIMPLE_SEGMENT|712,723|false|false|false|C1547992|Outside Lab|outside lab
Finding|Gene or Genome|SIMPLE_SEGMENT|720,723|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|720,723|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Event|Event|SIMPLE_SEGMENT|724,729|false|false|false|||value
Finding|Intellectual Product|SIMPLE_SEGMENT|724,729|false|false|false|C1554112|MDF Attribute Type - Value|value
Finding|Body Substance|SIMPLE_SEGMENT|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|749,758|false|false|false|||underwent
Event|Event|SIMPLE_SEGMENT|770,781|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|770,781|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|770,781|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|770,796|false|false|false|C0948143|Nephrostomy tube placement|nephrostomy tube placement
Event|Event|SIMPLE_SEGMENT|782,786|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|782,786|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|782,786|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|782,796|false|false|false|C0883304|placement of tube|tube placement
Event|Event|SIMPLE_SEGMENT|787,796|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|787,796|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|787,796|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|823,830|false|false|false|||started
Finding|Sign or Symptom|SIMPLE_SEGMENT|831,843|false|false|false|C3714552|Weakness|feeling weak
Event|Event|SIMPLE_SEGMENT|839,843|false|false|false|||weak
Finding|Intellectual Product|SIMPLE_SEGMENT|839,843|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|839,843|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|SIMPLE_SEGMENT|876,885|false|false|false|||exercises
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|876,885|false|false|false|C0015259|Exercise|exercises
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|876,885|false|false|false|C0452240|Physical therapy exercises|exercises
Event|Event|SIMPLE_SEGMENT|891,903|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|891,903|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|909,919|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|909,919|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|909,919|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|SIMPLE_SEGMENT|925,934|false|false|false|||tightness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|939,944|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|939,944|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|950,960|false|false|false|||ambulating
Event|Event|SIMPLE_SEGMENT|967,976|false|false|false|||yesterday
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|983,988|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|983,988|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|983,988|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|983,988|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|983,988|false|false|false|C0031765|Phototherapy|light
Event|Event|SIMPLE_SEGMENT|989,995|false|false|false|||headed
Event|Event|SIMPLE_SEGMENT|1002,1012|false|false|false|||ambulation
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1002,1012|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|SIMPLE_SEGMENT|1002,1012|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Event|Event|SIMPLE_SEGMENT|1018,1025|false|false|false|||noticed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1036,1045|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|1036,1045|false|false|false|||hematuria
Finding|Intellectual Product|SIMPLE_SEGMENT|1053,1056|false|false|false|C1552710|Bag Data Type|bag
Event|Event|SIMPLE_SEGMENT|1057,1063|false|false|false|||darker
Event|Event|SIMPLE_SEGMENT|1072,1075|false|false|false|||bag
Finding|Intellectual Product|SIMPLE_SEGMENT|1072,1075|false|false|false|C1552710|Bag Data Type|bag
Event|Event|SIMPLE_SEGMENT|1082,1091|false|false|false|||yesterday
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1097,1105|false|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1097,1105|false|false|false|C0856443|Urostomy procedure|Urostomy
Event|Event|SIMPLE_SEGMENT|1107,1113|false|false|false|||placed
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1127,1135|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|1127,1135|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|1127,1135|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|1127,1135|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|1127,1139|false|false|false|C1446409|Positive|positive for
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1140,1149|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|1140,1149|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|1159,1170|false|false|false|||transferred
Event|Event|SIMPLE_SEGMENT|1194,1204|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|1194,1204|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|1194,1204|false|false|false|C0376636|Disease Management|management
Finding|Idea or Concept|SIMPLE_SEGMENT|1218,1225|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|SIMPLE_SEGMENT|1226,1232|false|false|false|||vitals
Event|Event|SIMPLE_SEGMENT|1242,1246|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1242,1246|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1242,1246|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1291,1295|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1296,1303|false|false|false|||notable
Anatomy|Cell|SIMPLE_SEGMENT|1311,1314|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|1328,1337|false|false|false|C0005821|Blood Platelets|platelets
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1328,1337|false|false|false|C0443116|Platelets Product|platelets
Event|Event|SIMPLE_SEGMENT|1328,1337|false|false|false|||platelets
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1328,1337|false|false|false|C0032181|Platelet count (procedure)|platelets
Event|Event|SIMPLE_SEGMENT|1366,1372|false|false|false|||biacrb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1378,1381|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1378,1381|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|1378,1381|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1378,1381|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Event|Event|SIMPLE_SEGMENT|1394,1396|false|false|false|||UA
Event|Event|SIMPLE_SEGMENT|1412,1423|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|1412,1423|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1412,1423|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Event|Event|SIMPLE_SEGMENT|1424,1429|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|1424,1429|false|false|false|C1547937||tubes
Anatomy|Cell|SIMPLE_SEGMENT|1441,1444|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1446,1454|false|false|false|||moderate
Finding|Finding|SIMPLE_SEGMENT|1446,1454|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|SIMPLE_SEGMENT|1446,1454|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Cell|SIMPLE_SEGMENT|1456,1466|false|false|false|C0023516|Leukocytes|leukocytes
Event|Event|SIMPLE_SEGMENT|1456,1466|false|false|false|||leukocytes
Finding|Body Substance|SIMPLE_SEGMENT|1456,1466|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Finding|Intellectual Product|SIMPLE_SEGMENT|1456,1466|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Finding|Gene or Genome|SIMPLE_SEGMENT|1472,1477|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1478,1483|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|1478,1483|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|1478,1483|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|1488,1495|false|false|false|||Imaging
Finding|Finding|SIMPLE_SEGMENT|1488,1495|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1488,1495|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|SIMPLE_SEGMENT|1500,1507|false|false|false|||notable
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1514,1520|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1517,1520|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|1517,1520|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1521,1527|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1521,1527|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1521,1527|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Event|Event|SIMPLE_SEGMENT|1521,1527|false|false|false|||pelvis
Finding|Finding|SIMPLE_SEGMENT|1521,1527|false|false|false|C0812455|Pelvis problem|pelvis
Event|Event|SIMPLE_SEGMENT|1529,1530|false|false|false|||/
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1532,1540|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|1532,1540|false|false|false|||contrast
Finding|Intellectual Product|SIMPLE_SEGMENT|1542,1550|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|1551,1560|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|1551,1560|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1551,1560|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|SIMPLE_SEGMENT|1574,1586|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|SIMPLE_SEGMENT|1587,1605|false|false|false|||nephroureterostomy
Event|Event|SIMPLE_SEGMENT|1607,1612|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|1607,1612|false|false|false|C1547937||tubes
Finding|Conceptual Entity|SIMPLE_SEGMENT|1618,1626|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|SIMPLE_SEGMENT|1618,1626|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1627,1648|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Event|Event|SIMPLE_SEGMENT|1627,1648|false|false|false|||hydroureteronephrosis
Event|Event|SIMPLE_SEGMENT|1656,1664|true|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|1656,1664|true|false|false|C0018944|Hematoma|hematoma
Finding|Body Substance|SIMPLE_SEGMENT|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Activity|SIMPLE_SEGMENT|1700,1707|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|1700,1707|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|1700,1707|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1715,1720|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1730,1737|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1747,1754|false|false|false|||noticed
Event|Event|SIMPLE_SEGMENT|1756,1765|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1756,1775|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|1756,1775|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|1769,1775|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|1787,1794|false|false|false|||walking
Event|Event|SIMPLE_SEGMENT|1798,1809|false|false|false|||conjunction
Finding|Idea or Concept|SIMPLE_SEGMENT|1798,1809|false|false|false|C2699427|Conjunction|conjunction
Finding|Finding|SIMPLE_SEGMENT|1816,1822|false|false|false|C4554530|Bloody|bloody
Event|Event|SIMPLE_SEGMENT|1823,1829|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|1823,1829|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|1823,1829|false|false|false|C3251815|Measurement of fluid output|output
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1839,1845|false|false|false|C0029473|Ostomy|ostomy
Event|Event|SIMPLE_SEGMENT|1846,1851|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|1846,1851|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|1857,1862|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|1872,1878|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|1872,1878|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|1872,1878|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|1889,1900|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|1889,1900|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1889,1900|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Event|Event|SIMPLE_SEGMENT|1901,1906|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|1901,1906|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|1916,1922|false|false|false|||tinged
Finding|Idea or Concept|SIMPLE_SEGMENT|1942,1950|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Gene or Genome|SIMPLE_SEGMENT|1958,1961|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|SIMPLE_SEGMENT|1972,1980|false|false|false|||endorses
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1992,1997|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1992,1997|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1999,2008|false|false|false|||tightness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2016,2020|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2016,2020|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2016,2020|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2016,2020|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2024,2032|true|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|2024,2032|true|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|2038,2044|false|false|false|||denies
Drug|Organic Chemical|SIMPLE_SEGMENT|2045,2050|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2045,2050|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2045,2050|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2045,2050|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|2052,2057|true|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|2052,2057|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|2052,2057|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|2060,2066|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|2060,2066|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2068,2077|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|2068,2082|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2078,2082|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2078,2082|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2078,2082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2078,2082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|2087,2095|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|2087,2095|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2087,2095|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|2101,2106|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|2124,2130|true|false|false|||ostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2124,2130|true|false|false|C0029473|Ostomy|ostomy
Event|Event|SIMPLE_SEGMENT|2135,2153|true|false|false|||nephroureterostomy
Event|Event|SIMPLE_SEGMENT|2162,2171|true|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|2162,2171|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2162,2171|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2162,2171|true|false|false|C2229507|sensory exam|sensation
Event|Event|SIMPLE_SEGMENT|2175,2182|true|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|2175,2182|true|false|false|C0013428|Dysuria|dysuria
Finding|Body Substance|SIMPLE_SEGMENT|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|2193,2198|false|false|false|||notes
Event|Event|SIMPLE_SEGMENT|2199,2206|false|false|false|||feeling
Finding|Sign or Symptom|SIMPLE_SEGMENT|2199,2212|false|false|false|C0849959|feeling dizzy|feeling dizzy
Event|Event|SIMPLE_SEGMENT|2207,2212|false|false|false|||dizzy
Finding|Sign or Symptom|SIMPLE_SEGMENT|2207,2212|false|false|false|C0012833|Dizziness|dizzy
Event|Event|SIMPLE_SEGMENT|2217,2228|false|false|false|||lightheaded
Finding|Sign or Symptom|SIMPLE_SEGMENT|2217,2228|false|false|false|C0220870|Lightheadedness|lightheaded
Event|Event|SIMPLE_SEGMENT|2261,2273|false|false|false|||asymptomatic
Finding|Finding|SIMPLE_SEGMENT|2261,2273|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Finding|SIMPLE_SEGMENT|2279,2299|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2284,2291|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2284,2291|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2284,2291|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2284,2291|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2284,2291|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2284,2299|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2292,2299|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2292,2299|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2292,2299|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2303,2315|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|2303,2315|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2325,2328|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2325,2328|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|2325,2328|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|2325,2328|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|2325,2328|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|2325,2328|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2325,2328|false|false|false|C0031150|Laparoscopy|lap
Event|Event|SIMPLE_SEGMENT|2329,2334|false|false|false|||chole
Finding|Functional Concept|SIMPLE_SEGMENT|2344,2348|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2344,2353|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2344,2353|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2349,2353|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2349,2365|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2349,2365|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Event|Event|SIMPLE_SEGMENT|2354,2365|false|false|false|||replacement
Finding|Functional Concept|SIMPLE_SEGMENT|2354,2365|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|2354,2365|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2354,2365|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|SIMPLE_SEGMENT|2375,2386|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2375,2386|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2399,2402|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2399,2402|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|2399,2402|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2412,2419|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2412,2419|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2412,2419|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2412,2426|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder Cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2420,2426|false|false|false|C0006826|Malignant Neoplasms|Cancer
Event|Event|SIMPLE_SEGMENT|2420,2426|false|false|false|||Cancer
Finding|Finding|SIMPLE_SEGMENT|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|2427,2437|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|SIMPLE_SEGMENT|2427,2437|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|SIMPLE_SEGMENT|2432,2437|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|2432,2437|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|SIMPLE_SEGMENT|2438,2441|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2438,2441|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|SIMPLE_SEGMENT|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Event|Event|SIMPLE_SEGMENT|2438,2441|false|false|false|||TCC
Event|Event|SIMPLE_SEGMENT|2446,2455|false|false|false|||diagnosed
Finding|Intellectual Product|SIMPLE_SEGMENT|2464,2468|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2474,2480|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2474,2484|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Event|Event|SIMPLE_SEGMENT|2481,2484|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|2481,2484|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2481,2484|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|2481,2484|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2487,2495|false|false|false|C1269955|Tumor Cell Invasion|invasion
Event|Event|SIMPLE_SEGMENT|2487,2495|false|false|false|||invasion
Finding|Pathologic Function|SIMPLE_SEGMENT|2487,2495|false|false|false|C2699153|Cell Invasion|invasion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2501,2508|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2501,2508|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2501,2508|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2501,2513|false|false|false|C0458421|Wall of bladder|bladder wall
Event|Event|SIMPLE_SEGMENT|2515,2526|false|false|false|||perivesical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2528,2532|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2528,2539|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|2528,2539|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|2533,2539|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|2533,2539|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2544,2552|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2553,2560|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2553,2560|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|2553,2560|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|2553,2560|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2553,2565|false|false|false|C0447612|Vaginal wall|vaginal wall
Event|Event|SIMPLE_SEGMENT|2567,2568|false|false|false|||/
Event|Event|SIMPLE_SEGMENT|2573,2580|false|false|false|||staging
Finding|Functional Concept|SIMPLE_SEGMENT|2573,2580|false|false|false|C0332305|With staging|staging
Event|Event|SIMPLE_SEGMENT|2590,2602|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|2590,2602|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2590,2602|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2607,2629|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|SIMPLE_SEGMENT|2617,2629|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2617,2629|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|SIMPLE_SEGMENT|2634,2639|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|SIMPLE_SEGMENT|2634,2646|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2640,2646|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|SIMPLE_SEGMENT|2640,2646|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2640,2646|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2640,2646|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|SIMPLE_SEGMENT|2640,2646|false|false|false|||uterus
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2640,2646|false|false|false|C0869889|examination of uterus|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2650,2657|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|SIMPLE_SEGMENT|2650,2657|false|false|false|||fibroid
Event|Event|SIMPLE_SEGMENT|2676,2677|false|false|false|||b
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2680,2686|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2680,2697|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|SIMPLE_SEGMENT|2687,2692|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2687,2697|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|SIMPLE_SEGMENT|2698,2707|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2698,2707|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2714,2721|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2714,2732|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|2722,2732|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2722,2732|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2737,2745|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|2746,2757|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2746,2757|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2763,2770|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2763,2770|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|2763,2770|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|2763,2770|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|SIMPLE_SEGMENT|2772,2786|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|2772,2786|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2772,2786|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2792,2797|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2792,2805|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2792,2805|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|SIMPLE_SEGMENT|2806,2814|false|false|false|C1706214|Creation|creation
Event|Event|SIMPLE_SEGMENT|2806,2814|false|false|false|||creation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2806,2814|false|false|false|C0441513|Surgical construction|creation
Event|Event|SIMPLE_SEGMENT|2828,2839|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|2843,2853|false|false|false|||bacteremia
Finding|Finding|SIMPLE_SEGMENT|2843,2853|false|false|false|C0004610|Bacteremia|bacteremia
Event|Event|SIMPLE_SEGMENT|2858,2869|true|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|2858,2869|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|2858,2869|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Event|Event|SIMPLE_SEGMENT|2873,2888|true|false|false|||intra-abdominal
Finding|Functional Concept|SIMPLE_SEGMENT|2873,2888|true|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|SIMPLE_SEGMENT|2890,2895|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2890,2895|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|2896,2906|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|2896,2906|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|2896,2906|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|2896,2906|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|2896,2906|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|2915,2920|true|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|2915,2920|true|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2915,2930|true|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|2921,2930|true|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|2921,2930|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2921,2930|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|2948,2949|false|false|false|||/
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2955,2958|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2955,2958|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2955,2958|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|2955,2958|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|2963,2965|false|false|false|||PE
Drug|Organic Chemical|SIMPLE_SEGMENT|2969,2976|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2969,2976|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|2969,2976|false|false|false|||lovenox
Finding|Functional Concept|SIMPLE_SEGMENT|2982,2988|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2982,2996|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2989,2996|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2989,2996|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2989,2996|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2989,2996|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3002,3008|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3002,3008|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3002,3008|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3002,3008|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3002,3016|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3009,3016|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3009,3016|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3009,3016|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3009,3016|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|3018,3026|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|3018,3026|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|3018,3026|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3018,3026|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|SIMPLE_SEGMENT|3018,3030|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3031,3038|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3031,3038|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|3031,3038|true|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3031,3038|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3031,3041|true|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Event|Event|SIMPLE_SEGMENT|3046,3054|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3046,3054|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3046,3054|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3046,3054|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3046,3059|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3046,3059|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3055,3059|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3055,3059|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3055,3059|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3087,3096|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3097,3105|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3097,3105|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3097,3105|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3097,3105|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3097,3110|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3097,3110|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|3106,3110|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3106,3110|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3106,3110|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|SIMPLE_SEGMENT|3140,3145|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|VITAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3140,3151|false|false|false|C0488614;C0518766|Vital signs|VITAL SIGNS
Procedure|Health Care Activity|SIMPLE_SEGMENT|3140,3151|false|false|false|C0150404|Taking vital signs|VITAL SIGNS
Event|Event|SIMPLE_SEGMENT|3146,3151|false|false|false|||SIGNS
Finding|Finding|SIMPLE_SEGMENT|3146,3151|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|SIGNS
Finding|Functional Concept|SIMPLE_SEGMENT|3146,3151|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|SIGNS
Event|Event|SIMPLE_SEGMENT|3153,3157|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|3153,3157|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3153,3157|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3191,3195|false|false|false|C2317096|Saturation of Peripheral Oxygen|Spo2
Event|Event|SIMPLE_SEGMENT|3203,3210|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3203,3210|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3203,3210|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|3212,3216|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3217,3226|true|false|false|||appearing
Finding|Finding|SIMPLE_SEGMENT|3241,3261|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|3247,3252|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|3253,3261|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|3253,3261|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3253,3261|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3263,3270|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3263,3270|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|3272,3275|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|3280,3287|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|3280,3287|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3288,3293|true|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|3295,3300|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3295,3300|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|3304,3316|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3304,3316|false|false|false|C0004339|Auscultation|auscultation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3330,3337|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3330,3337|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3330,3337|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3330,3337|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3339,3343|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3339,3343|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3359,3368|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3359,3368|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3377,3382|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|3377,3389|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|3383,3389|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3383,3389|false|false|false|C0037709||sounds
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3392,3398|false|false|false|C0029473|Ostomy|Ostomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3408,3413|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Finding|Finding|SIMPLE_SEGMENT|3408,3419|false|false|false|C5880922|Brown color of stool|brown stool
Event|Event|SIMPLE_SEGMENT|3414,3419|false|false|false|||stool
Finding|Body Substance|SIMPLE_SEGMENT|3414,3419|false|false|false|C0015733|Feces|stool
Finding|Finding|SIMPLE_SEGMENT|3455,3458|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|3455,3458|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Finding|SIMPLE_SEGMENT|3459,3465|false|false|false|C4554530|Bloody|bloody
Finding|Finding|SIMPLE_SEGMENT|3459,3471|false|false|false|C0473237|Frank hematuria|bloody urine
Event|Event|SIMPLE_SEGMENT|3466,3471|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|3483,3494|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|3483,3494|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3483,3494|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Event|Event|SIMPLE_SEGMENT|3495,3500|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|3495,3500|false|false|false|C1547937||tubes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3510,3515|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|3510,3515|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|3510,3515|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|3517,3522|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3525,3536|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3541,3546|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3541,3546|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3541,3546|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3548,3552|true|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3548,3552|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3548,3552|true|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3557,3561|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3562,3570|true|false|false|||perfused
Finding|Body Substance|SIMPLE_SEGMENT|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3599,3608|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3609,3617|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3609,3617|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|3609,3617|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3609,3617|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|3609,3622|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3609,3622|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|3618,3622|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3618,3622|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3618,3622|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|3686,3693|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|3686,3693|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3686,3693|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|SIMPLE_SEGMENT|3695,3699|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3700,3709|true|false|false|||appearing
Finding|Finding|SIMPLE_SEGMENT|3724,3744|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|SIMPLE_SEGMENT|3730,3735|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|3736,3744|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|3736,3744|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|3736,3744|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3746,3753|true|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3746,3753|true|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|SIMPLE_SEGMENT|3755,3758|true|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|3763,3770|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|3763,3770|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3771,3776|true|false|false|C0024109|Lung|LUNGS
Event|Event|SIMPLE_SEGMENT|3778,3783|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3778,3783|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|3787,3799|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3787,3799|false|false|false|C0004339|Auscultation|auscultation
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3813,3820|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3813,3820|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|SIMPLE_SEGMENT|3813,3820|false|false|false|||ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3813,3820|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3822,3826|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3822,3826|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3842,3851|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3842,3851|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3860,3865|false|false|false|C0021853|Intestines|bowel
Finding|Finding|SIMPLE_SEGMENT|3860,3872|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|SIMPLE_SEGMENT|3866,3872|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3866,3872|false|false|false|C0037709||sounds
Finding|Finding|SIMPLE_SEGMENT|3909,3912|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|SIMPLE_SEGMENT|3909,3912|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Finding|SIMPLE_SEGMENT|3913,3919|false|false|false|C4554530|Bloody|bloody
Finding|Finding|SIMPLE_SEGMENT|3913,3925|false|false|false|C0473237|Frank hematuria|bloody urine
Event|Event|SIMPLE_SEGMENT|3920,3925|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|3938,3949|false|false|false|||nephrostomy
Finding|Finding|SIMPLE_SEGMENT|3938,3949|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3938,3949|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Event|Event|SIMPLE_SEGMENT|3950,3955|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|3950,3955|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|3956,3962|false|false|false|||capped
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3965,3976|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3981,3986|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3981,3986|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3981,3986|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3988,3992|true|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3988,3992|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3988,3992|true|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3997,4001|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|4002,4010|true|false|false|||perfused
Procedure|Health Care Activity|SIMPLE_SEGMENT|4050,4059|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|4060,4064|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4060,4064|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4094,4099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4094,4099|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4094,4099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4100,4103|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4108,4111|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4108,4111|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4108,4111|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4118,4121|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4118,4121|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4118,4121|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4118,4121|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4127,4130|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4127,4130|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4138,4141|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4138,4141|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4138,4141|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4145,4148|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4145,4148|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4145,4148|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4145,4148|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4145,4148|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4145,4148|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4154,4158|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4154,4158|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4186,4189|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4206,4211|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4206,4211|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4206,4211|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4212,4215|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4220,4223|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4220,4223|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4220,4223|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4230,4233|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4230,4233|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4230,4233|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4230,4233|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4239,4242|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4239,4242|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4250,4253|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4250,4253|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4250,4253|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4250,4253|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4250,4253|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4257,4260|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4257,4260|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4257,4260|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4257,4260|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4257,4260|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4257,4260|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4266,4270|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4266,4270|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4298,4301|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4318,4323|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4318,4323|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4318,4323|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|SIMPLE_SEGMENT|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4350,4353|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|4350,4353|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|4350,4353|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4453,4458|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4453,4458|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4453,4458|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4453,4466|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4453,4466|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4453,4466|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4459,4466|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4459,4466|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4459,4466|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4459,4466|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4459,4466|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4459,4466|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4513,4517|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4513,4517|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4513,4517|false|false|false|C0202059|Bicarbonate measurement|HCO3
Event|Event|SIMPLE_SEGMENT|4549,4556|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4549,4556|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4549,4556|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|4557,4564|false|false|false|||STUDIES
Procedure|Research Activity|SIMPLE_SEGMENT|4557,4564|false|false|false|C0947630|Scientific Study|STUDIES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4588,4594|false|false|false|C1644645||CT Abd
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4591,4594|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|4591,4594|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4595,4598|false|false|false|C0449203|PEL (body structure)|Pel
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4595,4598|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|Pel
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4595,4598|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|Pel
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|4603,4611|false|true|false|C0009924|Contrast Media|Contrast
Event|Event|SIMPLE_SEGMENT|4614,4624|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4614,4624|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4614,4624|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|4632,4640|false|false|false|||Interval
Finding|Intellectual Product|SIMPLE_SEGMENT|4632,4640|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|SIMPLE_SEGMENT|4641,4650|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|4641,4650|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4641,4650|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|4664,4676|false|false|false|||percutaneous
Finding|Functional Concept|SIMPLE_SEGMENT|4664,4676|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Event|Event|SIMPLE_SEGMENT|4697,4702|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|4697,4702|false|false|false|C1547937||tubes
Finding|Conceptual Entity|SIMPLE_SEGMENT|4708,4716|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|SIMPLE_SEGMENT|4708,4716|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4717,4738|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Event|Event|SIMPLE_SEGMENT|4717,4738|false|false|false|||hydroureteronephrosis
Event|Event|SIMPLE_SEGMENT|4748,4756|true|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|4748,4756|true|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|4787,4794|false|false|false|||opacity
Finding|Finding|SIMPLE_SEGMENT|4787,4794|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|SIMPLE_SEGMENT|4787,4794|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Functional Concept|SIMPLE_SEGMENT|4802,4807|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4802,4819|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|4808,4814|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4808,4819|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4815,4819|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|4815,4819|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|4843,4851|false|false|false|||assessed
Event|Event|SIMPLE_SEGMENT|4869,4878|false|false|false|||dedicated
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4879,4887|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4879,4887|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4882,4887|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Event|Event|SIMPLE_SEGMENT|4882,4887|false|false|false|||chest
Finding|Finding|SIMPLE_SEGMENT|4882,4887|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|4895,4898|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4895,4898|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|SIMPLE_SEGMENT|4911,4918|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|4911,4918|false|false|false|C1550585|Entity Handling - upright|upright
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4931,4936|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|4931,4936|false|false|false|C0741025|Chest problem|chest
Finding|Functional Concept|SIMPLE_SEGMENT|4940,4945|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4940,4961|false|false|false|C0230329|Right upper extremity|Right upper extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4946,4961|false|false|false|C1140618|Upper Extremity|upper extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4952,4961|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|SIMPLE_SEGMENT|4963,4969|false|false|false|C1554204|Role Class - access|access
Event|Event|SIMPLE_SEGMENT|4970,4974|false|false|false|||PICC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4970,4974|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|4976,4980|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|4976,4980|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|4984,4988|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|4998,5001|false|false|false|||tip
Finding|Gene or Genome|SIMPLE_SEGMENT|4998,5001|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4998,5001|false|false|false|C0673828|TIP regimen|tip
Event|Event|SIMPLE_SEGMENT|5015,5018|false|false|false|||SVC
Finding|Finding|SIMPLE_SEGMENT|5015,5018|false|false|false|C0231957|Slow vital capacity|SVC
Event|Event|SIMPLE_SEGMENT|5031,5034|false|false|false|||EKG
Finding|Intellectual Product|SIMPLE_SEGMENT|5031,5034|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5031,5034|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|SIMPLE_SEGMENT|5046,5053|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|5046,5053|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|5046,5053|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5056,5061|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|5066,5071|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|5066,5071|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|5107,5113|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|5107,5113|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|SIMPLE_SEGMENT|5116,5120|false|false|false|C0443157|Bony|Bony
Event|Event|SIMPLE_SEGMENT|5121,5131|false|false|false|||structures
Event|Event|SIMPLE_SEGMENT|5136,5142|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|5136,5142|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|5161,5173|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|5161,5173|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|5161,5173|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5161,5173|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|SIMPLE_SEGMENT|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5212,5216|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Event|Event|SIMPLE_SEGMENT|5217,5228|false|false|false|||NEPHROSTOMY
Finding|Finding|SIMPLE_SEGMENT|5217,5228|false|false|false|C0481713|Has nephrostomy|NEPHROSTOMY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5217,5228|false|false|false|C0278314|Nephrostomy (procedure)|NEPHROSTOMY
Event|Event|SIMPLE_SEGMENT|5229,5233|false|false|false|||TUBE
Finding|Functional Concept|SIMPLE_SEGMENT|5229,5233|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Finding|Gene or Genome|SIMPLE_SEGMENT|5229,5233|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Finding|Idea or Concept|SIMPLE_SEGMENT|5266,5271|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|5266,5278|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5272,5278|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|5272,5278|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|5272,5278|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|5272,5278|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|SIMPLE_SEGMENT|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5286,5299|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5292,5299|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|5292,5299|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|5292,5299|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|5292,5299|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5292,5299|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|5301,5306|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|5301,5306|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|5318,5324|true|false|false|||GROWTH
Finding|Finding|SIMPLE_SEGMENT|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|SIMPLE_SEGMENT|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|SIMPLE_SEGMENT|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5318,5324|true|false|false|C2911660|Growth action|GROWTH
Finding|Body Substance|SIMPLE_SEGMENT|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5345,5354|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|5355,5359|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5355,5359|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5389,5394|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5389,5394|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5389,5394|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5395,5398|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5403,5406|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5403,5406|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5403,5406|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5413,5416|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5413,5416|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5413,5416|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5413,5416|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5422,5425|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5422,5425|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5433,5436|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5433,5436|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5433,5436|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5433,5436|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5433,5436|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5440,5443|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5440,5443|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5440,5443|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5440,5443|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5440,5443|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5440,5443|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5449,5453|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5449,5453|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5481,5484|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5501,5506|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5501,5506|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5501,5506|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5501,5514|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5501,5514|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5501,5514|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5507,5514|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5507,5514|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5507,5514|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5507,5514|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5507,5514|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5507,5514|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5559,5563|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5559,5563|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5559,5563|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5588,5593|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5588,5593|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5588,5593|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5588,5601|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5594,5601|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5594,5601|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5594,5601|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Intellectual Product|SIMPLE_SEGMENT|5625,5630|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5631,5639|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5631,5646|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5631,5646|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Idea or Concept|SIMPLE_SEGMENT|5666,5670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|5666,5670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|5671,5674|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|5686,5693|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5686,5696|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|5697,5705|false|false|false|||provoked
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5707,5710|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5707,5710|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5707,5710|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|5707,5710|false|false|false|||DVT
Drug|Organic Chemical|SIMPLE_SEGMENT|5718,5725|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5718,5725|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|5718,5725|false|false|false|||lovenox
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5728,5735|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5728,5735|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|5728,5735|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5728,5735|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5728,5742|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5736,5742|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|5736,5742|false|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|5755,5758|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5755,5758|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|5759,5762|false|false|false|||BSO
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5764,5767|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5764,5767|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|5764,5767|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|5764,5767|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|5764,5767|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|5764,5767|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5764,5767|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5769,5776|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5769,5787|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|5777,5787|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5777,5787|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5793,5798|false|false|false|C0020885|ileum|ileal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5793,5803|false|false|false|C1550266|Ileal Loop|ileal loop
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5799,5813|false|false|false|C4489477|Loop diversion|loop diversion
Event|Event|SIMPLE_SEGMENT|5804,5813|false|false|false|||diversion
Finding|Finding|SIMPLE_SEGMENT|5804,5813|false|false|false|C0439843;C3840275|Diversion|diversion
Finding|Functional Concept|SIMPLE_SEGMENT|5804,5813|false|false|false|C0439843;C3840275|Diversion|diversion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5804,5813|false|false|false|C0185033|Diversion procedure|diversion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5818,5826|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|5818,5826|false|false|false|||anterior
Event|Event|SIMPLE_SEGMENT|5828,5839|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5828,5839|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5851,5860|false|false|false|C0000726|Abdomen|abdominal
Finding|Body Substance|SIMPLE_SEGMENT|5851,5866|false|false|false|C2699330|Abdominal Fluid|abdominal fluid
Drug|Substance|SIMPLE_SEGMENT|5861,5866|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|5861,5866|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5861,5866|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|5867,5876|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|5878,5887|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|5878,5887|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5878,5887|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|5891,5899|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|5891,5899|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|5891,5899|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5891,5899|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|5900,5909|false|false|false|||catheters
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5922,5936|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|5922,5936|false|false|false|||hydronephrosis
Event|Event|SIMPLE_SEGMENT|5938,5947|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|5948,5957|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|5948,5957|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5948,5957|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Drug|Organic Chemical|SIMPLE_SEGMENT|5971,5974|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5971,5974|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|SIMPLE_SEGMENT|5971,5974|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Event|Event|SIMPLE_SEGMENT|5975,5980|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|5975,5980|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|6006,6011|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6006,6011|false|false|false|C0034991|Rehabilitation therapy|rehab
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6017,6026|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|6017,6026|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|6031,6039|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6031,6039|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Activity|SIMPLE_SEGMENT|6045,6052|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|6045,6052|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|6045,6052|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|SIMPLE_SEGMENT|6061,6069|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|6061,6069|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|6061,6072|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6073,6078|false|false|false|C0398650|Immune thrombocytopenic purpura|frank
Finding|Finding|SIMPLE_SEGMENT|6073,6088|false|false|false|C0473237|Frank hematuria|frank hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6079,6088|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|6079,6088|false|false|false|||hematuria
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|6096,6104|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6096,6104|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Event|SIMPLE_SEGMENT|6106,6109|false|false|false|||bag
Finding|Intellectual Product|SIMPLE_SEGMENT|6106,6109|false|false|false|C1552710|Bag Data Type|bag
Drug|Organic Chemical|SIMPLE_SEGMENT|6114,6117|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6114,6117|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Event|Event|SIMPLE_SEGMENT|6114,6117|false|false|false|||PCN
Finding|Gene or Genome|SIMPLE_SEGMENT|6114,6117|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Event|Event|SIMPLE_SEGMENT|6118,6123|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|6118,6123|false|false|false|C1547937||tubes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|SIMPLE_SEGMENT|6129,6139|false|false|false|||hemoglobin
Finding|Finding|SIMPLE_SEGMENT|6129,6139|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6129,6139|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Event|Event|SIMPLE_SEGMENT|6179,6186|false|false|false|||dropped
Drug|Organic Chemical|SIMPLE_SEGMENT|6198,6205|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6198,6205|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|6198,6205|false|false|false|||lovenox
Event|Event|SIMPLE_SEGMENT|6210,6214|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|6229,6239|false|false|false|||transfused
Event|Event|SIMPLE_SEGMENT|6249,6253|false|false|false|||PRBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Event|Event|SIMPLE_SEGMENT|6274,6284|false|false|false|||hemoglobin
Finding|Finding|SIMPLE_SEGMENT|6274,6284|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6274,6284|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6299,6308|false|false|false|C0018965|Hematuria|Hematuria
Event|Event|SIMPLE_SEGMENT|6299,6308|false|false|false|||Hematuria
Finding|Finding|SIMPLE_SEGMENT|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|6320,6326|false|false|false|||caused
Finding|Mental Process|SIMPLE_SEGMENT|6361,6368|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|6372,6387|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|6372,6387|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|6372,6387|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6372,6387|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6393,6402|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|6393,6402|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|6403,6411|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|6425,6434|false|false|false|||dizziness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6425,6434|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|SIMPLE_SEGMENT|6435,6443|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6435,6443|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|6453,6462|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|6467,6479|false|false|false|||recommending
Event|Event|SIMPLE_SEGMENT|6481,6488|false|false|false|||capping
Drug|Organic Chemical|SIMPLE_SEGMENT|6493,6496|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6493,6496|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|SIMPLE_SEGMENT|6493,6496|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Event|Event|SIMPLE_SEGMENT|6497,6502|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|6497,6502|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|6510,6520|false|false|false|||discussion
Finding|Social Behavior|SIMPLE_SEGMENT|6510,6520|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6510,6520|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Body Substance|SIMPLE_SEGMENT|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6541,6553|false|false|false|||hematologist
Event|Event|SIMPLE_SEGMENT|6562,6569|false|false|false|||decided
Event|Event|SIMPLE_SEGMENT|6573,6577|false|false|false|||stop
Drug|Organic Chemical|SIMPLE_SEGMENT|6582,6589|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6582,6589|false|false|false|C0728963|Lovenox|lovenox
Event|Event|SIMPLE_SEGMENT|6590,6599|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|6590,6599|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|6590,6599|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|6590,6599|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6590,6599|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6616,6619|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6616,6619|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6616,6619|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|6616,6619|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|6628,6636|false|false|false|||provoked
Finding|Mental Process|SIMPLE_SEGMENT|6644,6651|false|false|false|C0542559|contextual factors|setting
Event|Activity|SIMPLE_SEGMENT|6659,6667|false|false|false|C0237820||recovery
Event|Event|SIMPLE_SEGMENT|6659,6667|false|false|false|||recovery
Finding|Organism Function|SIMPLE_SEGMENT|6659,6667|false|false|false|C2004454|Recovery - healing process|recovery
Event|Event|SIMPLE_SEGMENT|6674,6681|false|false|false|||surgery
Finding|Finding|SIMPLE_SEGMENT|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|SIMPLE_SEGMENT|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6674,6681|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|SIMPLE_SEGMENT|6729,6738|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|6729,6738|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|6729,6738|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|6729,6738|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6729,6738|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6741,6750|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|6741,6750|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6741,6750|false|false|false|C1522484|metastatic qualifier|Secondary
Finding|Finding|SIMPLE_SEGMENT|6762,6774|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|Asymptomatic
Event|Event|SIMPLE_SEGMENT|6775,6785|false|false|false|||bacteruria
Finding|Body Substance|SIMPLE_SEGMENT|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|SIMPLE_SEGMENT|6800,6812|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|SIMPLE_SEGMENT|6813,6823|false|false|false|||bacteruria
Finding|Mental Process|SIMPLE_SEGMENT|6828,6835|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|6857,6869|false|false|false|||manipulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6857,6869|false|false|false|C0185111;C0947647|Manipulation procedure;Surgical Manipulation|manipulation
Event|Event|SIMPLE_SEGMENT|6879,6887|true|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|6879,6887|true|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6901,6913|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|6901,6913|true|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|6901,6913|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|6918,6927|true|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|6918,6927|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|6918,6927|true|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|6918,6927|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6918,6927|true|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Antibiotic|SIMPLE_SEGMENT|6933,6944|true|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|6933,6944|true|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|6950,6958|false|false|false|||deferred
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6963,6977|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|6963,6977|false|false|false|||Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|6963,6977|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|6979,6988|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|6989,7001|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6989,7001|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|6989,7001|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7017,7031|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|7017,7031|false|false|false|||Hypothyroidism
Event|Event|SIMPLE_SEGMENT|7033,7041|false|false|false|||continue
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|7042,7055|false|false|false|||levothyroxine
Finding|Idea or Concept|SIMPLE_SEGMENT|7091,7103|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7131,7141|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Event|Event|SIMPLE_SEGMENT|7131,7141|false|false|false|||Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7131,7141|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Event|Event|SIMPLE_SEGMENT|7142,7149|false|false|false|||Changes
Finding|Functional Concept|SIMPLE_SEGMENT|7142,7149|false|false|false|C0392747|Changing|Changes
Drug|Organic Chemical|SIMPLE_SEGMENT|7151,7158|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7151,7158|false|false|false|C0728963|Lovenox|Lovenox
Event|Event|SIMPLE_SEGMENT|7159,7166|false|false|false|||stopped
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7172,7182|false|false|false|C1644645||CT Abdomen
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7172,7182|false|false|false|C0412620|CT of abdomen|CT Abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7175,7182|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7175,7182|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|7175,7182|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|7175,7182|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7183,7189|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7183,7189|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7183,7189|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|SIMPLE_SEGMENT|7183,7189|false|false|false|C0812455|Pelvis problem|Pelvis
Event|Event|SIMPLE_SEGMENT|7190,7196|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|7207,7213|false|false|false|||imaged
Event|Event|SIMPLE_SEGMENT|7222,7229|false|false|false|||opacity
Finding|Finding|SIMPLE_SEGMENT|7222,7229|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|SIMPLE_SEGMENT|7222,7229|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Functional Concept|SIMPLE_SEGMENT|7238,7243|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7238,7255|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|SIMPLE_SEGMENT|7244,7250|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7244,7255|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7251,7255|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|SIMPLE_SEGMENT|7251,7255|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|SIMPLE_SEGMENT|7277,7285|false|false|false|||assessed
Event|Event|SIMPLE_SEGMENT|7304,7313|false|false|false|||dedicated
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7314,7322|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7314,7322|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7317,7322|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Event|Event|SIMPLE_SEGMENT|7317,7322|false|false|false|||chest
Finding|Finding|SIMPLE_SEGMENT|7317,7322|false|false|false|C0741025|Chest problem|chest
Drug|Organic Chemical|SIMPLE_SEGMENT|7334,7337|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7334,7337|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|SIMPLE_SEGMENT|7334,7337|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Event|Event|SIMPLE_SEGMENT|7338,7343|false|false|false|||tubes
Finding|Intellectual Product|SIMPLE_SEGMENT|7338,7343|false|false|false|C1547937||tubes
Event|Event|SIMPLE_SEGMENT|7349,7355|false|false|false|||capped
Event|Event|SIMPLE_SEGMENT|7364,7378|false|false|false|||recommendation
Finding|Idea or Concept|SIMPLE_SEGMENT|7364,7378|false|false|false|C0034866|Recommendation|recommendation
Event|Event|SIMPLE_SEGMENT|7391,7406|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|7391,7406|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|7416,7426|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|7442,7450|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|7442,7450|false|false|false|C1522577|follow-up|followup
Event|Event|SIMPLE_SEGMENT|7455,7461|false|false|false|||decide
Finding|Idea or Concept|SIMPLE_SEGMENT|7470,7474|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|SIMPLE_SEGMENT|7470,7474|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Event|Event|SIMPLE_SEGMENT|7475,7485|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|7475,7485|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|7475,7485|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|7496,7504|false|false|false|||develops
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7505,7514|false|false|false|C0018965|Hematuria|hematuria
Event|Event|SIMPLE_SEGMENT|7505,7514|false|false|false|||hematuria
Event|Event|SIMPLE_SEGMENT|7522,7537|false|false|false|||lightheadedness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7522,7537|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|SIMPLE_SEGMENT|7548,7556|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7548,7556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7548,7556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7560,7566|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|7560,7566|false|false|false|||anemia
Anatomy|Cell Component|SIMPLE_SEGMENT|7570,7573|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|7570,7573|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7570,7573|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|SIMPLE_SEGMENT|7584,7593|false|false|false|||rechecked
Event|Event|SIMPLE_SEGMENT|7597,7603|false|false|false|||assess
Event|Event|SIMPLE_SEGMENT|7609,7617|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|7609,7617|false|false|false|C0019080|Hemorrhage|bleeding
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Organic Chemical|SIMPLE_SEGMENT|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Event|Event|SIMPLE_SEGMENT|7622,7632|false|false|false|||Hemoglobin
Finding|Finding|SIMPLE_SEGMENT|7622,7632|false|false|false|C1561562|Hemoglobin finding|Hemoglobin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7622,7632|false|false|false|C0518015|Hemoglobin measurement|Hemoglobin
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7633,7643|false|false|false|C1542366|hematocrit attribute|Hematocrit
Event|Event|SIMPLE_SEGMENT|7633,7643|false|false|false|||Hematocrit
Finding|Finding|SIMPLE_SEGMENT|7633,7643|false|false|false|C0518014|Hematocrit level|Hematocrit
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7633,7643|false|false|false|C0018935|Hematocrit Measurement|Hematocrit
Event|Event|SIMPLE_SEGMENT|7647,7656|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7647,7656|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|7670,7674|false|false|false|||CODE
Event|Occupational Activity|SIMPLE_SEGMENT|7670,7674|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|SIMPLE_SEGMENT|7670,7674|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Event|Activity|SIMPLE_SEGMENT|7692,7699|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|SIMPLE_SEGMENT|7692,7699|false|false|false|||CONTACT
Finding|Functional Concept|SIMPLE_SEGMENT|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|SIMPLE_SEGMENT|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|SIMPLE_SEGMENT|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7692,7699|false|false|false|C0392367|Physical contact|CONTACT
Anatomy|Cell|SIMPLE_SEGMENT|7715,7719|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|7715,7719|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Finding|Idea or Concept|SIMPLE_SEGMENT|7727,7731|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7727,7731|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7727,7731|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7737,7748|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7737,7748|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|7737,7748|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7737,7748|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|7737,7761|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|7752,7761|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7752,7761|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7780,7790|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7780,7790|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7780,7795|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|7791,7795|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|7791,7795|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|7799,7807|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|7812,7820|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|7812,7820|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|7812,7820|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|7825,7837|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7825,7837|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|7855,7865|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7855,7865|false|false|false|C0206460|enoxaparin|Enoxaparin
Event|Event|SIMPLE_SEGMENT|7855,7865|false|false|false|||Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|7855,7872|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7855,7872|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7866,7872|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7866,7872|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7866,7872|false|false|false|C0337443|Sodium measurement|Sodium
Event|Event|SIMPLE_SEGMENT|7888,7893|false|false|false|||Start
Finding|Idea or Concept|SIMPLE_SEGMENT|7912,7916|false|false|false|C1552851|next - HtmlLinkType|Next
Event|Event|SIMPLE_SEGMENT|7917,7924|false|false|false|||Routine
Finding|Idea or Concept|SIMPLE_SEGMENT|7917,7924|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|7917,7924|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7917,7924|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|SIMPLE_SEGMENT|7925,7939|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7925,7939|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7963,7969|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7963,7969|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7963,7969|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|7991,8004|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8007,8010|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8007,8010|false|false|false|||TAB
Anatomy|Body System|SIMPLE_SEGMENT|8034,8043|false|false|false|C0012240|Gastrointestinal system|Digestive
Finding|Organism Function|SIMPLE_SEGMENT|8034,8043|false|false|false|C0012238|Digestion|Digestive
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Enzyme|SIMPLE_SEGMENT|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8034,8051|false|false|false|C0863186|Digestive enzyme test|Digestive Enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Enzyme|SIMPLE_SEGMENT|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Event|Event|SIMPLE_SEGMENT|8044,8051|false|false|false|||Enzymes
Finding|Functional Concept|SIMPLE_SEGMENT|8044,8051|false|false|false|C0014445|enzymology|Enzymes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8068,8071|false|false|false|C1321878|Desmoplastic infantile ganglioglioma|dig
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8087,8091|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8087,8091|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|8087,8091|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|8087,8091|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|8102,8111|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8102,8111|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8102,8123|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8112,8123|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8112,8123|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8112,8123|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8112,8123|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8129,8141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8129,8141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|8175,8181|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|8175,8181|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8175,8181|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|8205,8218|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8221,8224|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|8221,8224|false|false|false|||TAB
Anatomy|Body System|SIMPLE_SEGMENT|8250,8259|false|false|false|C0012240|Gastrointestinal system|Digestive
Finding|Organism Function|SIMPLE_SEGMENT|8250,8259|false|false|false|C0012238|Digestion|Digestive
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Enzyme|SIMPLE_SEGMENT|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8250,8267|false|false|false|C0863186|Digestive enzyme test|Digestive Enzymes
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Enzyme|SIMPLE_SEGMENT|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Event|Event|SIMPLE_SEGMENT|8260,8267|false|false|false|||Enzymes
Finding|Functional Concept|SIMPLE_SEGMENT|8260,8267|false|false|false|C0014445|enzymology|Enzymes
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8284,8287|false|false|false|C1321878|Desmoplastic infantile ganglioglioma|dig
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8303,8307|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8303,8307|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|8303,8307|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|8303,8307|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|SIMPLE_SEGMENT|8319,8328|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8319,8328|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8319,8340|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|8319,8340|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8329,8340|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|8329,8340|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|8329,8340|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|8342,8350|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|8342,8350|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|8342,8355|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|8351,8355|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|8351,8355|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|8351,8355|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|8351,8355|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|8358,8366|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|8358,8366|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|8374,8383|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8374,8383|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8374,8393|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8384,8393|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|8384,8393|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|8384,8393|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|8384,8393|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8384,8393|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|SIMPLE_SEGMENT|8403,8412|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8403,8412|false|false|false|C0011900|Diagnosis|Diagnoses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8414,8423|false|false|false|C0018965|Hematuria|Hematuria
Event|Event|SIMPLE_SEGMENT|8414,8423|false|false|false|||Hematuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8425,8431|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|8425,8431|false|false|false|||anemia
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8433,8442|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|8433,8442|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|8433,8442|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|SIMPLE_SEGMENT|8443,8452|false|false|false|||Diagnoses
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8443,8452|false|false|false|C0011900|Diagnosis|Diagnoses
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8454,8461|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8454,8461|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8454,8461|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8454,8468|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8462,8468|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|8462,8468|false|false|false|||cancer
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8470,8484|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|8470,8484|false|false|false|||hydronephrosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8487,8501|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Event|Event|SIMPLE_SEGMENT|8487,8501|false|false|false|||hypothyroidism
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8503,8506|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8503,8506|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8503,8506|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|8503,8506|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|8513,8522|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8513,8522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8513,8522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8513,8522|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8513,8522|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8523,8532|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8523,8532|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|8523,8532|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|8523,8532|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|8534,8540|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8534,8547|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|8534,8547|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8541,8547|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8541,8547|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|8549,8554|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|8549,8554|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|8559,8567|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|8559,8567|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|8569,8574|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8569,8591|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|8569,8591|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|8578,8591|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|8578,8591|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|8578,8591|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8593,8598|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|8593,8598|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8593,8598|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|8593,8598|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|8603,8614|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|8603,8614|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|8616,8624|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8616,8624|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|8616,8624|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8625,8631|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|8625,8631|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|8625,8631|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|8633,8643|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|8633,8643|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|8646,8657|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|8646,8657|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|8646,8657|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|8662,8671|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8662,8671|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8662,8671|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8662,8671|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8662,8671|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8662,8684|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8662,8684|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|8662,8684|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8672,8684|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8672,8684|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8672,8684|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|8686,8690|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|8711,8719|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|8711,8719|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|8711,8719|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|8727,8731|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8727,8731|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8727,8731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8727,8731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8727,8734|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|SIMPLE_SEGMENT|8757,8760|false|false|false|||YOU
Event|Event|SIMPLE_SEGMENT|8761,8765|false|false|false|||COME
Event|Event|SIMPLE_SEGMENT|8773,8781|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|8773,8781|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|8787,8794|false|false|false|||noticed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8795,8800|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8795,8800|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8795,8800|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|8809,8814|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|8829,8836|false|false|false|||feeling
Finding|Mental Process|SIMPLE_SEGMENT|8829,8836|false|false|false|C1527305|Feelings|feeling
Finding|Intellectual Product|SIMPLE_SEGMENT|8838,8842|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|8838,8842|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|SIMPLE_SEGMENT|8843,8854|false|false|false|||lightheaded
Finding|Sign or Symptom|SIMPLE_SEGMENT|8843,8854|false|false|false|C0220870|Lightheadedness|lightheaded
Event|Activity|SIMPLE_SEGMENT|8862,8870|false|false|false|C1709305|Occur (action)|HAPPENED
Event|Event|SIMPLE_SEGMENT|8877,8880|false|false|false|||YOU
Event|Event|SIMPLE_SEGMENT|8881,8885|false|false|false|||WERE
Event|Event|SIMPLE_SEGMENT|8886,8890|false|false|false|||HERE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8917,8922|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8917,8922|true|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8917,8922|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8931,8941|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|8931,8941|true|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8931,8941|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|SIMPLE_SEGMENT|8943,8950|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8943,8950|false|false|false|C0728963|Lovenox|Lovenox
Event|Event|SIMPLE_SEGMENT|8961,8965|false|false|false|||gave
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8980,8985|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8980,8985|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8980,8985|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8991,8996|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|8991,8996|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|8991,8996|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|9005,9010|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|9011,9018|false|false|false|||cleared
Event|Event|SIMPLE_SEGMENT|9038,9041|false|false|false|||YOU
Event|Event|SIMPLE_SEGMENT|9054,9059|false|false|false|||LEAVE
Event|Event|SIMPLE_SEGMENT|9064,9072|false|false|false|||HOSPITAL
Finding|Idea or Concept|SIMPLE_SEGMENT|9064,9072|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Event|Event|SIMPLE_SEGMENT|9114,9121|true|false|false|||decided
Event|Event|SIMPLE_SEGMENT|9142,9146|true|false|false|||need
Event|Event|SIMPLE_SEGMENT|9150,9154|true|false|false|||take
Drug|Organic Chemical|SIMPLE_SEGMENT|9159,9166|true|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9159,9166|true|false|false|C0728963|Lovenox|Lovenox
Event|Event|SIMPLE_SEGMENT|9159,9166|true|false|false|||Lovenox
Event|Event|SIMPLE_SEGMENT|9179,9187|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|9192,9198|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|9212,9219|false|false|false|||doctors
Event|Event|SIMPLE_SEGMENT|9225,9229|false|false|false|||take
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9242,9253|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9242,9253|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|9242,9253|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9242,9253|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|9258,9268|false|false|false|||prescribed
Event|Event|SIMPLE_SEGMENT|9275,9283|false|false|false|||followup
Procedure|Health Care Activity|SIMPLE_SEGMENT|9275,9283|false|false|false|C1522577|follow-up|followup
Event|Activity|SIMPLE_SEGMENT|9284,9296|false|false|false|C0003629|Appointments|appointments
Event|Event|SIMPLE_SEGMENT|9284,9296|false|false|false|||appointments
Event|Event|SIMPLE_SEGMENT|9301,9307|false|false|false|||listed
Event|Event|SIMPLE_SEGMENT|9332,9340|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|9332,9340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|9332,9340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|9348,9352|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|9348,9352|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|9348,9352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9348,9352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9348,9355|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|SIMPLE_SEGMENT|9391,9399|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9400,9412|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9400,9412|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9400,9412|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

