 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
SURGERY|158,165
<EOL>|165,166
<EOL>|167,168
Allergies|168,177
:|177,178
<EOL>|179,180
Sulfonamides|180,192
/|193,194
Codeine|195,202
/|203,204
Bactrim|205,212
<EOL>|212,213
<EOL>|214,215
Attending|215,224
:|224,225
_|226,227
_|227,228
_|228,229
.|229,230
<EOL>|230,231
<EOL>|232,233
Chief|233,238
Complaint|239,248
:|248,249
<EOL>|249,250
abdominal|250,259
pain|260,264
and|265,268
vomiting|269,277
<EOL>|277,278
<EOL>|279,280
Major|280,285
Surgical|286,294
or|295,297
Invasive|298,306
Procedure|307,316
:|316,317
<EOL>|317,318
_|318,319
_|319,320
_|320,321
Exploratory|322,333
laparotomy|334,344
,|344,345
lysis|346,351
of|352,354
adhesions|355,364
,|364,365
small|366,371
<EOL>|371,372
bowel|372,377
resection|378,387
with|388,392
enteroenterostomy|393,410
.|410,411
<EOL>|411,412
<EOL>|412,413
<EOL>|414,415
History|415,422
of|423,425
Present|426,433
Illness|434,441
:|441,442
<EOL>|442,443
The|443,446
patient|447,454
is|455,457
a|458,459
_|460,461
_|461,462
_|462,463
year|464,468
old|469,472
woman|473,478
s|479,480
/|480,481
p|481,482
hysterectomy|483,495
for|496,499
uterine|500,507
<EOL>|508,509
fibroids|509,517
and|518,521
s|522,523
/|523,524
p|524,525
R|526,527
lung|528,532
resection|533,542
for|543,546
carcinoid|547,556
tumor|557,562
who|563,566
is|567,569
<EOL>|570,571
seen|571,575
in|576,578
surgical|579,587
consultation|588,600
for|601,604
abdominal|605,614
pain|615,619
,|619,620
nausea|621,627
,|627,628
and|629,632
<EOL>|633,634
vomiting|634,642
.|642,643
The|644,647
patient|648,655
was|656,659
feeling|660,667
well|668,672
until|673,678
early|679,684
this|685,689
morning|690,697
<EOL>|698,699
at|699,701
approximately|702,715
1|716,717
:|717,718
00am|718,722
,|722,723
when|724,728
she|729,732
developed|733,742
cramping|743,751
abdominal|752,761
<EOL>|762,763
pain|763,767
associated|768,778
with|779,783
nausea|784,790
and|791,794
bilious|795,802
emesis|803,809
without|810,817
blood|818,823
.|823,824
<EOL>|826,827
She|827,830
<EOL>|830,831
vomited|831,838
approximately|839,852
_|853,854
_|854,855
_|855,856
times|857,862
which|863,868
prompted|869,877
her|878,881
presentation|882,894
<EOL>|895,896
to|896,898
the|899,902
ED|903,905
.|905,906
At|908,910
the|911,914
time|915,919
of|920,922
her|923,926
emesis|927,933
,|933,934
she|935,938
had|939,942
diarrhea|943,951
and|952,955
<EOL>|956,957
moved|957,962
her|963,966
bowels|967,973
>|974,975
3|976,977
times|978,983
.|983,984
She|986,989
has|990,993
never|994,999
had|1000,1003
this|1004,1008
or|1009,1011
similar|1012,1019
<EOL>|1020,1021
pain|1021,1025
in|1026,1028
the|1029,1032
past|1033,1037
,|1037,1038
and|1039,1042
she|1043,1046
states|1047,1053
that|1054,1058
she|1059,1062
has|1063,1066
never|1067,1072
before|1073,1079
had|1080,1083
a|1084,1085
<EOL>|1086,1087
small|1087,1092
bowel|1093,1098
obstruction|1099,1110
.|1110,1111
She|1113,1116
has|1117,1120
never|1121,1126
had|1127,1130
a|1131,1132
colonoscopy|1133,1144
.|1144,1145
<EOL>|1146,1147
<EOL>|1147,1148
<EOL>|1149,1150
<EOL>|1150,1151
<EOL>|1152,1153
<EOL>|1153,1154
<EOL>|1155,1156
Past|1156,1160
Medical|1161,1168
History|1169,1176
:|1176,1177
<EOL>|1177,1178
PMH|1178,1181
:|1181,1182
<EOL>|1183,1184
carcinoid|1184,1193
tumor|1194,1199
as|1200,1202
above|1203,1208
<EOL>|1208,1209
Vitamin|1209,1216
B12|1217,1220
deficiency|1221,1231
<EOL>|1231,1232
depression|1232,1242
<EOL>|1242,1243
hyperlipidemia|1243,1257
<EOL>|1257,1258
<EOL>|1258,1259
PSH|1259,1262
:|1262,1263
<EOL>|1264,1265
s|1265,1266
/|1266,1267
p|1267,1268
R|1269,1270
lung|1271,1275
resection|1276,1285
in|1286,1288
_|1289,1290
_|1290,1291
_|1291,1292
at|1293,1295
_|1296,1297
_|1297,1298
_|1298,1299
<EOL>|1299,1300
s|1300,1301
/|1301,1302
p|1302,1303
hysterectomy|1304,1316
in|1317,1319
_|1320,1321
_|1321,1322
_|1322,1323
<EOL>|1323,1324
s|1324,1325
/|1325,1326
p|1326,1327
R|1328,1329
arm|1330,1333
surgery|1334,1341
<EOL>|1341,1342
<EOL>|1342,1343
<EOL>|1344,1345
Social|1345,1351
History|1352,1359
:|1359,1360
<EOL>|1360,1361
_|1361,1362
_|1362,1363
_|1363,1364
<EOL>|1364,1365
Family|1365,1371
History|1372,1379
:|1379,1380
<EOL>|1380,1381
non|1381,1384
contributory|1385,1397
<EOL>|1397,1398
<EOL>|1399,1400
Physical|1400,1408
Exam|1409,1413
:|1413,1414
<EOL>|1414,1415
Temp|1415,1419
96.9|1420,1424
HR|1426,1428
105|1429,1432
BP|1434,1436
108|1437,1440
/|1440,1441
92|1441,1443
100|1444,1447
%|1447,1448
RA|1448,1450
<EOL>|1450,1451
NAD|1451,1454
,|1454,1455
appears|1456,1463
non-toxic|1464,1473
but|1474,1477
uncomfortable|1478,1491
<EOL>|1491,1492
heart|1492,1497
tachycardic|1498,1509
but|1510,1513
regular|1514,1521
,|1521,1522
no|1523,1525
murmurs|1526,1533
appreciated|1534,1545
<EOL>|1545,1546
lungs|1546,1551
clear|1552,1557
to|1558,1560
auscultation|1561,1573
;|1573,1574
decreased|1575,1584
breath|1585,1591
sounds|1592,1598
on|1599,1601
R|1602,1603
;|1603,1604
<EOL>|1604,1605
well|1605,1609
-|1609,1610
healed|1610,1616
R|1617,1618
thoracotomy|1619,1630
scar|1631,1635
present|1636,1643
<EOL>|1643,1644
abdomen|1644,1651
soft|1652,1656
,|1656,1657
very|1658,1662
obese|1663,1668
,|1668,1669
minimally|1670,1679
distended|1680,1689
,|1689,1690
somewhat|1691,1699
tender|1700,1706
<EOL>|1707,1708
to|1708,1710
<EOL>|1710,1711
palpation|1711,1720
diffusely|1721,1730
across|1731,1737
abdomen|1738,1745
;|1745,1746
no|1747,1749
guarding|1750,1758
;|1758,1759
no|1760,1762
rebound|1763,1770
<EOL>|1770,1771
tenderness|1771,1781
,|1781,1782
low|1783,1786
midline|1787,1794
abdominal|1795,1804
wound|1805,1810
c|1811,1812
/|1812,1813
d|1813,1814
/|1814,1815
i|1815,1816
,|1816,1817
no|1818,1820
drainage|1821,1829
,|1829,1830
no|1831,1833
<EOL>|1834,1835
erythema|1835,1843
<EOL>|1843,1844
<EOL>|1844,1845
<EOL>|1846,1847
Pertinent|1847,1856
Results|1857,1864
:|1864,1865
<EOL>|1865,1866
_|1866,1867
_|1867,1868
_|1868,1869
04|1870,1872
:|1872,1873
40AM|1873,1877
WBC|1880,1883
-|1883,1884
12|1884,1886
.|1886,1887
5|1887,1888
*|1888,1889
#|1889,1890
RBC|1891,1894
-|1894,1895
4|1895,1896
.|1896,1897
46|1897,1899
HGB|1900,1903
-|1903,1904
13.6|1904,1908
HCT|1909,1912
-|1912,1913
39.7|1913,1917
MCV|1918,1921
-|1921,1922
89|1922,1924
<EOL>|1925,1926
MCH|1926,1929
-|1929,1930
30.5|1930,1934
MCHC|1935,1939
-|1939,1940
34.2|1940,1944
RDW|1945,1948
-|1948,1949
13.0|1949,1953
<EOL>|1953,1954
_|1954,1955
_|1955,1956
_|1956,1957
04|1958,1960
:|1960,1961
40AM|1961,1965
NEUTS|1968,1973
-|1973,1974
91|1974,1976
.|1976,1977
1|1977,1978
*|1978,1979
LYMPHS|1980,1986
-|1986,1987
7|1987,1988
.|1988,1989
4|1989,1990
*|1990,1991
MONOS|1992,1997
-|1997,1998
0|1998,1999
.|1999,2000
8|2000,2001
*|2001,2002
EOS|2003,2006
-|2006,2007
0.3|2007,2010
<EOL>|2011,2012
BASOS|2012,2017
-|2017,2018
0.2|2018,2021
<EOL>|2021,2022
_|2022,2023
_|2023,2024
_|2024,2025
04|2026,2028
:|2028,2029
40AM|2029,2033
PLT|2036,2039
COUNT|2040,2045
-|2045,2046
329|2046,2049
<EOL>|2049,2050
_|2050,2051
_|2051,2052
_|2052,2053
04|2054,2056
:|2056,2057
40AM|2057,2061
GLUCOSE|2064,2071
-|2071,2072
151|2072,2075
*|2075,2076
UREA|2077,2081
N|2082,2083
-|2083,2084
10|2084,2086
CREAT|2087,2092
-|2092,2093
0.8|2093,2096
SODIUM|2097,2103
-|2103,2104
142|2104,2107
<EOL>|2108,2109
POTASSIUM|2109,2118
-|2118,2119
3.8|2119,2122
CHLORIDE|2123,2131
-|2131,2132
105|2132,2135
TOTAL|2136,2141
CO2|2142,2145
-|2145,2146
28|2146,2148
ANION|2149,2154
GAP|2155,2158
-|2158,2159
13|2159,2161
<EOL>|2161,2162
_|2162,2163
_|2163,2164
_|2164,2165
04|2166,2168
:|2168,2169
40AM|2169,2173
ALT|2176,2179
(|2179,2180
SGPT|2180,2184
)|2184,2185
-|2185,2186
12|2186,2188
AST|2189,2192
(|2192,2193
SGOT|2193,2197
)|2197,2198
-|2198,2199
16|2199,2201
LD|2202,2204
(|2204,2205
LDH|2205,2208
)|2208,2209
-|2209,2210
180|2210,2213
ALK|2214,2217
<EOL>|2218,2219
PHOS|2219,2223
-|2223,2224
62|2224,2226
<EOL>|2227,2228
<EOL>|2228,2229
_|2229,2230
_|2230,2231
_|2231,2232
CT|2233,2235
of|2236,2238
abdomen|2239,2246
and|2247,2250
pelvis|2251,2257
:|2258,2259
1|2259,2260
.|2260,2261
Slightly|2262,2270
dilated|2271,2278
loops|2279,2284
of|2285,2287
<EOL>|2288,2289
small|2289,2294
bowel|2295,2300
with|2301,2305
fecalization|2306,2318
of|2319,2321
small|2322,2327
bowel|2328,2333
contents|2334,2342
and|2343,2346
distal|2347,2353
<EOL>|2354,2355
collapsed|2355,2364
loops|2365,2370
,|2370,2371
together|2372,2380
indicating|2381,2391
early|2392,2397
complete|2398,2406
or|2407,2409
partial|2410,2417
<EOL>|2418,2419
small|2419,2424
-|2424,2425
bowel|2425,2430
obstruction|2431,2442
.|2442,2443
<EOL>|2444,2445
2.|2445,2447
Post-surgical|2448,2461
changes|2462,2469
noted|2470,2475
at|2476,2478
the|2479,2482
right|2483,2488
ribs|2489,2493
as|2494,2496
detailed|2497,2505
<EOL>|2506,2507
above|2507,2512
.|2512,2513
<EOL>|2513,2514
<EOL>|2514,2515
_|2515,2516
_|2516,2517
_|2517,2518
CT|2519,2521
of|2522,2524
abdoman|2525,2532
and|2533,2536
pelvis|2537,2543
:|2544,2545
<EOL>|2547,2548
1.|2548,2550
Interval|2551,2559
worsening|2560,2569
of|2570,2572
small|2573,2578
bowel|2579,2584
obstruction|2585,2596
.|2596,2597
Transition|2598,2608
<EOL>|2609,2610
point|2610,2615
in|2616,2618
the|2619,2622
<EOL>|2623,2624
left|2624,2628
mid|2629,2632
abdomen.|2633,2641
(|2642,2643
The|2643,2646
patient|2647,2654
went|2655,2659
to|2660,2662
the|2663,2666
OR|2667,2669
on|2670,2672
the|2673,2676
evening|2677,2684
of|2685,2687
<EOL>|2688,2689
the|2689,2692
study|2693,2698
)|2698,2699
.|2699,2700
<EOL>|2701,2702
2.|2702,2704
Trace|2705,2710
free|2711,2715
fluid|2716,2721
in|2722,2724
the|2725,2728
pelvis|2729,2735
is|2736,2738
likely|2739,2745
physiologic|2746,2757
.|2757,2758
<EOL>|2760,2761
<EOL>|2761,2762
<EOL>|2764,2765
<EOL>|2765,2766
_|2766,2767
_|2767,2768
_|2768,2769
10|2770,2772
:|2772,2773
57PM|2773,2777
URINE|2778,2783
COLOR|2785,2790
-|2790,2791
Yellow|2791,2797
APPEAR|2798,2804
-|2804,2805
Hazy|2805,2809
SP|2810,2812
_|2813,2814
_|2814,2815
_|2815,2816
<EOL>|2816,2817
_|2817,2818
_|2818,2819
_|2819,2820
10|2821,2823
:|2823,2824
57PM|2824,2828
URINE|2829,2834
BLOOD|2836,2841
-|2841,2842
LG|2842,2844
NITRITE|2845,2852
-|2852,2853
NEG|2853,2856
PROTEIN|2857,2864
-|2864,2865
TR|2865,2867
<EOL>|2868,2869
GLUCOSE|2869,2876
-|2876,2877
NEG|2877,2880
KETONE|2881,2887
-|2887,2888
15|2888,2890
BILIRUBIN|2891,2900
-|2900,2901
NEG|2901,2904
UROBILNGN|2905,2914
-|2914,2915
NEG|2915,2918
PH|2919,2921
-|2921,2922
6.5|2922,2925
<EOL>|2926,2927
LEUK|2927,2931
-|2931,2932
NEG|2932,2935
<EOL>|2935,2936
_|2936,2937
_|2937,2938
_|2938,2939
10|2940,2942
:|2942,2943
57PM|2943,2947
URINE|2948,2953
RBC|2955,2958
-|2958,2959
>|2959,2960
50|2960,2962
_|2963,2964
_|2964,2965
_|2965,2966
BACTERIA|2967,2975
-|2975,2976
MOD|2976,2979
YEAST|2980,2985
-|2985,2986
NONE|2986,2990
<EOL>|2991,2992
EPI|2992,2995
-|2995,2996
0|2996,2997
<EOL>|2997,2998
_|2998,2999
_|2999,3000
_|3000,3001
10|3002,3004
:|3004,3005
57PM|3005,3009
URINE|3010,3015
MUCOUS|3017,3023
-|3023,3024
OCC|3024,3027
<EOL>|3027,3028
_|3028,3029
_|3029,3030
_|3030,3031
04|3032,3034
:|3034,3035
40AM|3035,3039
GLUCOSE|3042,3049
-|3049,3050
151|3050,3053
*|3053,3054
UREA|3055,3059
N|3060,3061
-|3061,3062
10|3062,3064
CREAT|3065,3070
-|3070,3071
0.8|3071,3074
SODIUM|3075,3081
-|3081,3082
142|3082,3085
<EOL>|3086,3087
POTASSIUM|3087,3096
-|3096,3097
3.8|3097,3100
CHLORIDE|3101,3109
-|3109,3110
105|3110,3113
TOTAL|3114,3119
CO2|3120,3123
-|3123,3124
28|3124,3126
ANION|3127,3132
GAP|3133,3136
-|3136,3137
13|3137,3139
<EOL>|3139,3140
_|3140,3141
_|3141,3142
_|3142,3143
04|3144,3146
:|3146,3147
40AM|3147,3151
estGFR|3154,3160
-|3160,3161
Using|3161,3166
this|3167,3171
<EOL>|3171,3172
_|3172,3173
_|3173,3174
_|3174,3175
04|3176,3178
:|3178,3179
40AM|3179,3183
ALT|3186,3189
(|3189,3190
SGPT|3190,3194
)|3194,3195
-|3195,3196
12|3196,3198
AST|3199,3202
(|3202,3203
SGOT|3203,3207
)|3207,3208
-|3208,3209
16|3209,3211
LD|3212,3214
(|3214,3215
LDH|3215,3218
)|3218,3219
-|3219,3220
180|3220,3223
ALK|3224,3227
<EOL>|3228,3229
PHOS|3229,3233
-|3233,3234
62|3234,3236
TOT|3237,3240
BILI|3241,3245
-|3245,3246
0.2|3246,3249
<EOL>|3249,3250
_|3250,3251
_|3251,3252
_|3252,3253
04|3254,3256
:|3256,3257
40AM|3257,3261
LIPASE|3264,3270
-|3270,3271
17|3271,3273
<EOL>|3273,3274
_|3274,3275
_|3275,3276
_|3276,3277
04|3278,3280
:|3280,3281
40AM|3281,3285
WBC|3288,3291
-|3291,3292
12|3292,3294
.|3294,3295
5|3295,3296
*|3296,3297
#|3297,3298
RBC|3299,3302
-|3302,3303
4|3303,3304
.|3304,3305
46|3305,3307
HGB|3308,3311
-|3311,3312
13.6|3312,3316
HCT|3317,3320
-|3320,3321
39.7|3321,3325
MCV|3326,3329
-|3329,3330
89|3330,3332
<EOL>|3333,3334
MCH|3334,3337
-|3337,3338
30.5|3338,3342
MCHC|3343,3347
-|3347,3348
34.2|3348,3352
RDW|3353,3356
-|3356,3357
13.0|3357,3361
<EOL>|3361,3362
_|3362,3363
_|3363,3364
_|3364,3365
04|3366,3368
:|3368,3369
40AM|3369,3373
NEUTS|3376,3381
-|3381,3382
91|3382,3384
.|3384,3385
1|3385,3386
*|3386,3387
LYMPHS|3388,3394
-|3394,3395
7|3395,3396
.|3396,3397
4|3397,3398
*|3398,3399
MONOS|3400,3405
-|3405,3406
0|3406,3407
.|3407,3408
8|3408,3409
*|3409,3410
EOS|3411,3414
-|3414,3415
0.3|3415,3418
<EOL>|3419,3420
BASOS|3420,3425
-|3425,3426
0.2|3426,3429
<EOL>|3429,3430
_|3430,3431
_|3431,3432
_|3432,3433
04|3434,3436
:|3436,3437
40AM|3437,3441
PLT|3444,3447
COUNT|3448,3453
-|3453,3454
329|3454,3457
<EOL>|3457,3458
<EOL>|3459,3460
Brief|3460,3465
Hospital|3466,3474
Course|3475,3481
:|3481,3482
<EOL>|3482,3483
This|3483,3487
_|3488,3489
_|3489,3490
_|3490,3491
year|3492,3496
old|3497,3500
female|3501,3507
was|3508,3511
admitted|3512,3520
to|3521,3523
the|3524,3527
hospital|3528,3536
and|3537,3540
was|3541,3544
<EOL>|3545,3546
made|3546,3550
NPO|3551,3554
,|3554,3555
IV|3556,3558
fluids|3559,3565
were|3566,3570
started|3571,3578
and|3579,3582
she|3583,3586
had|3587,3590
a|3591,3592
nasogastric|3593,3604
tube|3605,3609
<EOL>|3610,3611
placed|3611,3617
.|3617,3618
She|3620,3623
was|3624,3627
pan|3628,3631
cultured|3632,3640
for|3641,3644
a|3645,3646
temperature|3647,3658
of|3659,3661
101|3662,3665
and|3666,3669
was|3670,3673
<EOL>|3674,3675
followed|3675,3683
with|3684,3688
serial|3689,3695
KUB|3696,3699
's|3699,3701
and|3702,3705
physical|3706,3714
exam|3715,3719
.|3719,3720
Her|3721,3724
nasogastric|3725,3736
<EOL>|3737,3738
tube|3738,3742
was|3743,3746
clamped|3747,3754
on|3755,3757
hospital|3758,3766
day|3767,3770
2|3771,3772
and|3773,3776
she|3777,3780
soon|3781,3785
developed|3786,3795
<EOL>|3796,3797
increased|3797,3806
abdominal|3807,3816
pain|3817,3821
prompting|3822,3831
repeat|3832,3838
CT|3839,3841
of|3842,3844
abdomen|3845,3852
and|3853,3856
<EOL>|3857,3858
pelvis|3858,3864
.|3864,3865
This|3867,3871
demonstrated|3872,3884
an|3885,3887
increase|3888,3896
in|3897,3899
the|3900,3903
degree|3904,3910
of|3911,3913
<EOL>|3914,3915
obstruction|3915,3926
and|3927,3930
she|3931,3934
was|3935,3938
subsequently|3939,3951
taken|3952,3957
to|3958,3960
the|3961,3964
operating|3965,3974
room|3975,3979
<EOL>|3980,3981
for|3981,3984
the|3985,3988
aforementioned|3989,4003
procedure|4004,4013
.|4013,4014
<EOL>|4014,4015
<EOL>|4015,4016
She|4016,4019
tolerated|4020,4029
the|4030,4033
procedure|4034,4043
well|4044,4048
,|4048,4049
remained|4050,4058
NPO|4059,4062
with|4064,4068
nasogastric|4069,4080
<EOL>|4081,4082
tube|4082,4086
in|4087,4089
place|4090,4095
and|4096,4099
treated|4100,4107
with|4108,4112
IV|4113,4115
fluids|4116,4122
.|4122,4123
Her|4125,4128
pain|4129,4133
was|4134,4137
<EOL>|4138,4139
initially|4139,4148
controlled|4149,4159
with|4160,4164
a|4165,4166
morphine|4167,4175
PCA|4176,4179
.|4180,4181
Her|4183,4186
nasogastric|4187,4198
tube|4199,4203
<EOL>|4204,4205
was|4205,4208
removed|4209,4216
on|4217,4219
post|4220,4224
op|4225,4227
day|4228,4231
#|4232,4233
2|4233,4234
and|4235,4238
she|4239,4242
began|4243,4248
a|4249,4250
clear|4251,4256
liquid|4257,4263
diet|4264,4268
<EOL>|4269,4270
which|4270,4275
she|4276,4279
tolerated|4280,4289
well|4290,4294
.|4294,4295
This|4297,4301
was|4302,4305
gradually|4306,4315
advanced|4316,4324
over|4325,4329
36|4330,4332
<EOL>|4333,4334
hours|4334,4339
to|4340,4342
a|4343,4344
regular|4345,4352
diet|4353,4357
and|4358,4361
was|4362,4365
tolerated|4366,4375
well|4376,4380
.|4380,4381
She|4383,4386
was|4387,4390
having|4391,4397
<EOL>|4398,4399
bowel|4399,4404
movements|4405,4414
and|4415,4418
tolerated|4419,4428
oral|4429,4433
pain|4434,4438
medication|4439,4449
.|4449,4450
Her|4452,4455
<EOL>|4456,4457
incision|4457,4465
was|4466,4469
healing|4470,4477
well|4478,4482
and|4483,4486
staples|4487,4494
were|4495,4499
intact|4500,4506
.|4506,4507
After|4509,4514
an|4515,4517
<EOL>|4518,4519
uncomplicated|4519,4532
course|4533,4539
she|4540,4543
was|4544,4547
discharged|4548,4558
home|4559,4563
on|4564,4566
_|4567,4568
_|4568,4569
_|4569,4570
<EOL>|4570,4571
<EOL>|4572,4573
Medications|4573,4584
on|4585,4587
Admission|4588,4597
:|4597,4598
<EOL>|4598,4599
Albuteral|4599,4608
MDI|4609,4612
prn|4613,4616
wheezes|4617,4624
<EOL>|4624,4625
Flovent|4625,4632
inhaler|4633,4640
prn|4641,4644
wheezes|4645,4652
<EOL>|4652,4653
Srtraline|4653,4662
200|4663,4666
mg|4667,4669
oral|4670,4674
daily|4675,4680
<EOL>|4680,4681
Simvastatin|4681,4692
20|4693,4695
mg|4696,4698
oral|4699,4703
daily|4704,4709
<EOL>|4709,4710
Trazadone|4710,4719
100|4720,4723
mg|4724,4726
oral|4727,4731
daily|4732,4737
at|4738,4740
bedtime|4741,4748
<EOL>|4748,4749
Wellbutrin|4749,4759
75|4760,4762
mg|4763,4765
oral|4766,4770
twice|4771,4776
a|4777,4778
day|4779,4782
<EOL>|4782,4783
<EOL>|4784,4785
Discharge|4785,4794
Medications|4795,4806
:|4806,4807
<EOL>|4807,4808
1.|4808,4810
Albuterol|4811,4820
Sulfate|4821,4828
90|4829,4831
mcg|4832,4835
/|4835,4836
Actuation|4836,4845
HFA|4846,4849
Aerosol|4850,4857
Inhaler|4858,4865
Sig|4866,4869
:|4869,4870
<EOL>|4871,4872
Two|4872,4875
(|4876,4877
2|4877,4878
)|4878,4879
Puff|4880,4884
Inhalation|4885,4895
Q6H|4896,4899
(|4900,4901
every|4901,4906
6|4907,4908
hours|4909,4914
)|4914,4915
as|4916,4918
needed|4919,4925
for|4926,4929
<EOL>|4930,4931
wheezing|4931,4939
,|4939,4940
shortness|4941,4950
of|4951,4953
breath|4954,4960
.|4960,4961
<EOL>|4963,4964
2.|4964,4966
Fluticasone|4967,4978
110|4979,4982
mcg|4983,4986
/|4986,4987
Actuation|4987,4996
Aerosol|4997,5004
Sig|5005,5008
:|5008,5009
Two|5010,5013
(|5014,5015
2|5015,5016
)|5016,5017
Puff|5018,5022
<EOL>|5023,5024
Inhalation|5024,5034
BID|5035,5038
(|5039,5040
2|5040,5041
times|5042,5047
a|5048,5049
day|5050,5053
)|5053,5054
.|5054,5055
<EOL>|5057,5058
3.|5058,5060
Oxycodone|5061,5070
-|5070,5071
Acetaminophen|5071,5084
_|5085,5086
_|5086,5087
_|5087,5088
mg|5089,5091
Tablet|5092,5098
Sig|5099,5102
:|5102,5103
_|5104,5105
_|5105,5106
_|5106,5107
Tablets|5108,5115
PO|5116,5118
<EOL>|5119,5120
Q4H|5120,5123
(|5124,5125
every|5125,5130
4|5131,5132
hours|5133,5138
)|5138,5139
as|5140,5142
needed|5143,5149
for|5150,5153
pain|5154,5158
.|5158,5159
<EOL>|5159,5160
Disp|5160,5164
:|5164,5165
*|5165,5166
40|5166,5168
Tablet|5169,5175
(|5175,5176
s|5176,5177
)|5177,5178
*|5178,5179
Refills|5180,5187
:|5187,5188
*|5188,5189
0|5189,5190
*|5190,5191
<EOL>|5191,5192
4.|5192,5194
Docusate|5195,5203
Sodium|5204,5210
100|5211,5214
mg|5215,5217
Capsule|5218,5225
Sig|5226,5229
:|5229,5230
One|5231,5234
(|5235,5236
1|5236,5237
)|5237,5238
Capsule|5239,5246
PO|5247,5249
BID|5250,5253
(|5254,5255
2|5255,5256
<EOL>|5257,5258
times|5258,5263
a|5264,5265
day|5266,5269
)|5269,5270
.|5270,5271
<EOL>|5271,5272
Disp|5272,5276
:|5276,5277
*|5277,5278
60|5278,5280
Capsule|5281,5288
(|5288,5289
s|5289,5290
)|5290,5291
*|5291,5292
Refills|5293,5300
:|5300,5301
*|5301,5302
2|5302,5303
*|5303,5304
<EOL>|5304,5305
5.|5305,5307
Simvastatin|5308,5319
20|5320,5322
mg|5323,5325
Tablet|5326,5332
Sig|5333,5336
:|5336,5337
One|5338,5341
(|5342,5343
1|5343,5344
)|5344,5345
Tablet|5346,5352
PO|5353,5355
once|5356,5360
a|5361,5362
day|5363,5366
.|5366,5367
<EOL>|5367,5368
Disp|5368,5372
:|5372,5373
*|5373,5374
30|5374,5376
Tablet|5377,5383
(|5383,5384
s|5384,5385
)|5385,5386
*|5386,5387
Refills|5388,5395
:|5395,5396
*|5396,5397
2|5397,5398
*|5398,5399
<EOL>|5399,5400
6.|5400,5402
Trazodone|5403,5412
100|5413,5416
mg|5417,5419
Tablet|5420,5426
Sig|5427,5430
:|5430,5431
One|5432,5435
(|5436,5437
1|5437,5438
)|5438,5439
Tablet|5440,5446
PO|5447,5449
at|5450,5452
bedtime|5453,5460
.|5460,5461
<EOL>|5463,5464
7.|5464,5466
Wellbutrin|5467,5477
75|5478,5480
mg|5481,5483
Tablet|5484,5490
Sig|5491,5494
:|5494,5495
One|5496,5499
(|5500,5501
1|5501,5502
)|5502,5503
Tablet|5504,5510
PO|5511,5513
twice|5514,5519
a|5520,5521
day|5522,5525
.|5525,5526
<EOL>|5528,5529
<EOL>|5529,5530
<EOL>|5531,5532
Discharge|5532,5541
Disposition|5542,5553
:|5553,5554
<EOL>|5554,5555
Home|5555,5559
<EOL>|5559,5560
<EOL>|5561,5562
Discharge|5562,5571
Diagnosis|5572,5581
:|5581,5582
<EOL>|5582,5583
High|5583,5587
grade|5588,5593
small|5594,5599
bowel|5600,5605
obstruction|5606,5617
<EOL>|5617,5618
<EOL>|5618,5619
<EOL>|5620,5621
Discharge|5621,5630
Condition|5631,5640
:|5640,5641
<EOL>|5641,5642
Henodynamically|5642,5657
stable|5658,5664
,|5664,5665
tolerating|5666,5676
a|5677,5678
regular|5679,5686
diet|5687,5691
,|5691,5692
having|5693,5699
bowel|5700,5705
<EOL>|5706,5707
movements|5707,5716
,|5716,5717
adequate|5718,5726
pain|5727,5731
control|5732,5739
<EOL>|5739,5740
<EOL>|5740,5741
<EOL>|5742,5743
Discharge|5743,5752
Instructions|5753,5765
:|5765,5766
<EOL>|5766,5767
Please|5767,5773
call|5774,5778
your|5779,5783
doctor|5784,5790
or|5791,5793
nurse|5794,5799
practitioner|5800,5812
or|5813,5815
return|5816,5822
to|5823,5825
the|5826,5829
<EOL>|5830,5831
Emergency|5831,5840
Department|5841,5851
for|5852,5855
any|5856,5859
of|5860,5862
the|5863,5866
following|5867,5876
:|5876,5877
<EOL>|5877,5878
<EOL>|5878,5879
*|5879,5880
You|5880,5883
experience|5884,5894
new|5895,5898
chest|5899,5904
pain|5905,5909
,|5909,5910
pressure|5911,5919
,|5919,5920
squeezing|5921,5930
or|5931,5933
<EOL>|5934,5935
tightness|5935,5944
.|5944,5945
<EOL>|5945,5946
<EOL>|5946,5947
*|5947,5948
New|5948,5951
or|5952,5954
worsening|5955,5964
cough|5965,5970
,|5970,5971
shortness|5972,5981
of|5982,5984
breath|5985,5991
,|5991,5992
or|5993,5995
wheeze|5996,6002
.|6002,6003
<EOL>|6003,6004
<EOL>|6004,6005
*|6005,6006
If|6006,6008
you|6009,6012
are|6013,6016
vomiting|6017,6025
and|6026,6029
can|6030,6033
not|6033,6036
keep|6037,6041
down|6042,6046
fluids|6047,6053
or|6054,6056
your|6057,6061
<EOL>|6062,6063
medications|6063,6074
.|6074,6075
<EOL>|6075,6076
<EOL>|6076,6077
*|6077,6078
You|6078,6081
are|6082,6085
getting|6086,6093
dehydrated|6094,6104
due|6105,6108
to|6109,6111
continued|6112,6121
vomiting|6122,6130
,|6130,6131
diarrhea|6132,6140
,|6140,6141
<EOL>|6142,6143
or|6143,6145
other|6146,6151
reasons|6152,6159
.|6159,6160
Signs|6161,6166
of|6167,6169
dehydration|6170,6181
include|6182,6189
dry|6190,6193
mouth|6194,6199
,|6199,6200
rapid|6201,6206
<EOL>|6207,6208
heartbeat|6208,6217
,|6217,6218
or|6219,6221
feeling|6222,6229
dizzy|6230,6235
or|6236,6238
faint|6239,6244
when|6245,6249
standing|6250,6258
.|6258,6259
<EOL>|6259,6260
<EOL>|6260,6261
*|6261,6262
You|6262,6265
see|6266,6269
blood|6270,6275
or|6276,6278
dark|6279,6283
/|6283,6284
black|6284,6289
material|6290,6298
when|6299,6303
you|6304,6307
vomit|6308,6313
or|6314,6316
have|6317,6321
a|6322,6323
<EOL>|6324,6325
bowel|6325,6330
movement|6331,6339
.|6339,6340
<EOL>|6340,6341
<EOL>|6341,6342
*|6342,6343
You|6343,6346
experience|6347,6357
burning|6358,6365
when|6366,6370
you|6371,6374
urinate|6375,6382
,|6382,6383
have|6384,6388
blood|6389,6394
in|6395,6397
your|6398,6402
<EOL>|6403,6404
urine|6404,6409
,|6409,6410
or|6411,6413
experience|6414,6424
a|6425,6426
discharge|6427,6436
.|6436,6437
<EOL>|6437,6438
<EOL>|6438,6439
*|6439,6440
Your|6440,6444
pain|6445,6449
in|6450,6452
not|6453,6456
improving|6457,6466
within|6467,6473
_|6474,6475
_|6475,6476
_|6476,6477
hours|6478,6483
or|6484,6486
is|6487,6489
not|6490,6493
gone|6494,6498
<EOL>|6499,6500
within|6500,6506
24|6507,6509
hours|6510,6515
.|6515,6516
Call|6517,6521
or|6522,6524
return|6525,6531
immediately|6532,6543
if|6544,6546
your|6547,6551
pain|6552,6556
is|6557,6559
<EOL>|6560,6561
getting|6561,6568
worse|6569,6574
or|6575,6577
changes|6578,6585
location|6586,6594
or|6595,6597
moving|6598,6604
to|6605,6607
your|6608,6612
chest|6613,6618
or|6619,6621
<EOL>|6622,6623
back|6623,6627
.|6627,6628
<EOL>|6628,6629
<EOL>|6629,6630
*|6630,6631
You|6631,6634
have|6635,6639
shaking|6640,6647
chills|6648,6654
,|6654,6655
or|6656,6658
fever|6659,6664
greater|6665,6672
than|6673,6677
101.5|6678,6683
degrees|6684,6691
<EOL>|6692,6693
Fahrenheit|6693,6703
or|6704,6706
38|6707,6709
degrees|6710,6717
Celsius|6718,6725
.|6725,6726
<EOL>|6726,6727
<EOL>|6727,6728
*|6728,6729
Any|6729,6732
change|6733,6739
in|6740,6742
your|6743,6747
symptoms|6748,6756
,|6756,6757
or|6758,6760
any|6761,6764
new|6765,6768
symptoms|6769,6777
that|6778,6782
concern|6783,6790
<EOL>|6791,6792
you|6792,6795
.|6795,6796
<EOL>|6796,6797
<EOL>|6797,6798
Please|6798,6804
resume|6805,6811
all|6812,6815
regular|6816,6823
home|6824,6828
medications|6829,6840
,|6841,6842
unless|6843,6849
specifically|6850,6862
<EOL>|6863,6864
advised|6864,6871
not|6872,6875
to|6876,6878
take|6879,6883
a|6884,6885
particular|6886,6896
medication|6897,6907
.|6907,6908
Also|6909,6913
,|6913,6914
please|6915,6921
take|6922,6926
<EOL>|6927,6928
any|6928,6931
new|6932,6935
medications|6936,6947
as|6948,6950
prescribed|6951,6961
.|6961,6962
<EOL>|6962,6963
<EOL>|6963,6964
Please|6964,6970
get|6971,6974
plenty|6975,6981
of|6982,6984
rest|6985,6989
,|6989,6990
continue|6991,6999
to|7000,7002
ambulate|7003,7011
several|7012,7019
times|7020,7025
<EOL>|7026,7027
per|7027,7030
day|7031,7034
,|7034,7035
and|7036,7039
drink|7040,7045
adequate|7046,7054
amounts|7055,7062
of|7063,7065
fluids|7066,7072
.|7072,7073
Avoid|7074,7079
lifting|7080,7087
<EOL>|7088,7089
weights|7089,7096
greater|7097,7104
than|7105,7109
_|7110,7111
_|7111,7112
_|7112,7113
lbs|7114,7117
until|7118,7123
you|7124,7127
follow|7128,7134
-|7134,7135
up|7135,7137
with|7138,7142
your|7143,7147
<EOL>|7148,7149
surgeon|7149,7156
.|7156,7157
<EOL>|7157,7158
<EOL>|7158,7159
Avoid|7159,7164
driving|7165,7172
or|7173,7175
operating|7176,7185
heavy|7186,7191
machinery|7192,7201
while|7202,7207
taking|7208,7214
pain|7215,7219
<EOL>|7220,7221
medications|7221,7232
.|7232,7233
<EOL>|7233,7234
<EOL>|7234,7235
Incision|7235,7243
Care|7244,7248
:|7248,7249
<EOL>|7249,7250
<EOL>|7250,7251
*|7251,7252
Please|7252,7258
call|7259,7263
your|7264,7268
doctor|7269,7275
or|7276,7278
nurse|7279,7284
practitioner|7285,7297
if|7298,7300
you|7301,7304
have|7305,7309
<EOL>|7310,7311
increased|7311,7320
pain|7321,7325
,|7325,7326
swelling|7327,7335
,|7335,7336
redness|7337,7344
,|7344,7345
or|7346,7348
drainage|7349,7357
from|7358,7362
the|7363,7366
incision|7367,7375
<EOL>|7376,7377
site|7377,7381
.|7381,7382
<EOL>|7382,7383
<EOL>|7383,7384
*|7384,7385
Avoid|7385,7390
swimming|7391,7399
and|7400,7403
baths|7404,7409
until|7410,7415
your|7416,7420
follow|7421,7427
-|7427,7428
up|7428,7430
appointment|7431,7442
.|7442,7443
<EOL>|7443,7444
<EOL>|7444,7445
*|7445,7446
You|7446,7449
may|7450,7453
shower|7454,7460
,|7460,7461
and|7462,7465
wash|7466,7470
surgical|7471,7479
incisions|7480,7489
with|7490,7494
a|7495,7496
mild|7497,7501
soap|7502,7506
<EOL>|7507,7508
and|7508,7511
warm|7512,7516
water|7517,7522
.|7522,7523
Gently|7524,7530
pat|7531,7534
the|7535,7538
area|7539,7543
dry|7544,7547
.|7547,7548
<EOL>|7548,7549
<EOL>|7549,7550
*|7550,7551
If|7551,7553
you|7554,7557
have|7558,7562
staples|7563,7570
,|7570,7571
they|7572,7576
will|7577,7581
be|7582,7584
removed|7585,7592
at|7593,7595
your|7596,7600
follow|7601,7607
-|7607,7608
up|7608,7610
<EOL>|7611,7612
appointment|7612,7623
.|7623,7624
<EOL>|7624,7625
<EOL>|7625,7626
*|7626,7627
If|7627,7629
you|7630,7633
have|7634,7638
steri|7639,7644
-|7644,7645
strips|7645,7651
,|7651,7652
they|7653,7657
will|7658,7662
fall|7663,7667
off|7668,7671
on|7672,7674
their|7675,7680
own|7681,7684
.|7684,7685
<EOL>|7686,7687
Please|7687,7693
remove|7694,7700
any|7701,7704
remaining|7705,7714
strips|7715,7721
_|7722,7723
_|7723,7724
_|7724,7725
days|7726,7730
after|7731,7736
surgery|7737,7744
.|7744,7745
<EOL>|7745,7746
<EOL>|7746,7747
*|7747,7748
Please|7748,7754
look|7755,7759
at|7760,7762
the|7763,7766
site|7767,7771
every|7772,7777
day|7778,7781
for|7782,7785
signs|7786,7791
of|7792,7794
infection|7795,7804
<EOL>|7805,7806
(|7806,7807
increased|7807,7816
redness|7817,7824
or|7825,7827
pain|7828,7832
,|7832,7833
swelling|7834,7842
,|7842,7843
odor|7844,7848
,|7848,7849
yellow|7850,7856
or|7857,7859
bloody|7860,7866
<EOL>|7867,7868
<EOL>|7868,7869
<EOL>|7870,7871
Followup|7871,7879
Instructions|7880,7892
:|7892,7893
<EOL>|7893,7894
_|7894,7895
_|7895,7896
_|7896,7897
<EOL>|7897,7898

