 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|152,162|false|false|false|||OBSTETRICS
Procedure|Health Care Activity|SIMPLE_SEGMENT|152,162|false|false|false|C0587597|Obstetrics service|OBSTETRICS
Event|Event|SIMPLE_SEGMENT|163,173|false|false|false|||GYNECOLOGY
Drug|Organic Chemical|Allergies|188,195|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|188,195|false|false|false|C0009214|codeine|Codeine
Event|Event|Allergies|188,195|false|false|false|||Codeine
Drug|Organic Chemical|Allergies|198,208|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Allergies|198,208|false|false|false|C0060926|gabapentin|gabapentin
Event|Event|Allergies|198,208|false|false|false|||gabapentin
Drug|Organic Chemical|Allergies|211,219|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|Allergies|211,219|false|false|false|C0026549|morphine|morphine
Event|Event|Allergies|211,219|false|false|false|||morphine
Drug|Antibiotic|Allergies|222,233|false|false|false|C0002645|amoxicillin|Amoxicillin
Drug|Organic Chemical|Allergies|222,233|false|false|false|C0002645|amoxicillin|Amoxicillin
Event|Event|Allergies|222,233|false|false|false|||Amoxicillin
Drug|Organic Chemical|Allergies|236,249|false|false|false|C0025872|metronidazole|metronidazole
Drug|Pharmacologic Substance|Allergies|236,249|false|false|false|C0025872|metronidazole|metronidazole
Event|Event|Allergies|236,249|false|false|false|||metronidazole
Drug|Organic Chemical|Allergies|253,265|false|false|false|C0033493|propoxyphene|propoxyphene
Drug|Pharmacologic Substance|Allergies|253,265|false|false|false|C0033493|propoxyphene|propoxyphene
Event|Event|Allergies|253,265|false|false|false|||propoxyphene
Procedure|Laboratory Procedure|Allergies|253,265|false|false|false|C0202458|Propoxyphene measurement|propoxyphene
Drug|Organic Chemical|Allergies|268,277|false|false|false|C0762662|rofecoxib|rofecoxib
Drug|Pharmacologic Substance|Allergies|268,277|false|false|false|C0762662|rofecoxib|rofecoxib
Event|Event|Allergies|268,277|false|false|false|||rofecoxib
Drug|Organic Chemical|Allergies|280,288|false|false|false|C0591750|Macrobid|Macrobid
Drug|Pharmacologic Substance|Allergies|280,288|false|false|false|C0591750|Macrobid|Macrobid
Event|Event|Allergies|280,288|false|false|false|||Macrobid
Drug|Organic Chemical|Allergies|291,301|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Allergies|291,301|false|false|false|C0016860|furosemide|furosemide
Event|Event|Allergies|291,301|false|false|false|||furosemide
Drug|Organic Chemical|Allergies|304,311|false|false|false|C1699150|Amitiza|Amitiza
Drug|Pharmacologic Substance|Allergies|304,311|false|false|false|C1699150|Amitiza|Amitiza
Drug|Pharmacologic Substance|Allergies|315,320|false|false|false|C0749139|sulfa|Sulfa
Event|Event|Allergies|315,320|false|false|false|||Sulfa
Drug|Antibiotic|Allergies|322,333|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Organic Chemical|Allergies|322,333|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Pharmacologic Substance|Allergies|322,333|false|false|false|C0038760;C0599503;C3536763|Sulfonamide Anti-Infective Agents;Sulfonamide [EPC];Sulfonamides|Sulfonamide
Drug|Antibiotic|Allergies|334,345|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|Antibiotics
Event|Event|Allergies|334,345|false|false|false|||Antibiotics
Drug|Organic Chemical|Allergies|349,356|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|Allergies|349,356|false|false|false|C0699142|Tylenol|Tylenol
Drug|Organic Chemical|Allergies|359,372|false|false|false|C0012306|hydromorphone|Hydromorphone
Drug|Pharmacologic Substance|Allergies|359,372|false|false|false|C0012306|hydromorphone|Hydromorphone
Event|Event|Allergies|359,372|false|false|false|||Hydromorphone
Drug|Organic Chemical|Allergies|376,383|false|false|false|C0146226|Toradol|Toradol
Drug|Pharmacologic Substance|Allergies|376,383|false|false|false|C0146226|Toradol|Toradol
Event|Event|Allergies|386,395|false|false|false|||Attending
Finding|Functional Concept|Allergies|386,395|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|424,433|false|false|false|||admission
Procedure|Health Care Activity|Chief Complaint|424,433|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Functional Concept|Chief Complaint|435,443|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Finding|Intellectual Product|Chief Complaint|435,443|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|444,463|false|false|false|C0038902|Gynecologic Surgical Procedures|gynecologic surgery
Event|Event|Chief Complaint|456,463|false|false|false|||surgery
Finding|Finding|Chief Complaint|456,463|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Chief Complaint|456,463|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Chief Complaint|456,463|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|456,463|false|false|false|C0543467|Operative Surgical Procedures|surgery
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|468,475|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|Chief Complaint|477,486|false|false|false|C1318143|Retention - dental|retention
Event|Event|Chief Complaint|477,486|false|false|false|||retention
Finding|Cell Function|Chief Complaint|477,486|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|Chief Complaint|477,486|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|Chief Complaint|477,486|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Event|Event|Chief Complaint|496,504|false|false|false|||transfer
Finding|Functional Concept|Chief Complaint|496,504|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|Chief Complaint|496,504|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|Chief Complaint|496,504|false|false|false|C4706767|Transfer (immobility management)|transfer
Disorder|Disease or Syndrome|Chief Complaint|506,517|false|false|false|C0850803|Anaphylaxis;non medication|Anaphylaxis
Event|Event|Chief Complaint|506,517|false|false|false|||Anaphylaxis
Finding|Pathologic Function|Chief Complaint|506,517|false|false|false|C0002792;C4316895|Anaphylactic shock;anaphylaxis|Anaphylaxis
Finding|Classification|Chief Complaint|520,525|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|526,534|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|526,534|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|538,556|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|547,556|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|547,556|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|547,556|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|547,556|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|547,556|false|false|false|C0184661|Interventional procedure|Procedure
Attribute|Clinical Attribute|Chief Complaint|558,563|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Chief Complaint|558,565|false|false|false|C0441767|Stage level 2|Stage 2
Event|Event|Chief Complaint|566,575|false|false|false|||interstim
Disorder|Disease or Syndrome|Chief Complaint|579,588|false|false|false|C0751438|Posterior pituitary disease|posterior
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|579,601|false|false|false|C0195230;C5574717|Posterior repair of vagina;Repair of rectocele|posterior colporrhaphy
Event|Event|Chief Complaint|589,601|false|false|false|||colporrhaphy
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|589,601|false|false|false|C0009416|Suture of vagina|colporrhaphy
Disorder|Acquired Abnormality|Chief Complaint|606,615|false|false|false|C0149771|Rectocele|rectocele
Event|Event|Chief Complaint|606,615|false|false|false|||rectocele
Disorder|Anatomical Abnormality|Chief Complaint|619,629|false|false|false|C0205792|Enterocele|enterocele
Event|Event|Chief Complaint|619,629|false|false|false|||enterocele
Event|Event|History of Present Illness|664,671|false|false|false|||History
Finding|Conceptual Entity|History of Present Illness|664,671|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|History of Present Illness|664,671|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|History of Present Illness|664,671|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|History of Present Illness|664,674|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|History of Present Illness|664,690|false|false|false|C0488508||History of Present Illness
Finding|Finding|History of Present Illness|664,690|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|History of Present Illness|675,682|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|History of Present Illness|675,682|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|History of Present Illness|675,690|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|History of Present Illness|683,690|false|false|false|C0221423|Illness (finding)|Illness
Anatomy|Body Location or Region|History of Present Illness|720,728|false|false|false|C0027530|Neck|cervical
Disorder|Neoplastic Process|History of Present Illness|720,731|false|false|false|C4048328|cervical cancer|cervical CA
Event|Event|History of Present Illness|729,731|false|false|false|||CA
Drug|Chemical Viewed Structurally|History of Present Illness|736,743|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|736,756|false|false|false|C2987682|Radical hysterectomy|radical hysterectomy
Event|Event|History of Present Illness|744,756|false|false|false|||hysterectomy
Finding|Finding|History of Present Illness|744,756|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|744,756|false|false|false|C0020699|Hysterectomy|hysterectomy
Event|Event|History of Present Illness|761,768|false|false|false|||chronic
Finding|Intellectual Product|History of Present Illness|761,768|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|761,768|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|History of Present Illness|774,784|false|false|false|C0024236|Lymphedema|lymphedema
Event|Event|History of Present Illness|774,784|false|false|false|||lymphedema
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|789,796|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|History of Present Illness|789,806|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|History of Present Illness|789,806|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|History of Present Illness|797,806|false|false|false|C1318143|Retention - dental|retention
Event|Event|History of Present Illness|797,806|false|false|false|||retention
Finding|Cell Function|History of Present Illness|797,806|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|History of Present Illness|797,806|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|History of Present Illness|797,806|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Idea or Concept|History of Present Illness|834,838|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|History of Present Illness|834,838|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Disorder|Disease or Syndrome|History of Present Illness|846,852|false|false|false|C0004096|Asthma|Asthma
Event|Event|History of Present Illness|846,852|false|false|false|||Asthma
Disorder|Disease or Syndrome|History of Present Illness|854,858|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|History of Present Illness|854,858|false|false|false|||GERD
Disorder|Congenital Abnormality|History of Present Illness|860,863|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Disorder|Disease or Syndrome|History of Present Illness|860,863|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Event|Event|History of Present Illness|860,863|false|false|false|||IBS
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|865,872|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|865,872|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|865,872|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|873,883|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|History of Present Illness|873,883|false|false|false|||depression
Finding|Functional Concept|History of Present Illness|873,883|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|History of Present Illness|873,883|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|History of Present Illness|885,897|false|false|false|C0016053|Fibromyalgia|fibromyalgia
Event|Event|History of Present Illness|885,897|false|false|false|||fibromyalgia
Event|Event|History of Present Illness|909,915|false|false|false|||issues
Event|Event|History of Present Illness|924,932|false|false|false|||admitted
Finding|Functional Concept|History of Present Illness|940,948|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Finding|Intellectual Product|History of Present Illness|940,948|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Event|Event|History of Present Illness|949,960|false|false|false|||gynecologic
Event|Event|History of Present Illness|962,969|false|false|false|||surgery
Finding|Finding|History of Present Illness|962,969|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|962,969|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|962,969|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|962,969|false|false|false|C0543467|Operative Surgical Procedures|surgery
Attribute|Clinical Attribute|History of Present Illness|971,976|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|History of Present Illness|971,978|false|false|false|C0441767|Stage level 2|stage 2
Disorder|Disease or Syndrome|History of Present Illness|993,1002|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|History of Present Illness|993,1002|false|false|false|||posterior
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|993,1015|false|false|false|C0195230;C5574717|Posterior repair of vagina;Repair of rectocele|posterior colporrhaphy
Event|Event|History of Present Illness|1003,1015|false|false|false|||colporrhaphy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1003,1015|false|false|false|C0009416|Suture of vagina|colporrhaphy
Anatomy|Tissue|History of Present Illness|1019,1024|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|History of Present Illness|1019,1024|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|History of Present Illness|1019,1024|false|false|false|||graft
Finding|Intellectual Product|History of Present Illness|1019,1024|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1019,1024|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1031,1038|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|History of Present Illness|1031,1048|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|History of Present Illness|1031,1048|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|History of Present Illness|1039,1048|false|false|false|C1318143|Retention - dental|retention
Event|Event|History of Present Illness|1039,1048|false|false|false|||retention
Finding|Cell Function|History of Present Illness|1039,1048|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|History of Present Illness|1039,1048|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|History of Present Illness|1039,1048|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Disorder|Acquired Abnormality|History of Present Illness|1053,1062|false|false|false|C0149771|Rectocele|rectocele
Event|Event|History of Present Illness|1053,1062|false|false|false|||rectocele
Disorder|Anatomical Abnormality|History of Present Illness|1065,1075|false|false|false|C0205792|Enterocele|enterocele
Event|Event|History of Present Illness|1065,1075|false|false|false|||enterocele
Anatomy|Body Location or Region|Past Medical History|1103,1111|false|false|false|C0027530|Neck|Cervical
Disorder|Neoplastic Process|Past Medical History|1103,1114|false|true|false|C4048328|cervical cancer|Cervical CA
Event|Event|Past Medical History|1112,1114|false|false|false|||CA
Drug|Chemical Viewed Structurally|Past Medical History|1119,1126|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1119,1139|false|false|false|C2987682|Radical hysterectomy|radical hysterectomy
Event|Event|Past Medical History|1127,1139|false|false|false|||hysterectomy
Finding|Finding|Past Medical History|1127,1139|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1127,1139|false|false|false|C0020699|Hysterectomy|hysterectomy
Event|Event|Past Medical History|1144,1151|false|false|false|||chronic
Finding|Intellectual Product|Past Medical History|1144,1151|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Past Medical History|1144,1151|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Past Medical History|1156,1166|false|false|false|C0024236|Lymphedema|lymphedema
Event|Event|Past Medical History|1156,1166|false|false|false|||lymphedema
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1167,1171|false|false|false|C1263846|Attention deficit hyperactivity disorder|ADHD
Event|Event|Past Medical History|1167,1171|false|false|false|||ADHD
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1172,1179|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Past Medical History|1172,1179|false|false|false|||Anxiety
Finding|Sign or Symptom|Past Medical History|1172,1179|false|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1180,1190|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Event|Event|Past Medical History|1180,1190|false|false|false|||Depression
Finding|Functional Concept|Past Medical History|1180,1190|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|Past Medical History|1180,1190|false|false|false|C0460137;C1579931|Depression - motion|Depression
Disorder|Disease or Syndrome|Past Medical History|1191,1197|false|false|false|C0004096|Asthma|Asthma
Event|Event|Past Medical History|1191,1197|false|false|false|||Asthma
Drug|Pharmacologic Substance|Past Medical History|1198,1206|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Past Medical History|1198,1206|false|false|false|||Insomnia
Finding|Sign or Symptom|Past Medical History|1198,1206|false|false|false|C0917801|Sleeplessness|Insomnia
Disorder|Disease or Syndrome|Past Medical History|1207,1211|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1207,1211|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|1212,1219|false|false|false|C0034734|Raynaud Disease|Raynaud
Disorder|Congenital Abnormality|Past Medical History|1222,1225|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Disorder|Disease or Syndrome|Past Medical History|1222,1225|false|false|false|C0022104;C0432306|Ichthyosis Bullosa of Siemens;Irritable Bowel Syndrome|IBS
Event|Event|Past Medical History|1222,1225|false|false|false|||IBS
Disorder|Disease or Syndrome|Past Medical History|1226,1238|false|false|false|C0016053|Fibromyalgia|Fibromyalgia
Event|Event|Past Medical History|1226,1238|false|false|false|||Fibromyalgia
Event|Event|Family Medical History|1287,1292|false|false|false|||atopy
Finding|Gene or Genome|Family Medical History|1287,1292|false|false|false|C0392707;C3539705|Atopy;MS4A2 wt Allele|atopy
Finding|Pathologic Function|Family Medical History|1287,1292|false|false|false|C0392707;C3539705|Atopy;MS4A2 wt Allele|atopy
Finding|Gene or Genome|Family Medical History|1296,1299|false|false|false|C1420310|SON gene|son
Finding|Finding|Family Medical History|1328,1335|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|Family Medical History|1328,1335|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|Family Medical History|1328,1335|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|Family Medical History|1328,1335|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Event|Event|Family Medical History|1336,1340|false|false|false|||rxns
Event|Event|Family Medical History|1342,1351|false|false|false|||requiring
Disorder|Disease or Syndrome|Family Medical History|1352,1355|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1352,1355|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|Family Medical History|1352,1355|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|Family Medical History|1352,1355|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|Family Medical History|1352,1355|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|Family Medical History|1352,1355|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|Family Medical History|1352,1355|false|false|false|||epi
Finding|Gene or Genome|Family Medical History|1352,1355|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|Family Medical History|1352,1355|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|Family Medical History|1352,1355|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Event|Event|Family Medical History|1356,1360|false|false|false|||pens
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1356,1360|false|false|false|C1527077|Peripheral Electronic Nerve Stimulation|pens
Procedure|Health Care Activity|General Exam|1383,1392|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|1393,1397|false|false|false|||EXAM
Finding|Functional Concept|General Exam|1393,1397|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|1393,1397|false|false|false|C0582103|Medical Examination|EXAM
Finding|Finding|General Exam|1479,1483|true|false|false|C5575035|Well (answer to question)|Well
Finding|Finding|General Exam|1501,1521|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|1507,1512|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|1513,1521|true|false|false|||distress
Finding|Finding|General Exam|1513,1521|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|1513,1521|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Finding|General Exam|1533,1546|true|false|false|C1846018|Muffled voice|muffled voice
Event|Event|General Exam|1541,1546|true|false|false|||voice
Finding|Idea or Concept|General Exam|1541,1546|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|1541,1546|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|1541,1546|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Finding|General Exam|1548,1556|false|false|false|C2984079|Somewhat|somewhat
Finding|Sign or Symptom|General Exam|1557,1564|false|false|false|C0016382|Flushing|flushed
Finding|Sign or Symptom|General Exam|1557,1569|false|false|false|C0016382|Flushing|flushed skin
Anatomy|Body System|General Exam|1565,1569|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|1565,1569|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|1565,1569|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|General Exam|1565,1569|false|false|false|||skin
Finding|Body Substance|General Exam|1565,1569|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|1565,1569|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Location or Region|General Exam|1570,1575|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|1577,1599|true|false|false|C0517391|Moist mucous membranes|Moist mucous membranes
Finding|Body Substance|General Exam|1583,1589|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|General Exam|1583,1599|true|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|General Exam|1583,1599|true|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|General Exam|1590,1599|true|false|false|C0025255|Membrane Tissue|membranes
Finding|Intellectual Product|General Exam|1601,1605|true|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|1606,1609|true|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|General Exam|1606,1609|true|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|General Exam|1606,1609|true|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|General Exam|1606,1609|true|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Finding|Sign or Symptom|General Exam|1606,1618|true|false|false|C0240211|Lip swelling|lip swelling
Event|Event|General Exam|1610,1618|true|false|false|||swelling
Finding|Finding|General Exam|1610,1618|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|1610,1618|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Part, Organ, or Organ Component|General Exam|1620,1626|true|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|1620,1626|true|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|General Exam|1620,1626|true|false|false|C0872394|Procedure on tongue|tongue
Event|Event|General Exam|1640,1649|true|false|false|||edematous
Finding|Pathologic Function|General Exam|1640,1649|true|false|false|C0013604|Edema|edematous
Event|Event|General Exam|1654,1664|true|false|false|||angioedema
Finding|Pathologic Function|General Exam|1654,1664|true|false|false|C0002994|Angioedema|angioedema
Anatomy|Body Location or Region|General Exam|1665,1669|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1665,1669|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1665,1669|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1671,1674|false|false|false|||JVP
Finding|Finding|General Exam|1671,1674|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Activity|General Exam|1700,1704|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|1700,1704|false|false|false|||rate
Finding|Idea or Concept|General Exam|1700,1704|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|1709,1715|true|false|false|||rhythm
Finding|Finding|General Exam|1709,1715|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|1709,1715|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|1734,1741|true|false|false|||murmurs
Finding|Finding|General Exam|1734,1741|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|1742,1747|true|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|1749,1754|true|false|false|||Clear
Finding|Idea or Concept|General Exam|1749,1754|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|1758,1770|true|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|1758,1770|true|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|1788,1795|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|1788,1795|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|1796,1801|true|false|false|||rales
Finding|Finding|General Exam|1796,1801|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|1802,1809|true|false|false|||rhonchi
Finding|Finding|General Exam|1802,1809|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|1810,1817|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|1810,1817|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|1810,1817|false|false|false|||Abdomen
Finding|Finding|General Exam|1810,1817|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|1819,1823|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|1819,1823|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|1837,1842|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|1837,1849|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|1843,1849|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|1843,1849|true|false|false|C0037709||sounds
Event|Event|General Exam|1851,1860|true|false|false|||nontender
Event|Event|General Exam|1863,1875|true|false|false|||nondistended
Event|Event|General Exam|1880,1887|true|false|false|||rebound
Event|Event|General Exam|1891,1899|true|false|false|||guarding
Finding|Finding|General Exam|1891,1899|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Activity|General Exam|1913,1918|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|1913,1918|false|false|false|||place
Finding|Functional Concept|General Exam|1913,1918|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|1913,1918|false|false|false|C1533810||place
Disorder|Congenital Abnormality|General Exam|1919,1922|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|1919,1922|false|false|false|||Ext
Finding|Gene or Genome|General Exam|1919,1922|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|1925,1929|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1925,1929|false|false|false|C0687712|warming process|Warm
Finding|Functional Concept|General Exam|1931,1936|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|General Exam|1941,1946|false|false|false|C1717255||edema
Event|Event|General Exam|1941,1946|false|false|false|||edema
Finding|Pathologic Function|General Exam|1941,1946|false|false|false|C0013604|Edema|edema
Finding|Pathologic Function|General Exam|1941,1958|false|false|false|C0085649|Peripheral edema|edema, peripheral
Finding|Organ or Tissue Function|General Exam|1948,1965|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|General Exam|1959,1965|false|false|false|C5890763||pulses
Event|Event|General Exam|1959,1965|false|false|false|||pulses
Finding|Physiologic Function|General Exam|1959,1965|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|1959,1965|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|1980,1985|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|1980,1985|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|1980,1985|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|1980,1985|false|false|false|||alert
Finding|Finding|General Exam|1980,1985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|1980,1985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|1980,1985|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|1990,1998|false|false|false|||oriented
Finding|Finding|General Exam|1990,1998|false|false|false|C1961028|Oriented to place|oriented
Finding|Finding|General Exam|1990,2008|false|false|false|C1961030|Oriented to person|oriented to person
Attribute|Clinical Attribute|General Exam|2002,2008|false|false|false|C5890614||person
Finding|Intellectual Product|General Exam|2002,2008|false|false|false|C1522390|Person Info|person
Finding|Idea or Concept|General Exam|2010,2018|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|General Exam|2035,2044|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|2035,2044|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2035,2044|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2035,2044|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2035,2044|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|2045,2049|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2045,2049|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2045,2049|false|false|false|C0582103|Medical Examination|EXAM
Finding|Finding|General Exam|2131,2135|true|false|false|C5575035|Well (answer to question)|Well
Finding|Finding|General Exam|2153,2173|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|2159,2164|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|2165,2173|true|false|false|||distress
Finding|Finding|General Exam|2165,2173|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2165,2173|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|General Exam|2175,2181|true|false|false|||normal
Event|Event|General Exam|2183,2188|true|false|false|||voice
Finding|Idea or Concept|General Exam|2183,2188|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|2183,2188|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|2183,2188|true|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Finding|General Exam|2190,2198|false|false|false|C2984079|Somewhat|somewhat
Finding|Sign or Symptom|General Exam|2199,2206|false|false|false|C0016382|Flushing|flushed
Finding|Sign or Symptom|General Exam|2199,2211|false|false|false|C0016382|Flushing|flushed skin
Anatomy|Body System|General Exam|2207,2211|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|2207,2211|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|2207,2211|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|2207,2211|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|2207,2211|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Event|Event|General Exam|2218,2227|false|false|false|||prominent
Anatomy|Body Part, Organ, or Organ Component|General Exam|2231,2236|false|false|false|C0043539|Zygomatic bone|malar
Event|Event|General Exam|2238,2250|false|false|false|||distribution
Finding|Cell Function|General Exam|2238,2250|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|General Exam|2238,2250|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Anatomy|Body Location or Region|General Exam|2254,2258|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|General Exam|2254,2258|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|General Exam|2254,2258|false|false|false|||face
Finding|Gene or Genome|General Exam|2254,2258|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Location or Region|General Exam|2259,2264|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2266,2288|false|false|false|C0517391|Moist mucous membranes|Moist mucous membranes
Finding|Body Substance|General Exam|2272,2278|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|mucous
Anatomy|Tissue|General Exam|2272,2288|false|false|false|C0026724|Mucous Membrane|mucous membranes
Finding|Finding|General Exam|2272,2288|false|false|false|C2230150|moisture of mucous membranes (physical finding)|mucous membranes
Anatomy|Tissue|General Exam|2279,2288|false|false|false|C0025255|Membrane Tissue|membranes
Attribute|Clinical Attribute|General Exam|2290,2300|false|false|false|C0550215||appearance
Event|Event|General Exam|2290,2300|false|false|false|||appearance
Procedure|Health Care Activity|General Exam|2290,2300|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Anatomy|Body Location or Region|General Exam|2304,2308|true|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|General Exam|2304,2308|true|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|General Exam|2304,2308|true|false|false|||face
Finding|Gene or Genome|General Exam|2304,2308|true|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|General Exam|2309,2318|true|false|false|||unchanged
Finding|Finding|General Exam|2309,2318|true|false|false|C0442739||unchanged
Anatomy|Body Part, Organ, or Organ Component|General Exam|2336,2342|true|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|2336,2342|true|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|General Exam|2336,2342|true|false|false|C0872394|Procedure on tongue|tongue
Event|Event|General Exam|2347,2356|true|false|false|||edematous
Finding|Pathologic Function|General Exam|2347,2356|true|false|false|C0013604|Edema|edematous
Event|Event|General Exam|2361,2371|true|false|false|||angioedema
Finding|Pathologic Function|General Exam|2361,2371|true|false|false|C0002994|Angioedema|angioedema
Anatomy|Body Location or Region|General Exam|2372,2376|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|2372,2376|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|2372,2376|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|2378,2381|false|false|false|||JVP
Finding|Finding|General Exam|2378,2381|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Activity|General Exam|2407,2411|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|2407,2411|false|false|false|||rate
Finding|Idea or Concept|General Exam|2407,2411|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|2416,2422|true|false|false|||rhythm
Finding|Finding|General Exam|2416,2422|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2416,2422|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|2441,2448|true|false|false|||murmurs
Finding|Finding|General Exam|2441,2448|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2449,2454|true|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|2456,2461|true|false|false|||Clear
Finding|Idea or Concept|General Exam|2456,2461|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|2465,2477|true|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|2465,2477|true|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|2495,2502|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|2495,2502|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|2503,2508|true|false|false|||rales
Finding|Finding|General Exam|2503,2508|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Event|General Exam|2509,2516|true|false|false|||rhonchi
Finding|Finding|General Exam|2509,2516|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|2517,2524|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2517,2524|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|2517,2524|false|false|false|||Abdomen
Finding|Finding|General Exam|2517,2524|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2526,2530|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|2526,2530|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|2544,2549|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|2544,2556|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|2550,2556|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|2550,2556|true|false|false|C0037709||sounds
Event|Event|General Exam|2558,2567|true|false|false|||nontender
Event|Event|General Exam|2570,2582|true|false|false|||nondistended
Event|Event|General Exam|2587,2594|true|false|false|||rebound
Event|Event|General Exam|2598,2606|true|false|false|||guarding
Finding|Finding|General Exam|2598,2606|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Activity|General Exam|2620,2625|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|2620,2625|false|false|false|||place
Finding|Functional Concept|General Exam|2620,2625|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|2620,2625|false|false|false|C1533810||place
Disorder|Congenital Abnormality|General Exam|2626,2629|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|2626,2629|false|false|false|||Ext
Finding|Gene or Genome|General Exam|2626,2629|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|2632,2636|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2632,2636|false|false|false|C0687712|warming process|Warm
Finding|Functional Concept|General Exam|2638,2643|false|false|false|C1883002|Sequence Chromatogram|trace
Attribute|Clinical Attribute|General Exam|2648,2653|false|false|false|C1717255||edema
Event|Event|General Exam|2648,2653|false|false|false|||edema
Finding|Pathologic Function|General Exam|2648,2653|false|false|false|C0013604|Edema|edema
Finding|Pathologic Function|General Exam|2648,2665|false|false|false|C0085649|Peripheral edema|edema, peripheral
Finding|Organ or Tissue Function|General Exam|2655,2672|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|General Exam|2666,2672|false|false|false|C5890763||pulses
Event|Event|General Exam|2666,2672|false|false|false|||pulses
Finding|Physiologic Function|General Exam|2666,2672|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|2666,2672|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|2687,2692|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|2687,2692|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|2687,2692|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|2687,2692|false|false|false|||alert
Finding|Finding|General Exam|2687,2692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|2687,2692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|2687,2692|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|2697,2705|false|false|false|||oriented
Finding|Finding|General Exam|2697,2705|false|false|false|C1961028|Oriented to place|oriented
Finding|Finding|General Exam|2697,2715|false|false|false|C1961030|Oriented to person|oriented to person
Attribute|Clinical Attribute|General Exam|2709,2715|false|false|false|C5890614||person
Finding|Intellectual Product|General Exam|2709,2715|false|false|false|C1522390|Person Info|person
Finding|Idea or Concept|General Exam|2717,2725|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Anatomical Structure|General Exam|2741,2746|false|false|false|C3714591|Floor (anatomic)|Floor
Event|Event|General Exam|2747,2756|false|false|false|||discharge
Finding|Body Substance|General Exam|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|2747,2756|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|2747,2756|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|General Exam|2757,2761|false|false|false|||exam
Finding|Functional Concept|General Exam|2757,2761|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|2757,2761|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|2763,2766|false|false|false|||VSS
Finding|Classification|General Exam|2771,2774|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|2771,2774|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Disorder|Disease or Syndrome|General Exam|2776,2779|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2776,2779|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2776,2779|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2776,2779|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2776,2779|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|2776,2779|false|false|false|||NAD
Finding|Finding|General Exam|2776,2779|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|2780,2781|false|false|false|||A
Attribute|Clinical Attribute|General Exam|2788,2792|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|2788,2792|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|General Exam|2788,2792|false|false|false|||Resp
Attribute|Clinical Attribute|General Exam|2805,2816|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|General Exam|2805,2816|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|General Exam|2805,2816|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|General Exam|2805,2816|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|General Exam|2805,2825|true|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|General Exam|2817,2825|true|false|false|||distress
Finding|Finding|General Exam|2817,2825|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2817,2825|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|General Exam|2827,2835|true|false|false|||speaking
Event|Event|General Exam|2845,2854|false|false|false|||sentences
Finding|Intellectual Product|General Exam|2845,2854|false|false|false|C0876929|Sentence|sentences
Anatomy|Body Location or Region|General Exam|2855,2858|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|2855,2858|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|General Exam|2860,2864|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|2860,2864|false|false|false|||soft
Disorder|Congenital Abnormality|General Exam|2872,2875|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|2872,2875|false|false|false|||Ext
Finding|Gene or Genome|General Exam|2872,2875|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|2877,2883|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|General Exam|2890,2901|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Health Care Activity|General Exam|2929,2938|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2939,2943|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|2939,2943|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|2958,2963|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2958,2963|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2958,2963|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|2964,2967|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|2974,2977|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|2974,2977|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|2974,2977|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|2983,2986|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|2983,2986|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|2983,2986|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|2983,2986|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|2992,2995|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|2992,2995|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3002,3005|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3002,3005|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3002,3005|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3002,3005|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3002,3005|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3009,3012|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3009,3012|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3009,3012|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3009,3012|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3009,3012|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3009,3012|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3019,3023|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3039,3042|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3059,3064|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3059,3064|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3059,3064|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3077,3083|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3089,3094|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3089,3094|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3089,3094|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3101,3104|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|3101,3104|false|false|false|||Eos
Finding|Gene or Genome|General Exam|3101,3104|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3130,3135|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3130,3135|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3130,3135|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3140,3143|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|3140,3143|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|3140,3143|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3165,3170|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3165,3170|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3165,3170|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3165,3178|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3165,3178|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3165,3178|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3171,3178|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3171,3178|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3171,3178|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3171,3178|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3171,3178|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3171,3178|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3224,3228|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3224,3228|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3224,3228|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3253,3258|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3253,3258|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3253,3258|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3253,3266|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3259,3266|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3259,3266|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3259,3266|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3259,3266|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3259,3266|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3259,3266|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3259,3266|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3259,3266|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3300,3305|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3300,3305|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3300,3305|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3300,3314|false|false|false|C1328414|Blood tryptase|BLOOD TRYPTASE
Drug|Amino Acid, Peptide, or Protein|General Exam|3306,3314|false|false|false|C0147080|TRYPTASE|TRYPTASE
Drug|Enzyme|General Exam|3306,3314|false|false|false|C0147080|TRYPTASE|TRYPTASE
Event|Event|General Exam|3306,3314|false|false|false|||TRYPTASE
Procedure|Laboratory Procedure|General Exam|3306,3314|false|false|false|C1328729|Tryptase measurement|TRYPTASE
Disorder|Disease or Syndrome|General Exam|3315,3318|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|General Exam|3315,3318|false|false|false|||PND
Finding|Gene or Genome|General Exam|3315,3318|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|General Exam|3325,3334|false|false|false|||DISCHARGE
Finding|Body Substance|General Exam|3325,3334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3325,3334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3325,3334|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3325,3334|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3335,3339|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|3335,3339|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3354,3359|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3354,3359|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3354,3359|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3360,3363|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3370,3373|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3370,3373|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3370,3373|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3380,3383|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3380,3383|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3380,3383|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3380,3383|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3389,3392|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3389,3392|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3399,3402|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3399,3402|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3399,3402|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3399,3402|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3399,3402|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3406,3409|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3406,3409|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3406,3409|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3406,3409|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3406,3409|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3406,3409|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|3415,3419|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|3415,3419|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3434,3437|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3454,3459|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3454,3459|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3454,3459|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3460,3463|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3480,3485|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3480,3485|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3480,3485|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3480,3493|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3480,3493|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3480,3493|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3486,3493|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3486,3493|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3486,3493|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3486,3493|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3486,3493|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3486,3493|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3539,3543|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3539,3543|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3539,3543|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3568,3573|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3568,3573|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3568,3573|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3568,3581|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3574,3581|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3574,3581|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3574,3581|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3574,3581|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3574,3581|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3574,3581|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3574,3581|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3574,3581|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Amino Acid, Peptide, or Protein|General Exam|3595,3599|false|false|false|C1431987|MCOLN1 protein, human|Mg-2
Drug|Biologically Active Substance|General Exam|3595,3599|false|false|false|C1431987|MCOLN1 protein, human|Mg-2
Finding|Gene or Genome|General Exam|3595,3599|false|false|false|C5890919|MCOLN1 wt Allele|Mg-2
Event|Event|General Exam|3614,3618|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|3614,3618|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3633,3638|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3633,3638|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3633,3638|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3639,3642|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3649,3652|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3649,3652|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3649,3652|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3658,3661|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3658,3661|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3658,3661|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3658,3661|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3667,3670|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3667,3670|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3677,3680|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3677,3680|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3677,3680|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3677,3680|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3677,3680|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3684,3687|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3684,3687|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3684,3687|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3684,3687|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3684,3687|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3684,3687|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3694,3698|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3714,3717|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3734,3739|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3734,3739|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3734,3739|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3752,3758|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3764,3769|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3764,3769|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3764,3769|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3776,3779|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|3776,3779|false|false|false|||Eos
Finding|Gene or Genome|General Exam|3776,3779|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3805,3810|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3805,3810|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3805,3810|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3815,3818|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|3815,3818|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|3815,3818|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3840,3845|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3840,3845|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3840,3845|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3840,3853|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3840,3853|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3840,3853|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3846,3853|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3846,3853|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3846,3853|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3846,3853|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3846,3853|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3846,3853|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3899,3903|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3899,3903|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3899,3903|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3928,3933|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3928,3933|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3928,3933|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3928,3941|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|3934,3941|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|3934,3941|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|3934,3941|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|3934,3941|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|3934,3941|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|3934,3941|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|3934,3941|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|3934,3941|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|3975,3980|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3975,3980|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3975,3980|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|3975,3989|false|false|false|C1328414|Blood tryptase|BLOOD TRYPTASE
Drug|Amino Acid, Peptide, or Protein|General Exam|3981,3989|false|false|false|C0147080|TRYPTASE|TRYPTASE
Drug|Enzyme|General Exam|3981,3989|false|false|false|C0147080|TRYPTASE|TRYPTASE
Event|Event|General Exam|3981,3989|false|false|false|||TRYPTASE
Procedure|Laboratory Procedure|General Exam|3981,3989|false|false|false|C1328729|Tryptase measurement|TRYPTASE
Disorder|Disease or Syndrome|General Exam|3990,3993|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|General Exam|3990,3993|false|false|false|||PND
Finding|Gene or Genome|General Exam|3990,3993|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Event|Event|General Exam|4005,4012|false|false|false|||IMAGING
Finding|Finding|General Exam|4005,4012|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4005,4012|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|4031,4036|true|false|false|||MICRO
Finding|Conceptual Entity|General Exam|4031,4036|true|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|General Exam|4031,4036|true|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|General Exam|4031,4036|true|false|false|C0085672|Microbiology procedure|MICRO
Anatomy|Body Location or Region|Hospital Course|4101,4109|false|false|false|C0027530|Neck|cervical
Disorder|Neoplastic Process|Hospital Course|4101,4112|false|true|false|C4048328|cervical cancer|cervical CA
Event|Event|Hospital Course|4110,4112|false|false|false|||CA
Drug|Chemical Viewed Structurally|Hospital Course|4117,4124|false|false|false|C0302912|Radicals (chemistry)|radical
Event|Event|Hospital Course|4126,4138|false|false|false|||hysterectomy
Finding|Finding|Hospital Course|4126,4138|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4126,4138|false|false|false|C0020699|Hysterectomy|hysterectomy
Event|Event|Hospital Course|4143,4150|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|4143,4150|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|4143,4150|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|4155,4165|false|false|false|C0024236|Lymphedema|lymphedema
Event|Event|Hospital Course|4155,4165|false|false|false|||lymphedema
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4170,4177|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|Hospital Course|4170,4187|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|Hospital Course|4170,4187|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|Hospital Course|4178,4187|false|false|false|C1318143|Retention - dental|retention
Event|Event|Hospital Course|4178,4187|false|false|false|||retention
Finding|Cell Function|Hospital Course|4178,4187|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|Hospital Course|4178,4187|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|Hospital Course|4178,4187|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Disorder|Disease or Syndrome|Hospital Course|4190,4196|false|false|false|C0004096|Asthma|Asthma
Event|Event|Hospital Course|4190,4196|false|false|false|||Asthma
Disorder|Disease or Syndrome|Hospital Course|4198,4202|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Hospital Course|4198,4202|false|false|false|||GERD
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4204,4211|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|4204,4211|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|4204,4211|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4212,4222|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|4212,4222|false|false|false|||depression
Finding|Functional Concept|Hospital Course|4212,4222|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|4212,4222|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|Hospital Course|4224,4236|false|false|false|C0016053|Fibromyalgia|fibromyalgia
Event|Event|Hospital Course|4224,4236|false|false|false|||fibromyalgia
Finding|Intellectual Product|Hospital Course|4259,4275|false|false|false|C1269801|Operative report|operative report
Attribute|Clinical Attribute|Hospital Course|4269,4275|false|false|false|C4255046||report
Event|Event|Hospital Course|4269,4275|false|false|false|||report
Finding|Intellectual Product|Hospital Course|4269,4275|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Hospital Course|4269,4275|false|false|false|C0700287|Reporting|report
Event|Event|Hospital Course|4285,4292|false|false|false|||details
Event|Event|Hospital Course|4314,4320|false|false|false|||course
Event|Event|Hospital Course|4325,4338|false|false|false|||uncomplicated
Attribute|Clinical Attribute|Hospital Course|4366,4370|false|false|false|C2598155||pain
Event|Event|Hospital Course|4366,4370|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4366,4370|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4366,4370|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|4375,4385|false|false|false|||controlled
Drug|Organic Chemical|Hospital Course|4394,4402|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|Hospital Course|4394,4402|false|false|false|C0728755|Dilaudid|dilaudid
Event|Event|Hospital Course|4394,4402|false|false|false|||dilaudid
Drug|Organic Chemical|Hospital Course|4407,4414|false|false|false|C0146226|Toradol|toradol
Drug|Pharmacologic Substance|Hospital Course|4407,4414|false|false|false|C0146226|Toradol|toradol
Event|Event|Hospital Course|4407,4414|false|false|false|||toradol
Finding|Body Substance|Hospital Course|4443,4450|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4443,4450|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4443,4450|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4451,4458|false|false|false|||started
Event|Event|Hospital Course|4459,4466|false|false|false|||feeling
Event|Event|Hospital Course|4467,4472|false|false|false|||itchy
Finding|Sign or Symptom|Hospital Course|4467,4472|false|false|false|C0033774|Pruritus|itchy
Finding|Intellectual Product|Hospital Course|4475,4479|false|false|false|C1720092|Once - dosing instruction fragment|Once
Event|Event|Hospital Course|4488,4496|false|false|false|||returned
Anatomy|Anatomical Structure|Hospital Course|4504,4509|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|4515,4520|false|false|false|||noted
Event|Event|Hospital Course|4521,4530|false|false|false|||sensation
Finding|Finding|Hospital Course|4521,4530|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Hospital Course|4521,4530|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Hospital Course|4521,4530|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4534,4540|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|Hospital Course|4534,4540|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Event|Event|Hospital Course|4534,4540|false|false|false|||tongue
Procedure|Health Care Activity|Hospital Course|4534,4540|false|false|false|C0872394|Procedure on tongue|tongue
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4544,4547|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|Hospital Course|4544,4547|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|Hospital Course|4544,4547|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|Hospital Course|4544,4547|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Finding|Sign or Symptom|Hospital Course|4544,4556|false|false|false|C0240211|Lip swelling|lip swelling
Event|Event|Hospital Course|4548,4556|false|false|false|||swelling
Finding|Finding|Hospital Course|4548,4556|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|4548,4556|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Hospital Course|4558,4568|false|false|false|||difficulty
Finding|Finding|Hospital Course|4558,4568|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Hospital Course|4580,4590|false|false|false|||secretions
Finding|Body Substance|Hospital Course|4580,4590|false|false|false|C0036537|Bodily secretions|secretions
Event|Event|Hospital Course|4598,4604|false|false|false|||change
Finding|Functional Concept|Hospital Course|4598,4604|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4598,4604|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Hospital Course|4598,4607|false|false|false|C0392747|Changing|change in
Event|Event|Hospital Course|4613,4618|false|false|false|||voice
Finding|Idea or Concept|Hospital Course|4613,4618|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|Hospital Course|4613,4618|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|Hospital Course|4613,4618|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Event|Event|Hospital Course|4624,4627|true|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|4624,4627|true|false|false|C0013404|Dyspnea|SOB
Event|Event|Hospital Course|4632,4640|true|false|false|||flushing
Finding|Sign or Symptom|Hospital Course|4632,4640|true|false|false|C0016382|Flushing|flushing
Event|Event|Hospital Course|4645,4652|true|false|false|||stridor
Finding|Sign or Symptom|Hospital Course|4645,4652|true|false|false|C0038450|Stridor|stridor
Event|Event|Hospital Course|4656,4662|true|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|4656,4662|true|false|false|C0043144|Wheezing|wheeze
Event|Event|Hospital Course|4674,4686|false|false|false|||administered
Disorder|Disease or Syndrome|Hospital Course|4690,4693|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4690,4693|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|Hospital Course|4690,4693|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|Hospital Course|4690,4693|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|Hospital Course|4690,4693|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|Hospital Course|4690,4693|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|Hospital Course|4690,4693|false|false|false|||Epi
Finding|Gene or Genome|Hospital Course|4690,4693|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|Hospital Course|4690,4693|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|Hospital Course|4690,4693|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Drug|Organic Chemical|Hospital Course|4694,4697|false|false|false|C0070220|penclomedine|pen
Drug|Pharmacologic Substance|Hospital Course|4694,4697|false|false|false|C0070220|penclomedine|pen
Event|Event|Hospital Course|4694,4697|false|false|false|||pen
Finding|Gene or Genome|Hospital Course|4694,4697|false|false|false|C1424886;C1428887;C1823520|PCSK1N gene;PUM3 gene;TSPAN33 gene|pen
Drug|Organic Chemical|Hospital Course|4699,4709|false|false|false|C0701466|Solu-Medrol|Solumedrol
Drug|Pharmacologic Substance|Hospital Course|4699,4709|false|false|false|C0701466|Solu-Medrol|Solumedrol
Event|Event|Hospital Course|4699,4709|false|false|false|||Solumedrol
Drug|Organic Chemical|Hospital Course|4721,4731|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|4721,4731|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|Hospital Course|4747,4758|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Drug|Pharmacologic Substance|Hospital Course|4747,4758|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Event|Event|Hospital Course|4747,4758|false|false|false|||Hydroxyzine
Event|Event|Hospital Course|4778,4789|false|false|false|||transferred
Event|Event|Hospital Course|4797,4801|false|false|false|||MICU
Event|Activity|Hospital Course|4814,4824|false|false|false|C1283169||monitoring
Event|Event|Hospital Course|4814,4824|false|false|false|||monitoring
Procedure|Health Care Activity|Hospital Course|4814,4824|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Body Substance|Hospital Course|4832,4839|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4832,4839|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4832,4839|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|4832,4843|false|false|false|C0332310|Has patient|patient has
Drug|Pharmacologic Substance|Hospital Course|4853,4857|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Hospital Course|4853,4857|false|false|false|C0740721|Drug problem|drug
Finding|Pathologic Function|Hospital Course|4853,4867|false|false|false|C0013182|Drug Allergy|drug allergies
Attribute|Clinical Attribute|Hospital Course|4858,4867|false|false|false|C1717415||allergies
Event|Event|Hospital Course|4858,4867|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|4858,4867|false|false|false|C0020517|Hypersensitivity|allergies
Event|Event|Hospital Course|4876,4888|false|false|false|||administered
Attribute|Clinical Attribute|Hospital Course|4904,4915|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4904,4915|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|4904,4915|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|4904,4915|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|4935,4944|false|false|false|C0026056|midazolam|Midazolam
Drug|Pharmacologic Substance|Hospital Course|4935,4944|false|false|false|C0026056|midazolam|Midazolam
Event|Event|Hospital Course|4935,4944|false|false|false|||Midazolam
Drug|Organic Chemical|Hospital Course|4946,4956|false|false|false|C0209337|rocuronium|Rocuronium
Drug|Pharmacologic Substance|Hospital Course|4946,4956|false|false|false|C0209337|rocuronium|Rocuronium
Event|Event|Hospital Course|4946,4956|false|false|false|||Rocuronium
Drug|Organic Chemical|Hospital Course|4959,4967|false|false|false|C0015846|fentanyl|Fentanyl
Drug|Pharmacologic Substance|Hospital Course|4959,4967|false|false|false|C0015846|fentanyl|Fentanyl
Event|Event|Hospital Course|4959,4967|false|false|false|||Fentanyl
Procedure|Laboratory Procedure|Hospital Course|4959,4967|false|false|false|C0524136|Fentanyl measurement|Fentanyl
Drug|Organic Chemical|Hospital Course|4969,4982|false|false|false|C0011777|dexamethasone|Dexamethasone
Drug|Pharmacologic Substance|Hospital Course|4969,4982|false|false|false|C0011777|dexamethasone|Dexamethasone
Event|Event|Hospital Course|4969,4982|false|false|false|||Dexamethasone
Drug|Organic Chemical|Hospital Course|4984,4997|false|false|false|C0012306|hydromorphone|Hydromorphone
Drug|Pharmacologic Substance|Hospital Course|4984,4997|false|false|false|C0012306|hydromorphone|Hydromorphone
Event|Event|Hospital Course|4984,4997|false|false|false|||Hydromorphone
Drug|Organic Chemical|Hospital Course|4999,5010|false|false|false|C0061851|ondansetron|Ondansetron
Drug|Pharmacologic Substance|Hospital Course|4999,5010|false|false|false|C0061851|ondansetron|Ondansetron
Event|Event|Hospital Course|4999,5010|false|false|false|||Ondansetron
Drug|Organic Chemical|Hospital Course|5012,5021|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|5012,5021|false|false|false|C0023660|lidocaine|Lidocaine
Event|Event|Hospital Course|5012,5021|false|false|false|||Lidocaine
Procedure|Laboratory Procedure|Hospital Course|5012,5021|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Organic Chemical|Hospital Course|5024,5032|false|false|false|C0033487|propofol|Propofol
Drug|Pharmacologic Substance|Hospital Course|5024,5032|false|false|false|C0033487|propofol|Propofol
Drug|Antibiotic|Hospital Course|5034,5043|false|false|false|C0007546|cefazolin|Cefazolin
Drug|Organic Chemical|Hospital Course|5034,5043|false|false|false|C0007546|cefazolin|Cefazolin
Event|Event|Hospital Course|5034,5043|false|false|false|||Cefazolin
Drug|Organic Chemical|Hospital Course|5045,5059|false|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Drug|Pharmacologic Substance|Hospital Course|5045,5059|false|false|false|C0017970|glycopyrrolate|Glycopyrrolate
Event|Event|Hospital Course|5045,5059|false|false|false|||Glycopyrrolate
Drug|Organic Chemical|Hospital Course|5061,5074|false|false|false|C0031469|phenylephrine|Phenylephrine
Drug|Pharmacologic Substance|Hospital Course|5061,5074|false|false|false|C0031469|phenylephrine|Phenylephrine
Event|Event|Hospital Course|5061,5074|false|false|false|||Phenylephrine
Drug|Organic Chemical|Hospital Course|5081,5090|false|false|false|C0073631|ketorolac|Ketorolac
Drug|Pharmacologic Substance|Hospital Course|5081,5090|false|false|false|C0073631|ketorolac|Ketorolac
Event|Event|Hospital Course|5081,5090|false|false|false|||Ketorolac
Finding|Idea or Concept|Hospital Course|5106,5113|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|Hospital Course|5114,5116|false|false|false|||VS
Event|Event|Hospital Course|5122,5124|false|false|false|||HR
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5129,5135|false|false|false|C2715713|BP 100|BP 100
Drug|Biologically Active Substance|Hospital Course|5129,5135|false|false|false|C2715713|BP 100|BP 100
Finding|Body Substance|Hospital Course|5165,5172|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5165,5172|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5165,5172|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|5180,5183|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Hospital Course|5180,5183|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Hospital Course|5180,5183|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|5180,5183|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Hospital Course|5180,5183|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Hospital Course|5180,5183|true|false|false|||NAD
Finding|Finding|Hospital Course|5180,5183|true|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|Hospital Course|5193,5199|true|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|5193,5199|true|false|false|C0043144|Wheezing|wheeze
Finding|Intellectual Product|Hospital Course|5203,5207|true|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|Hospital Course|5208,5211|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|5208,5211|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|5208,5211|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Hospital Course|5208,5211|true|false|false|||air
Finding|Finding|Hospital Course|5208,5211|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|5208,5211|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|5208,5211|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Hospital Course|5213,5221|true|false|false|||movement
Finding|Organism Function|Hospital Course|5213,5221|true|false|false|C0026649|Movement|movement
Event|Event|Hospital Course|5225,5229|false|false|false|||exam
Finding|Functional Concept|Hospital Course|5225,5229|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|5225,5229|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|5235,5245|false|false|false|||complained
Finding|Idea or Concept|Hospital Course|5260,5265|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|Hospital Course|5260,5265|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|Hospital Course|5260,5265|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5260,5272|false|false|false|C1527344|Dysphonia|voice change
Finding|Sign or Symptom|Hospital Course|5260,5272|false|false|false|C0518179|Change in voice (finding)|voice change
Event|Event|Hospital Course|5266,5272|false|false|false|||change
Finding|Functional Concept|Hospital Course|5266,5272|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5266,5272|false|false|false|C4319952|Change - procedure|change
Event|Event|Hospital Course|5278,5288|false|false|false|||difficulty
Finding|Finding|Hospital Course|5278,5288|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Hospital Course|5289,5299|false|false|false|||swallowing
Event|Event|Hospital Course|5315,5323|false|false|false|||required
Disorder|Disease or Syndrome|Hospital Course|5331,5334|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5331,5334|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|Hospital Course|5331,5334|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|Hospital Course|5331,5334|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|Hospital Course|5331,5334|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|Hospital Course|5331,5334|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|Hospital Course|5331,5334|false|false|false|||epi
Finding|Gene or Genome|Hospital Course|5331,5334|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|Hospital Course|5331,5334|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|Hospital Course|5331,5334|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Event|Event|Hospital Course|5335,5339|false|false|false|||pens
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5335,5339|false|false|false|C1527077|Peripheral Electronic Nerve Stimulation|pens
Event|Event|Hospital Course|5347,5355|true|false|false|||remained
Finding|Finding|Hospital Course|5356,5378|true|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|Hospital Course|5372,5378|true|false|false|||stable
Finding|Intellectual Product|Hospital Course|5372,5378|true|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|5391,5402|true|false|false|C0231832|Respiratory rate|respiratory
Event|Event|Hospital Course|5391,5402|true|false|false|||respiratory
Finding|Body Substance|Hospital Course|5391,5402|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|5391,5402|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|5391,5402|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|Hospital Course|5404,5414|true|false|false|||compromise
Finding|Social Behavior|Hospital Course|5404,5414|true|false|false|C2945640|compromise|compromise
Event|Event|Hospital Course|5424,5430|false|false|false|||ISSUES
Finding|Gene or Genome|Hospital Course|5436,5440|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|Post
Finding|Finding|Hospital Course|5436,5450|false|false|false|C0241311|post operative (finding)|Post operative
Event|Activity|Hospital Course|5451,5455|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|5451,5455|false|false|false|||care
Finding|Finding|Hospital Course|5451,5455|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|5451,5455|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|Hospital Course|5460,5464|false|false|false|C2598155||pain
Event|Event|Hospital Course|5460,5464|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5460,5464|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5460,5464|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|5469,5479|false|false|false|||controlled
Event|Event|Hospital Course|5492,5499|false|false|false|||post-op
Drug|Organic Chemical|Hospital Course|5508,5516|false|false|false|C0728755|Dilaudid|dilaudid
Drug|Pharmacologic Substance|Hospital Course|5508,5516|false|false|false|C0728755|Dilaudid|dilaudid
Event|Event|Hospital Course|5508,5516|false|false|false|||dilaudid
Drug|Organic Chemical|Hospital Course|5522,5529|false|false|false|C0146226|Toradol|toradol
Drug|Pharmacologic Substance|Hospital Course|5522,5529|false|false|false|C0146226|Toradol|toradol
Event|Event|Hospital Course|5522,5529|false|false|false|||toradol
Event|Event|Hospital Course|5540,5552|false|false|false|||transitioned
Drug|Organic Chemical|Hospital Course|5559,5568|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|5559,5568|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|5559,5568|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|5559,5568|false|false|false|C0524222|Oxycodone measurement|oxycodone
Event|Event|Hospital Course|5580,5589|false|false|false|||difficult
Finding|Finding|Hospital Course|5580,5589|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|Hospital Course|5593,5602|false|false|false|||determine
Event|Event|Hospital Course|5612,5619|false|false|false|||causing
Finding|Functional Concept|Hospital Course|5623,5631|false|false|false|C0700624|Allergic|allergic
Finding|Pathologic Function|Hospital Course|5623,5640|false|false|false|C0020517;C1527304|Allergic Reaction;Hypersensitivity|allergic reaction
Event|Event|Hospital Course|5632,5640|false|false|false|||reaction
Finding|Functional Concept|Hospital Course|5632,5640|false|false|false|C0443286|Reaction|reaction
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5659,5666|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Hospital Course|5659,5666|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Hospital Course|5659,5666|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Hospital Course|5659,5666|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5659,5674|false|false|false|C1270937|Insertion of pack into vagina|vaginal packing
Drug|Biomedical or Dental Material|Hospital Course|5667,5674|false|false|false|C1706363|Packing Dosage Form|packing
Event|Activity|Hospital Course|5667,5674|false|false|false|C2828395|Packing (action)|packing
Event|Event|Hospital Course|5667,5674|false|false|false|||packing
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5667,5674|false|false|false|C0184967|Insertion of pack (procedure)|packing
Event|Event|Hospital Course|5679,5686|false|false|false|||removed
Event|Event|Hospital Course|5715,5718|false|false|false|||day
Finding|Idea or Concept|Hospital Course|5715,5718|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5715,5718|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|Hospital Course|5727,5732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|5727,5732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|5727,5732|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|Hospital Course|5727,5739|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5727,5739|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|Hospital Course|5733,5739|false|false|false|||output
Finding|Conceptual Entity|Hospital Course|5733,5739|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|5733,5739|false|false|false|C3251815|Measurement of fluid output|output
Event|Event|Hospital Course|5744,5752|false|false|false|||adequate
Event|Event|Hospital Course|5771,5778|false|false|false|||removed
Finding|Body Substance|Hospital Course|5785,5792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5785,5792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5785,5792|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5797,5801|false|false|false|||able
Finding|Finding|Hospital Course|5797,5801|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|5833,5840|false|false|false|||require
Finding|Idea or Concept|Hospital Course|5842,5846|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Finding|Intellectual Product|Hospital Course|5842,5846|false|false|false|C0036588;C1551994|Self;subscriber - self|self
Event|Event|Hospital Course|5847,5862|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5847,5862|false|false|false|C0007430|Catheterization|catheterization
Disorder|Disease or Syndrome|Hospital Course|5867,5872|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5875,5878|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5875,5878|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5890,5899|false|false|false|||sensation
Finding|Finding|Hospital Course|5890,5899|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Hospital Course|5890,5899|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Hospital Course|5890,5899|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5904,5911|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|5904,5911|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|Hospital Course|5904,5911|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5904,5911|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Disease or Syndrome|Hospital Course|5927,5938|false|false|false|C0850803|Anaphylaxis;non medication|Anaphylaxis
Event|Event|Hospital Course|5927,5938|false|false|false|||Anaphylaxis
Finding|Pathologic Function|Hospital Course|5927,5938|false|false|false|C0002792;C4316895|Anaphylactic shock;anaphylaxis|Anaphylaxis
Finding|Body Substance|Hospital Course|5957,5964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5957,5964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5957,5964|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|5965,5970|false|false|false|||awoke
Event|Event|Hospital Course|5975,5982|false|false|false|||started
Event|Event|Hospital Course|5991,5999|false|false|false|||pruritis
Finding|Sign or Symptom|Hospital Course|5991,5999|false|false|false|C0033774|Pruritus|pruritis
Finding|Intellectual Product|Hospital Course|6001,6005|false|false|false|C1720092|Once - dosing instruction fragment|Once
Event|Event|Hospital Course|6011,6018|false|false|false|||arrived
Anatomy|Anatomical Structure|Hospital Course|6026,6031|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|Hospital Course|6037,6044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6037,6044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6037,6044|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6045,6050|false|false|false|||noted
Event|Event|Hospital Course|6051,6061|false|false|false|||difficulty
Finding|Finding|Hospital Course|6051,6061|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Hospital Course|6062,6069|false|false|false|||talking
Finding|Finding|Hospital Course|6085,6092|false|false|false|C0038999|Swelling|swollen
Finding|Sign or Symptom|Hospital Course|6085,6097|false|false|false|C0240211|Lip swelling|swollen lips
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6093,6097|false|false|false|C0023759|Lip structure|lips
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6098,6104|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|Hospital Course|6098,6104|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|Hospital Course|6098,6104|false|false|false|C0872394|Procedure on tongue|tongue
Finding|Functional Concept|Hospital Course|6110,6115|false|false|false|C0205382|vocal|vocal
Event|Event|Hospital Course|6116,6123|false|false|false|||changes
Finding|Functional Concept|Hospital Course|6116,6123|false|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|6128,6131|true|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|6128,6131|true|false|false|C0013404|Dyspnea|SOB
Event|Event|Hospital Course|6137,6145|true|false|false|||flushing
Finding|Sign or Symptom|Hospital Course|6137,6145|true|false|false|C0016382|Flushing|flushing
Event|Event|Hospital Course|6150,6157|true|false|false|||stridor
Finding|Sign or Symptom|Hospital Course|6150,6157|true|false|false|C0038450|Stridor|stridor
Event|Event|Hospital Course|6161,6167|true|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|6161,6167|true|false|false|C0043144|Wheezing|wheeze
Attribute|Clinical Attribute|Hospital Course|6171,6178|false|false|false|C0032930|Precipitating Factors|trigger
Event|Event|Hospital Course|6183,6189|false|false|false|||called
Event|Event|Hospital Course|6195,6207|false|false|false|||anaphyllaxis
Event|Event|Hospital Course|6216,6224|false|false|false|||recieved
Disorder|Disease or Syndrome|Hospital Course|6228,6231|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6228,6231|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|Hospital Course|6228,6231|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|Hospital Course|6228,6231|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|Hospital Course|6228,6231|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|Hospital Course|6228,6231|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|Hospital Course|6228,6231|false|false|false|||Epi
Finding|Gene or Genome|Hospital Course|6228,6231|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|Hospital Course|6228,6231|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|Hospital Course|6228,6231|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Drug|Organic Chemical|Hospital Course|6232,6235|false|false|false|C0070220|penclomedine|pen
Drug|Pharmacologic Substance|Hospital Course|6232,6235|false|false|false|C0070220|penclomedine|pen
Event|Event|Hospital Course|6232,6235|false|false|false|||pen
Finding|Gene or Genome|Hospital Course|6232,6235|false|false|false|C1424886;C1428887;C1823520|PCSK1N gene;PUM3 gene;TSPAN33 gene|pen
Drug|Organic Chemical|Hospital Course|6237,6247|false|false|false|C0701466|Solu-Medrol|Solumedrol
Drug|Pharmacologic Substance|Hospital Course|6237,6247|false|false|false|C0701466|Solu-Medrol|Solumedrol
Event|Event|Hospital Course|6237,6247|false|false|false|||Solumedrol
Drug|Organic Chemical|Hospital Course|6260,6270|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|Hospital Course|6260,6270|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|Hospital Course|6285,6296|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Drug|Pharmacologic Substance|Hospital Course|6285,6296|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Event|Event|Hospital Course|6285,6296|false|false|false|||Hydroxyzine
Event|Event|Hospital Course|6317,6328|false|false|false|||transferred
Event|Event|Hospital Course|6336,6340|false|false|false|||MICU
Event|Activity|Hospital Course|6352,6362|false|false|false|C1283169||monitoring
Event|Event|Hospital Course|6352,6362|false|false|false|||monitoring
Procedure|Health Care Activity|Hospital Course|6352,6362|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Idea or Concept|Hospital Course|6379,6386|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|Hospital Course|6387,6389|false|false|false|||VS
Event|Event|Hospital Course|6395,6397|false|false|false|||HR
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6402,6408|false|false|false|C2715713|BP 100|BP 100
Drug|Biologically Active Substance|Hospital Course|6402,6408|false|false|false|C2715713|BP 100|BP 100
Finding|Body Substance|Hospital Course|6438,6445|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6438,6445|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6438,6445|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|6453,6456|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Hospital Course|6453,6456|true|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Hospital Course|6453,6456|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|6453,6456|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Hospital Course|6453,6456|true|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Hospital Course|6453,6456|true|false|false|||NAD
Finding|Finding|Hospital Course|6453,6456|true|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|Hospital Course|6466,6472|true|false|false|||wheeze
Finding|Sign or Symptom|Hospital Course|6466,6472|true|false|false|C0043144|Wheezing|wheeze
Finding|Intellectual Product|Hospital Course|6476,6480|true|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|Hospital Course|6481,6484|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|6481,6484|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|6481,6484|true|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Hospital Course|6481,6484|true|false|false|||air
Finding|Finding|Hospital Course|6481,6484|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|6481,6484|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|6481,6484|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Hospital Course|6486,6494|true|false|false|||movement
Finding|Organism Function|Hospital Course|6486,6494|true|false|false|C0026649|Movement|movement
Event|Event|Hospital Course|6498,6502|false|false|false|||exam
Finding|Functional Concept|Hospital Course|6498,6502|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|6498,6502|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|6508,6518|false|false|false|||complained
Finding|Idea or Concept|Hospital Course|6533,6538|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|Hospital Course|6533,6538|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|Hospital Course|6533,6538|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6533,6545|false|false|false|C1527344|Dysphonia|voice change
Finding|Sign or Symptom|Hospital Course|6533,6545|false|false|false|C0518179|Change in voice (finding)|voice change
Event|Event|Hospital Course|6539,6545|false|false|false|||change
Finding|Functional Concept|Hospital Course|6539,6545|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6539,6545|false|false|false|C4319952|Change - procedure|change
Event|Event|Hospital Course|6551,6561|false|false|false|||difficulty
Finding|Finding|Hospital Course|6551,6561|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Hospital Course|6562,6572|false|false|false|||swallowing
Event|Event|Hospital Course|6588,6596|false|false|false|||required
Disorder|Disease or Syndrome|Hospital Course|6604,6607|false|false|false|C0267963|Exocrine pancreatic insufficiency|epi
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6604,6607|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Biologically Active Substance|Hospital Course|6604,6607|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Hormone|Hospital Course|6604,6607|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Organic Chemical|Hospital Course|6604,6607|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Drug|Pharmacologic Substance|Hospital Course|6604,6607|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|epi
Event|Event|Hospital Course|6604,6607|false|false|false|||epi
Finding|Gene or Genome|Hospital Course|6604,6607|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Finding|Intellectual Product|Hospital Course|6604,6607|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|epi
Procedure|Diagnostic Procedure|Hospital Course|6604,6607|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|epi
Event|Event|Hospital Course|6608,6612|false|false|false|||pens
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6608,6612|false|false|false|C1527077|Peripheral Electronic Nerve Stimulation|pens
Event|Event|Hospital Course|6620,6628|true|false|false|||remained
Finding|Finding|Hospital Course|6629,6651|true|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Event|Event|Hospital Course|6645,6651|true|false|false|||stable
Finding|Intellectual Product|Hospital Course|6645,6651|true|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|6664,6675|true|false|false|C0231832|Respiratory rate|respiratory
Event|Event|Hospital Course|6664,6675|true|false|false|||respiratory
Finding|Body Substance|Hospital Course|6664,6675|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|6664,6675|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|6664,6675|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Event|Event|Hospital Course|6677,6687|true|false|false|||compromise
Finding|Social Behavior|Hospital Course|6677,6687|true|false|false|C2945640|compromise|compromise
Finding|Body Substance|Hospital Course|6700,6707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6700,6707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6700,6707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|6712,6717|false|false|false|||lying
Event|Event|Hospital Course|6718,6729|false|false|false|||comfortable
Finding|Finding|Hospital Course|6718,6729|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|Hospital Course|6733,6736|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|Hospital Course|6733,6736|false|false|false|||bed
Finding|Intellectual Product|Hospital Course|6733,6736|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|Hospital Course|6754,6764|false|false|false|||continuing
Event|Event|Hospital Course|6768,6775|false|false|false|||inquire
Disorder|Disease or Syndrome|Hospital Course|6787,6790|false|false|false|C0267963|Exocrine pancreatic insufficiency|Epi
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6787,6790|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Biologically Active Substance|Hospital Course|6787,6790|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Hormone|Hospital Course|6787,6790|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Organic Chemical|Hospital Course|6787,6790|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Drug|Pharmacologic Substance|Hospital Course|6787,6790|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|Epi
Event|Event|Hospital Course|6787,6790|false|false|false|||Epi
Finding|Gene or Genome|Hospital Course|6787,6790|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Finding|Intellectual Product|Hospital Course|6787,6790|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|Epi
Procedure|Diagnostic Procedure|Hospital Course|6787,6790|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|Epi
Event|Event|Hospital Course|6791,6795|false|false|false|||pens
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6791,6795|false|false|false|C1527077|Peripheral Electronic Nerve Stimulation|pens
Drug|Hormone|Hospital Course|6799,6810|false|false|false|C0014563|epinephrine|epinephrine
Drug|Organic Chemical|Hospital Course|6799,6810|false|false|false|C0014563|epinephrine|epinephrine
Drug|Pharmacologic Substance|Hospital Course|6799,6810|false|false|false|C0014563|epinephrine|epinephrine
Event|Event|Hospital Course|6799,6810|false|false|false|||epinephrine
Procedure|Laboratory Procedure|Hospital Course|6799,6810|false|false|false|C0201998|Epinephrine measurement|epinephrine
Disorder|Neoplastic Process|Hospital Course|6811,6814|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|6811,6814|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|Hospital Course|6811,6814|false|false|false|||gtt
Procedure|Laboratory Procedure|Hospital Course|6811,6814|false|false|false|C0017741|Glucose tolerance test|gtt
Finding|Finding|Hospital Course|6824,6835|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|Hospital Course|6836,6847|false|false|false|||respiration
Finding|Cell Function|Hospital Course|6836,6847|false|false|false|C0035203;C0282636|Cell Respiration;Respiration|respiration
Finding|Physiologic Function|Hospital Course|6836,6847|false|false|false|C0035203;C0282636|Cell Respiration;Respiration|respiration
Phenomenon|Biologic Function|Hospital Course|6836,6847|false|false|false|C1160636|respiratory system process|respiration
Event|Event|Hospital Course|6849,6861|false|false|false|||vocalization
Finding|Finding|Hospital Course|6849,6861|false|false|false|C0564182|Vocalization (finding)|vocalization
Anatomy|Body Space or Junction|Hospital Course|6878,6882|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|6878,6882|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|6878,6882|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|6878,6882|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|6883,6893|false|false|false|||structures
Event|Event|Hospital Course|6904,6916|false|false|false|||perseverated
Drug|Organic Chemical|Hospital Course|6927,6933|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|Hospital Course|6927,6933|false|false|false|C0699194|Ativan|Ativan
Drug|Organic Chemical|Hospital Course|6939,6945|false|false|false|C0487782|Ambien|Ambien
Drug|Pharmacologic Substance|Hospital Course|6939,6945|false|false|false|C0487782|Ambien|Ambien
Event|Event|Hospital Course|6939,6945|false|false|false|||Ambien
Finding|Finding|Hospital Course|6950,6954|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|Hospital Course|6962,6973|false|false|false|C0033497|propranolol|propranolol
Drug|Pharmacologic Substance|Hospital Course|6962,6973|false|false|false|C0033497|propranolol|propranolol
Event|Event|Hospital Course|6962,6973|false|false|false|||propranolol
Disorder|Disease or Syndrome|Hospital Course|6978,6994|false|true|false|C0270736|Essential Tremor|essential tremor
Finding|Sign or Symptom|Hospital Course|6988,6994|false|true|false|C0040822|Tremor|tremor
Event|Event|Hospital Course|6995,7002|false|false|false|||despite
Event|Event|Hospital Course|7004,7015|false|false|false|||explanation
Finding|Intellectual Product|Hospital Course|7004,7015|false|false|false|C0681841|Explanation|explanation
Finding|Intellectual Product|Hospital Course|7021,7025|false|false|false|C0439096|Greek letter beta|beta
Drug|Pharmacologic Substance|Hospital Course|7021,7034|false|false|false|C0001645|Adrenergic beta-Antagonists|beta blockers
Event|Event|Hospital Course|7026,7034|false|false|false|||blockers
Event|Event|Hospital Course|7046,7065|false|false|false|||bronchoconstriction
Finding|Organ or Tissue Function|Hospital Course|7046,7065|false|false|false|C0079043;C3536811|Bronchoconstriction;Bronchoconstriction [PE]|bronchoconstriction
Attribute|Clinical Attribute|Hospital Course|7071,7082|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|7071,7082|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|7071,7082|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|7071,7082|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Finding|Hospital Course|7071,7093|false|false|false|C5208132|Respiratory compromise|respiratory compromise
Event|Event|Hospital Course|7083,7093|false|false|false|||compromise
Finding|Social Behavior|Hospital Course|7083,7093|false|false|false|C2945640|compromise|compromise
Disorder|Disease or Syndrome|Hospital Course|7097,7108|false|false|false|C0850803|Anaphylaxis;non medication|anaphylaxis
Event|Event|Hospital Course|7097,7108|false|false|false|||anaphylaxis
Finding|Pathologic Function|Hospital Course|7097,7108|false|false|false|C0002792;C4316895|Anaphylactic shock;anaphylaxis|anaphylaxis
Finding|Idea or Concept|Hospital Course|7118,7121|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7118,7121|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|7130,7136|false|false|false|||called
Anatomy|Anatomical Structure|Hospital Course|7148,7153|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|7162,7172|false|false|false|||complained
Anatomy|Body Location or Region|Hospital Course|7188,7194|false|false|false|C0015450|Face|facial
Finding|Sign or Symptom|Hospital Course|7188,7203|false|false|false|C0016382;C5848177|Face goes red;Flushing|facial flushing
Event|Event|Hospital Course|7195,7203|false|false|false|||flushing
Finding|Sign or Symptom|Hospital Course|7195,7203|false|false|false|C0016382|Flushing|flushing
Event|Event|Hospital Course|7214,7222|true|false|false|||afebrile
Finding|Finding|Hospital Course|7214,7222|true|false|false|C0277797|Apyrexial|afebrile
Event|Event|Hospital Course|7241,7247|true|false|false|||stable
Finding|Intellectual Product|Hospital Course|7241,7247|true|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|7261,7272|true|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Hospital Course|7261,7272|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Hospital Course|7261,7272|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Hospital Course|7261,7272|true|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Finding|Hospital Course|7261,7283|true|false|false|C5208132|Respiratory compromise|respiratory compromise
Event|Event|Hospital Course|7273,7283|true|false|false|||compromise
Finding|Social Behavior|Hospital Course|7273,7283|true|false|false|C2945640|compromise|compromise
Finding|Functional Concept|Hospital Course|7287,7295|true|false|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Finding|Sign or Symptom|Hospital Course|7287,7304|true|false|false|C2039684|systemic symptoms|systemic symptoms
Event|Event|Hospital Course|7296,7304|true|false|false|||symptoms
Finding|Functional Concept|Hospital Course|7296,7304|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|7296,7304|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|Hospital Course|7308,7319|false|false|false|C0231220|Symptomatic|Symptomatic
Event|Activity|Hospital Course|7320,7324|false|false|false|C1947933|care activity|care
Event|Event|Hospital Course|7320,7324|false|false|false|||care
Finding|Finding|Hospital Course|7320,7324|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Hospital Course|7320,7324|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Drug|Organic Chemical|Hospital Course|7330,7341|false|false|false|C0020404|hydroxyzine|hydroxyzine
Drug|Pharmacologic Substance|Hospital Course|7330,7341|false|false|false|C0020404|hydroxyzine|hydroxyzine
Event|Event|Hospital Course|7330,7341|false|false|false|||hydroxyzine
Drug|Organic Chemical|Hospital Course|7346,7353|false|false|false|C0164056|eucerin|eucerin
Drug|Pharmacologic Substance|Hospital Course|7346,7353|false|false|false|C0164056|eucerin|eucerin
Drug|Biomedical or Dental Material|Hospital Course|7354,7360|false|false|false|C0544341|Lotion|lotion
Event|Event|Hospital Course|7354,7360|false|false|false|||lotion
Event|Event|Hospital Course|7366,7374|false|false|false|||provided
Event|Event|Hospital Course|7382,7386|false|false|false|||step
Finding|Conceptual Entity|Hospital Course|7382,7386|false|false|false|C1261552;C1419107;C1704379|PTPN5 gene;Step (specific stage);Treatment Step|step
Finding|Functional Concept|Hospital Course|7382,7386|false|false|false|C1261552;C1419107;C1704379|PTPN5 gene;Step (specific stage);Treatment Step|step
Finding|Gene or Genome|Hospital Course|7382,7386|false|false|false|C1261552;C1419107;C1704379|PTPN5 gene;Step (specific stage);Treatment Step|step
Anatomy|Anatomical Structure|Hospital Course|7399,7404|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|Hospital Course|7410,7417|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7410,7417|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7410,7417|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7424,7432|false|false|false|||reported
Event|Event|Hospital Course|7437,7444|false|false|false|||nursing
Finding|Organism Function|Hospital Course|7437,7444|false|false|false|C0006147|Breast Feeding|nursing
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7437,7444|false|false|false|C0028678|RNAx nursing therapy actions|nursing
Event|Event|Hospital Course|7454,7458|false|false|false|||felt
Anatomy|Body Location or Region|Hospital Course|7459,7465|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7459,7465|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Hospital Course|7459,7465|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|Hospital Course|7459,7465|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Hospital Course|7459,7465|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Finding|Hospital Course|7459,7478|false|false|false|C0236071|Constriction in throat|throat constriction
Anatomy|Cell Component|Hospital Course|7466,7478|false|false|false|C1760025|constriction location|constriction
Event|Event|Hospital Course|7466,7478|false|false|false|||constriction
Finding|Pathologic Function|Hospital Course|7466,7478|false|false|false|C1261287|Stenosis|constriction
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7466,7478|false|false|false|C0009813|Constriction procedure|constriction
Drug|Hormone|Hospital Course|7480,7491|false|false|false|C0014563|epinephrine|Epinephrine
Drug|Organic Chemical|Hospital Course|7480,7491|false|false|false|C0014563|epinephrine|Epinephrine
Drug|Pharmacologic Substance|Hospital Course|7480,7491|false|false|false|C0014563|epinephrine|Epinephrine
Event|Event|Hospital Course|7480,7491|false|false|false|||Epinephrine
Procedure|Laboratory Procedure|Hospital Course|7480,7491|false|false|false|C0201998|Epinephrine measurement|Epinephrine
Drug|Organic Chemical|Hospital Course|7497,7507|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Pharmacologic Substance|Hospital Course|7497,7507|false|false|false|C0701466|Solu-Medrol|solumedrol
Event|Event|Hospital Course|7497,7507|false|false|false|||solumedrol
Event|Event|Hospital Course|7513,7518|false|false|false|||given
Finding|Body Substance|Hospital Course|7527,7534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7527,7534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7527,7534|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|7540,7546|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|Hospital Course|7540,7546|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|Hospital Course|7540,7546|false|false|false|||relief
Finding|Finding|Hospital Course|7540,7546|false|false|false|C0564405|Feeling relief|relief
Finding|Finding|Hospital Course|7548,7555|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Idea or Concept|Hospital Course|7548,7555|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Pathologic Function|Hospital Course|7548,7555|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Physiologic Function|Hospital Course|7548,7555|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Event|Event|Hospital Course|7561,7570|false|false|false|||consulted
Event|Event|Hospital Course|7581,7586|false|false|false|||asked
Event|Event|Hospital Course|7593,7597|false|false|false|||stop
Finding|Finding|Hospital Course|7602,7605|false|false|true|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|7602,7605|false|false|true|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Hospital Course|7602,7617|false|false|true|C1718097|New medications|new medications
Attribute|Clinical Attribute|Hospital Course|7606,7617|false|false|true|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|7606,7617|false|false|true|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|7606,7617|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|7606,7617|false|false|true|C4284232|Medications|medications
Finding|Idea or Concept|Hospital Course|7645,7653|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|7662,7668|false|false|false|||report
Attribute|Clinical Attribute|Hospital Course|7685,7694|false|false|false|C1717415||allergies
Event|Event|Hospital Course|7685,7694|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|7685,7694|false|false|false|C0020517|Hypersensitivity|allergies
Finding|Functional Concept|Hospital Course|7699,7707|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Event|Event|Hospital Course|7712,7716|false|false|false|||sent
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7723,7731|false|false|false|C0147080|TRYPTASE|tryptase
Drug|Enzyme|Hospital Course|7723,7731|false|false|false|C0147080|TRYPTASE|tryptase
Procedure|Laboratory Procedure|Hospital Course|7723,7731|false|false|false|C1328729|Tryptase measurement|tryptase
Event|Event|Hospital Course|7732,7737|false|false|false|||level
Finding|Finding|Hospital Course|7742,7746|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|7751,7762|false|false|false|||coordinated
Event|Event|Hospital Course|7763,7773|false|false|false|||outpatient
Finding|Classification|Hospital Course|7763,7773|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7763,7773|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|7774,7780|false|false|false|||follow
Finding|Functional Concept|Hospital Course|7774,7780|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|7774,7780|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|7774,7783|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|7774,7783|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|7798,7805|false|false|false|||Chronic
Finding|Intellectual Product|Hospital Course|7798,7805|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|7798,7805|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Attribute|Clinical Attribute|Hospital Course|7810,7815|false|false|false|C1717255||edema
Event|Event|Hospital Course|7810,7815|false|false|false|||edema
Finding|Pathologic Function|Hospital Course|7810,7815|false|false|false|C0013604|Edema|edema
Event|Event|Hospital Course|7817,7825|false|false|false|||Continue
Finding|Idea or Concept|Hospital Course|7826,7830|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7826,7830|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7826,7830|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7831,7841|false|false|false|C0025854|metolazone|Metolazone
Drug|Pharmacologic Substance|Hospital Course|7831,7841|false|false|false|C0025854|metolazone|Metolazone
Event|Event|Hospital Course|7831,7841|false|false|false|||Metolazone
Drug|Organic Chemical|Hospital Course|7843,7857|true|false|false|C0037982|spironolactone|spironolactone
Drug|Pharmacologic Substance|Hospital Course|7843,7857|true|false|false|C0037982|spironolactone|spironolactone
Event|Event|Hospital Course|7843,7857|true|false|false|||spironolactone
Drug|Biologically Active Substance|Hospital Course|7860,7869|true|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Hospital Course|7860,7869|true|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Hospital Course|7860,7869|true|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Hospital Course|7860,7869|true|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Hospital Course|7860,7869|true|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Hospital Course|7860,7869|true|false|false|||potassium
Finding|Physiologic Function|Hospital Course|7860,7869|true|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Hospital Course|7860,7869|true|false|false|C0202194|Potassium measurement|potassium
Event|Event|Hospital Course|7870,7879|true|false|false|||repletion
Event|Event|Hospital Course|7887,7898|true|false|false|||hypotensive
Finding|Pathologic Function|Hospital Course|7887,7898|true|false|false|C0857353|Hypotensive|hypotensive
Event|Event|Hospital Course|7904,7913|false|false|false|||monitored
Event|Event|Hospital Course|7932,7936|false|false|false|||stay
Event|Event|Hospital Course|7948,7951|false|false|false|||WNL
Disorder|Disease or Syndrome|Hospital Course|7955,7961|false|false|false|C0004096|Asthma|Asthma
Event|Event|Hospital Course|7955,7961|false|false|false|||Asthma
Event|Event|Hospital Course|7963,7967|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|7963,7967|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|7963,7967|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|7963,7967|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|7968,7977|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|7968,7977|false|false|false|C0001927|albuterol|Albuterol
Event|Event|Hospital Course|7978,7981|false|false|false|||use
Finding|Functional Concept|Hospital Course|7978,7981|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|7978,7981|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Hospital Course|7990,7994|true|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|8004,8011|true|false|false|||require
Event|Event|Hospital Course|8020,8024|true|false|false|||MICU
Disorder|Disease or Syndrome|Hospital Course|8029,8033|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Hospital Course|8029,8033|false|false|false|||GERD
Drug|Organic Chemical|Hospital Course|8035,8041|false|false|false|C0939400|Nexium|Nexium
Drug|Pharmacologic Substance|Hospital Course|8035,8041|false|false|false|C0939400|Nexium|Nexium
Event|Event|Hospital Course|8035,8041|false|false|false|||Nexium
Event|Event|Hospital Course|8057,8061|false|false|false|||held
Event|Event|Hospital Course|8065,8074|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8065,8074|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Activity|Hospital Course|8088,8095|false|false|false|C1272683||request
Event|Event|Hospital Course|8088,8095|false|false|false|||request
Finding|Idea or Concept|Hospital Course|8088,8095|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Finding|Intellectual Product|Hospital Course|8088,8095|false|false|false|C1522634;C1553397;C1553888|Question (inquiry);Request - ActReason;request - ActMood|request
Event|Event|Hospital Course|8100,8105|false|false|false|||given
Drug|Food|Hospital Course|8132,8136|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|8132,8136|false|false|false|||diet
Finding|Functional Concept|Hospital Course|8132,8136|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|8132,8136|false|false|false|C0012159|Diet therapy|diet
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8140,8144|false|false|false|C1263846|Attention deficit hyperactivity disorder|ADHD
Event|Event|Hospital Course|8140,8144|false|false|false|||ADHD
Drug|Organic Chemical|Hospital Course|8149,8157|false|false|false|C0290795|Adderall|Adderall
Drug|Pharmacologic Substance|Hospital Course|8149,8157|false|false|false|C0290795|Adderall|Adderall
Event|Event|Hospital Course|8159,8163|false|false|false|||held
Event|Event|Hospital Course|8167,8176|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|8167,8176|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8180,8187|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|8180,8187|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|8180,8187|false|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8188,8198|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Hospital Course|8188,8198|false|false|false|||depression
Finding|Functional Concept|Hospital Course|8188,8198|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Hospital Course|8188,8198|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|Hospital Course|8199,8211|false|false|false|C0016053|Fibromyalgia|fibromyalgia
Event|Event|Hospital Course|8199,8211|false|false|false|||fibromyalgia
Drug|Organic Chemical|Hospital Course|8213,8222|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|8213,8222|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|8213,8222|false|false|false|||lorazepam
Drug|Pharmacologic Substance|Hospital Course|8227,8235|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|8227,8235|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|8227,8235|false|false|false|C0917801|Sleeplessness|Insomnia
Drug|Organic Chemical|Hospital Course|8237,8245|false|false|false|C0078839|zolpidem|zolpidem
Drug|Pharmacologic Substance|Hospital Course|8237,8245|false|false|false|C0078839|zolpidem|zolpidem
Event|Event|Hospital Course|8237,8245|false|false|false|||zolpidem
Finding|Idea or Concept|Hospital Course|8265,8268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8265,8268|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|8280,8290|false|false|false|||tolerating
Finding|Daily or Recreational Activity|Hospital Course|8293,8305|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|8301,8305|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|8301,8305|false|false|false|||diet
Finding|Functional Concept|Hospital Course|8301,8305|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|8301,8305|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|8308,8318|false|false|false|||ambulating
Attribute|Clinical Attribute|Hospital Course|8338,8342|false|false|false|C2598155||pain
Event|Event|Hospital Course|8338,8342|false|false|false|||pain
Finding|Functional Concept|Hospital Course|8338,8342|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8338,8342|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|8347,8357|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|8363,8367|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8363,8367|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8363,8367|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8363,8367|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Attribute|Clinical Attribute|Hospital Course|8369,8380|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|8369,8380|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Hospital Course|8369,8380|false|false|false|||medications
Finding|Intellectual Product|Hospital Course|8369,8380|false|false|false|C4284232|Medications|medications
Event|Event|Hospital Course|8406,8410|false|false|false|||home
Finding|Idea or Concept|Hospital Course|8406,8410|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8406,8410|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8406,8410|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|Hospital Course|8414,8420|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|8421,8430|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|8421,8430|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|8421,8430|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|8421,8430|false|false|false|C1705253|Logical Condition|condition
Event|Event|Hospital Course|8437,8447|false|false|false|||outpatient
Finding|Classification|Hospital Course|8437,8447|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|8437,8447|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|8448,8454|false|false|false|||follow
Finding|Functional Concept|Hospital Course|8448,8454|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|8448,8454|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|8448,8457|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|8448,8457|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|8458,8467|false|false|false|||scheduled
Event|Event|Hospital Course|8482,8491|false|false|false|||scheduled
Event|Activity|Hospital Course|8504,8515|false|false|false|C0003629|Appointments|appointment
Event|Event|Hospital Course|8504,8515|false|false|false|||appointment
Event|Event|Hospital Course|8521,8528|false|false|false|||Allergy
Finding|Finding|Hospital Course|8521,8528|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Idea or Concept|Hospital Course|8521,8528|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Pathologic Function|Hospital Course|8521,8528|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Finding|Physiologic Function|Hospital Course|8521,8528|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|Allergy
Event|Event|Hospital Course|8533,8543|false|false|false|||Immunology
Finding|Intellectual Product|Hospital Course|8533,8543|false|false|false|C1547987|Diagnostic Service Section ID - Immunology|Immunology
Attribute|Clinical Attribute|Hospital Course|8548,8559|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8548,8559|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|8548,8559|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|8548,8559|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8548,8572|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|8563,8572|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|8563,8572|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|8574,8583|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8574,8583|false|false|false|C0001927|albuterol|Albuterol
Drug|Organic Chemical|Hospital Course|8574,8591|false|false|false|C0543495|albuterol sulfate|Albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|8574,8591|false|false|false|C0543495|albuterol sulfate|Albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8584,8591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|8584,8591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|8584,8591|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|8584,8591|false|false|false|||sulfate
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8614,8617|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|8614,8617|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|8614,8617|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|8614,8617|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|8614,8617|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Event|Event|Hospital Course|8622,8625|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|8622,8625|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8626,8635|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|8626,8635|false|false|false|C0001927|albuterol|Albuterol
Drug|Organic Chemical|Hospital Course|8636,8642|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|8636,8642|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|8636,8646|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|8636,8646|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|8643,8646|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Hospital Course|8643,8646|false|false|false|||HFA
Procedure|Diagnostic Procedure|Hospital Course|8643,8646|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|8654,8657|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|8654,8657|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|8654,8657|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|8654,8657|false|false|false|||INH
Finding|Functional Concept|Hospital Course|8654,8657|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8665,8668|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8665,8668|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8665,8668|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8665,8668|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8665,8668|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|8669,8672|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|8669,8672|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Antibiotic|Hospital Course|8674,8684|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Organic Chemical|Hospital Course|8674,8684|false|false|false|C0007716|cephalexin|Cephalexin
Drug|Organic Chemical|Hospital Course|8696,8704|false|false|false|C0290795|Adderall|Adderall
Drug|Pharmacologic Substance|Hospital Course|8696,8704|false|false|false|C0290795|Adderall|Adderall
Event|Event|Hospital Course|8696,8704|false|false|false|||Adderall
Drug|Organic Chemical|Hospital Course|8696,8707|false|false|false|C1170024|Adderall-XR|Adderall XR
Drug|Pharmacologic Substance|Hospital Course|8696,8707|false|false|false|C1170024|Adderall-XR|Adderall XR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8714,8717|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8714,8717|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8714,8717|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8714,8717|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8714,8717|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8718,8732|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|Ergocalciferol
Drug|Pharmacologic Substance|Hospital Course|8718,8732|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|Ergocalciferol
Drug|Vitamin|Hospital Course|8718,8732|false|false|false|C0014695;C3714696|Ergocalciferol Drug Product;ergocalciferol|Ergocalciferol
Event|Event|Hospital Course|8718,8732|false|false|false|||Ergocalciferol
Drug|Organic Chemical|Hospital Course|8718,8745|false|false|false|C0014695|ergocalciferol|Ergocalciferol (vitamin D2)
Drug|Pharmacologic Substance|Hospital Course|8718,8745|false|false|false|C0014695|ergocalciferol|Ergocalciferol (vitamin D2)
Drug|Vitamin|Hospital Course|8718,8745|false|false|false|C0014695|ergocalciferol|Ergocalciferol (vitamin D2)
Drug|Organic Chemical|Hospital Course|8734,8741|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|8734,8741|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|8734,8741|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|Hospital Course|8734,8744|false|false|false|C0014695|ergocalciferol|vitamin D2
Drug|Pharmacologic Substance|Hospital Course|8734,8744|false|false|false|C0014695|ergocalciferol|vitamin D2
Drug|Vitamin|Hospital Course|8734,8744|false|false|false|C0014695|ergocalciferol|vitamin D2
Event|Event|Hospital Course|8734,8744|false|false|false|||vitamin D2
Finding|Intellectual Product|Hospital Course|8757,8761|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|Hospital Course|8762,8768|false|false|false|C0939400|Nexium|Nexium
Drug|Pharmacologic Substance|Hospital Course|8762,8768|false|false|false|C0939400|Nexium|Nexium
Event|Event|Hospital Course|8762,8768|false|false|false|||Nexium
Event|Event|Hospital Course|8779,8782|false|false|false|||QAM
Drug|Hormone|Hospital Course|8783,8790|false|false|false|C0724374|Vivelle|Vivelle
Drug|Organic Chemical|Hospital Course|8783,8790|false|false|false|C0724374|Vivelle|Vivelle
Drug|Pharmacologic Substance|Hospital Course|8783,8790|false|false|false|C0724374|Vivelle|Vivelle
Drug|Biomedical or Dental Material|Hospital Course|8816,8821|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|8816,8821|false|false|false|||Patch
Finding|Finding|Hospital Course|8816,8821|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Intellectual Product|Hospital Course|8827,8831|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|Hospital Course|8833,8841|false|false|false|C0699601|Diflucan|Diflucan
Drug|Pharmacologic Substance|Hospital Course|8833,8841|false|false|false|C0699601|Diflucan|Diflucan
Drug|Organic Chemical|Hospital Course|8856,8867|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Drug|Pharmacologic Substance|Hospital Course|8856,8867|false|false|false|C0020404|hydroxyzine|Hydroxyzine
Drug|Organic Chemical|Hospital Course|8856,8871|false|false|false|C0600110|hydroxyzine hydrochloride|Hydroxyzine HCl
Drug|Pharmacologic Substance|Hospital Course|8856,8871|false|false|false|C0600110|hydroxyzine hydrochloride|Hydroxyzine HCl
Disorder|Neoplastic Process|Hospital Course|8868,8871|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|8868,8871|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|8868,8871|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|8868,8871|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|8868,8871|false|false|false|||HCl
Event|Event|Hospital Course|8881,8884|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|8881,8884|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8886,8895|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Hospital Course|8886,8895|false|false|false|C0020740|ibuprofen|Ibuprofen
Event|Event|Hospital Course|8907,8910|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|8907,8910|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8911,8918|false|false|false|C3496839|Linzess|Linzess
Drug|Pharmacologic Substance|Hospital Course|8911,8918|false|false|false|C3496839|Linzess|Linzess
Drug|Organic Chemical|Hospital Course|8944,8950|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|Hospital Course|8944,8950|false|false|false|C0699194|Ativan|Ativan
Event|Event|Hospital Course|8959,8962|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|8959,8962|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|8964,8974|false|false|false|C0025854|metolazone|Metolazone
Drug|Pharmacologic Substance|Hospital Course|8964,8974|false|false|false|C0025854|metolazone|Metolazone
Drug|Organic Chemical|Hospital Course|8985,8991|false|false|false|C0206046|Zofran|Zofran
Drug|Pharmacologic Substance|Hospital Course|8985,8991|false|false|false|C0206046|Zofran|Zofran
Event|Event|Hospital Course|9000,9003|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|9000,9003|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|9005,9014|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Hospital Course|9005,9014|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Hospital Course|9005,9014|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Hospital Course|9005,9014|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Event|Event|Hospital Course|9027,9030|false|false|false|||PRN
Finding|Gene or Genome|Hospital Course|9027,9030|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Biologically Active Substance|Hospital Course|9032,9041|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|9032,9041|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|9032,9041|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|9032,9041|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|9032,9041|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|9032,9041|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|9032,9041|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|9032,9041|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|9032,9050|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Pharmacologic Substance|Hospital Course|9032,9050|false|false|false|C0032825|potassium chloride|Potassium chloride
Drug|Element, Ion, or Isotope|Hospital Course|9042,9050|false|false|false|C0008203;C0596019|Chlorides;chloride ion|chloride
Event|Event|Hospital Course|9042,9050|false|false|false|||chloride
Finding|Physiologic Function|Hospital Course|9042,9050|false|false|false|C4553021|Chloride metabolic function|chloride
Procedure|Laboratory Procedure|Hospital Course|9042,9050|false|false|false|C0201952|Chloride measurement|chloride
Anatomy|Body Space or Junction|Hospital Course|9056,9060|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|9056,9060|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|9056,9060|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|9056,9060|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biomedical or Dental Material|Hospital Course|9056,9067|false|false|false|C1273619|Oral Liquid Product|Oral Liquid
Drug|Biomedical or Dental Material|Hospital Course|9061,9067|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|Hospital Course|9061,9067|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|Hospital Course|9061,9067|false|false|false|||Liquid
Finding|Finding|Hospital Course|9061,9067|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9061,9067|false|false|false|C0301571|Liquid diet|Liquid
Drug|Organic Chemical|Hospital Course|9080,9091|false|false|false|C0033497|propranolol|Propranolol
Drug|Pharmacologic Substance|Hospital Course|9080,9091|false|false|false|C0033497|propranolol|Propranolol
Event|Event|Hospital Course|9104,9107|false|false|false|||QHS
Drug|Organic Chemical|Hospital Course|9108,9122|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|Hospital Course|9108,9122|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Antibiotic|Hospital Course|9133,9145|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|9133,9145|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|Hospital Course|9153,9159|false|false|false|C0039225|Tablet Dosage Form|tablet
Drug|Organic Chemical|Hospital Course|9163,9169|false|false|false|C0487782|Ambien|Ambien
Drug|Pharmacologic Substance|Hospital Course|9163,9169|false|false|false|C0487782|Ambien|Ambien
Event|Event|Hospital Course|9188,9196|false|false|false|||catheter
Finding|Intellectual Product|Hospital Course|9188,9196|false|false|false|C1546572||catheter
Drug|Organic Chemical|Hospital Course|9198,9206|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9198,9206|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|9198,9213|false|false|false|C0243237|docusate sodium|Docusate sodium
Drug|Pharmacologic Substance|Hospital Course|9198,9213|false|false|false|C0243237|docusate sodium|Docusate sodium
Drug|Biologically Active Substance|Hospital Course|9207,9213|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|9207,9213|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|9207,9213|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|9207,9213|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|9207,9213|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|9207,9213|false|false|false|C0337443|Sodium measurement|sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9221,9224|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9221,9224|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9221,9224|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9221,9224|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9221,9224|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|9239,9250|false|false|false|C3811910|combination - answer to question|COMBINATION
Event|Event|Hospital Course|9253,9262|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9253,9262|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9253,9262|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9253,9262|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9253,9262|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9253,9274|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9263,9274|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9263,9274|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9263,9274|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9263,9274|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9279,9287|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9279,9287|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|9279,9294|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|9279,9294|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|9288,9294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9288,9294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9288,9294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|9288,9294|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|9288,9294|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9288,9294|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Biomedical or Dental Material|Hospital Course|9296,9302|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Drug|Substance|Hospital Course|9296,9302|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|Liquid
Event|Event|Hospital Course|9296,9302|false|false|false|||Liquid
Finding|Finding|Hospital Course|9296,9302|false|false|false|C1304698|Liquid (finding)|Liquid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9296,9302|false|false|false|C0301571|Liquid diet|Liquid
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9314,9317|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9314,9317|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9314,9317|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9314,9317|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9314,9317|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9323,9331|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|9323,9331|false|false|false|C1692318|docusate|docusate
Drug|Organic Chemical|Hospital Course|9323,9338|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|9323,9338|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|9332,9338|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|9332,9338|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|9332,9338|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|9332,9338|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|9332,9338|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|9332,9338|false|false|false|C0337443|Sodium measurement|sodium
Drug|Biomedical or Dental Material|Hospital Course|9348,9354|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|9348,9354|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|9355,9363|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9358,9363|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9358,9363|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Hospital Course|9372,9375|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|9372,9375|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|9376,9380|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|9376,9380|false|false|false|C2828567|PRSS30P gene|Disp
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9387,9394|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|9387,9394|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|9387,9394|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Hospital Course|9395,9402|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9395,9402|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9409,9418|false|false|false|C0005632|bisacodyl|Bisacodyl
Drug|Pharmacologic Substance|Hospital Course|9409,9418|false|false|false|C0005632|bisacodyl|Bisacodyl
Finding|Gene or Genome|Hospital Course|9437,9440|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9441,9453|false|false|false|||Constipation
Finding|Sign or Symptom|Hospital Course|9441,9453|false|false|false|C0009806|Constipation|Constipation
Event|Event|Hospital Course|9455,9457|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|9459,9468|false|false|false|C0005632|bisacodyl|bisacodyl
Drug|Pharmacologic Substance|Hospital Course|9459,9468|false|false|false|C0005632|bisacodyl|bisacodyl
Drug|Biomedical or Dental Material|Hospital Course|9478,9484|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|9478,9484|false|false|false|||tablet
Event|Event|Hospital Course|9485,9492|false|false|false|||delayed
Event|Event|Hospital Course|9493,9500|false|false|false|||release
Finding|Functional Concept|Hospital Course|9493,9500|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|release
Procedure|Health Care Activity|Hospital Course|9493,9500|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9493,9500|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|release
Anatomy|Body Location or Region|Hospital Course|9511,9516|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9511,9516|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|9517,9529|false|false|false|||constipation
Finding|Sign or Symptom|Hospital Course|9517,9529|false|false|false|C0009806|Constipation|constipation
Drug|Biomedical or Dental Material|Hospital Course|9540,9546|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9547,9554|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9547,9554|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9561,9571|false|false|false|C0025854|metolazone|Metolazone
Drug|Pharmacologic Substance|Hospital Course|9561,9571|false|false|false|C0025854|metolazone|Metolazone
Drug|Organic Chemical|Hospital Course|9592,9598|false|false|false|C0939400|Nexium|NexIUM
Drug|Pharmacologic Substance|Hospital Course|9592,9598|false|false|false|C0939400|Nexium|NexIUM
Event|Event|Hospital Course|9592,9598|false|false|false|||NexIUM
Drug|Organic Chemical|Hospital Course|9600,9612|false|false|false|C0937846|esomeprazole|esomeprazole
Drug|Pharmacologic Substance|Hospital Course|9600,9612|false|false|false|C0937846|esomeprazole|esomeprazole
Drug|Organic Chemical|Hospital Course|9600,9622|false|false|false|C0937622|esomeprazole magnesium|esomeprazole magnesium
Drug|Pharmacologic Substance|Hospital Course|9600,9622|false|false|false|C0937622|esomeprazole magnesium|esomeprazole magnesium
Drug|Biologically Active Substance|Hospital Course|9613,9622|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Element, Ion, or Isotope|Hospital Course|9613,9622|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Inorganic Chemical|Hospital Course|9613,9622|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Drug|Pharmacologic Substance|Hospital Course|9613,9622|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|magnesium
Event|Event|Hospital Course|9613,9622|false|false|false|||magnesium
Procedure|Laboratory Procedure|Hospital Course|9613,9622|false|false|false|C0373675|Magnesium measurement|magnesium
Anatomy|Body Space or Junction|Hospital Course|9630,9634|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|Hospital Course|9630,9634|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|Hospital Course|9630,9634|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|Hospital Course|9630,9634|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Intellectual Product|Hospital Course|9635,9639|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|9640,9648|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|9640,9648|false|false|false|||Duration
Drug|Organic Chemical|Hospital Course|9662,9671|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|9662,9671|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|9662,9671|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|9662,9671|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|9673,9682|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|9673,9682|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|9673,9690|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|9683,9690|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9683,9690|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9683,9690|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9683,9690|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|9707,9710|true|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9711,9715|true|false|false|C2598155||pain
Event|Event|Hospital Course|9711,9715|true|false|false|||pain
Finding|Functional Concept|Hospital Course|9711,9715|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9711,9715|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9724,9729|true|false|false|||drive
Event|Event|Hospital Course|9734,9739|true|false|false|||drink
Drug|Pharmacologic Substance|Hospital Course|9748,9758|true|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|9748,9758|true|false|false|||medication
Finding|Intellectual Product|Hospital Course|9748,9758|true|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|9760,9762|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|9764,9773|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|9764,9773|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|9764,9773|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|9764,9773|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|9783,9789|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|9783,9789|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|9793,9801|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9796,9801|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9796,9801|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|9810,9813|false|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9810,9813|false|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|Hospital Course|9810,9813|false|false|false|C1568891|HGS protein, human|hrs
Event|Event|Hospital Course|9810,9813|false|false|false|||hrs
Finding|Gene or Genome|Hospital Course|9810,9813|false|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Drug|Biomedical or Dental Material|Hospital Course|9825,9831|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|9832,9839|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|9832,9839|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9846,9857|false|false|false|C0033497|propranolol|Propranolol
Drug|Pharmacologic Substance|Hospital Course|9846,9857|false|false|false|C0033497|propranolol|Propranolol
Event|Event|Hospital Course|9846,9857|false|false|false|||Propranolol
Drug|Organic Chemical|Hospital Course|9880,9894|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|Hospital Course|9880,9894|false|false|false|C0037982|spironolactone|Spironolactone
Event|Event|Hospital Course|9880,9894|false|false|false|||Spironolactone
Drug|Organic Chemical|Hospital Course|9915,9923|false|false|false|C0078839|zolpidem|Zolpidem
Drug|Pharmacologic Substance|Hospital Course|9915,9923|false|false|false|C0078839|zolpidem|Zolpidem
Drug|Organic Chemical|Hospital Course|9915,9932|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Pharmacologic Substance|Hospital Course|9915,9932|false|false|false|C0724725|zolpidem tartrate|Zolpidem Tartrate
Drug|Organic Chemical|Hospital Course|9924,9932|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|9924,9932|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|Hospital Course|9924,9932|false|false|false|||Tartrate
Drug|Antibiotic|Hospital Course|9948,9960|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|Hospital Course|9948,9960|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Hormone|Hospital Course|9982,9989|false|false|false|C0724374|Vivelle|Vivelle
Drug|Organic Chemical|Hospital Course|9982,9989|false|false|false|C0724374|Vivelle|Vivelle
Drug|Pharmacologic Substance|Hospital Course|9982,9989|false|false|false|C0724374|Vivelle|Vivelle
Drug|Hormone|Hospital Course|9991,10000|false|false|false|C0014912|estradiol|estradiol
Drug|Organic Chemical|Hospital Course|9991,10000|false|false|false|C0014912|estradiol|estradiol
Drug|Pharmacologic Substance|Hospital Course|9991,10000|false|false|false|C0014912|estradiol|estradiol
Event|Event|Hospital Course|9991,10000|false|false|false|||estradiol
Procedure|Laboratory Procedure|Hospital Course|9991,10000|false|false|false|C0337434|Estradiol measurement|estradiol
Event|Event|Hospital Course|10017,10028|false|false|false|||Transdermal
Finding|Finding|Hospital Course|10017,10028|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Finding|Functional Concept|Hospital Course|10017,10028|false|false|false|C0040652;C0694643;C4521342|Transdermal (intended site);Transdermal Route of Administration;transdermal|Transdermal
Finding|Intellectual Product|Hospital Course|10035,10039|false|false|false|C1561540|Transaction counts and value totals - week|week
Drug|Organic Chemical|Hospital Course|10045,10054|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|10045,10054|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|10069,10072|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10073,10080|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|10073,10080|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|10073,10080|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Biologically Active Substance|Hospital Course|10086,10095|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|10086,10095|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|10086,10095|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|10086,10095|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|10086,10095|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|10086,10095|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|10086,10095|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|10086,10095|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Inorganic Chemical|Hospital Course|10086,10104|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Pharmacologic Substance|Hospital Course|10086,10104|false|false|false|C0032825|potassium chloride|Potassium Chloride
Drug|Element, Ion, or Isotope|Hospital Course|10096,10104|false|false|false|C0008203;C0596019|Chlorides;chloride ion|Chloride
Event|Event|Hospital Course|10096,10104|false|false|false|||Chloride
Finding|Physiologic Function|Hospital Course|10096,10104|false|false|false|C4553021|Chloride metabolic function|Chloride
Procedure|Laboratory Procedure|Hospital Course|10096,10104|false|false|false|C0201952|Chloride measurement|Chloride
Event|Event|Hospital Course|10108,10111|false|false|false|||mEq
Drug|Pharmacologic Substance|Hospital Course|10121,10129|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|10121,10129|false|false|false|||Duration
Event|Activity|Hospital Course|10141,10145|false|false|false|C1948035|Hold (action)|Hold
Event|Event|Hospital Course|10141,10145|false|false|false|||Hold
Finding|Functional Concept|Hospital Course|10141,10145|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|Hold
Finding|Intellectual Product|Hospital Course|10141,10145|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|Hold
Event|Event|Hospital Course|10158,10167|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10158,10167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10158,10167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10158,10167|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10158,10167|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10158,10179|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10158,10179|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10168,10179|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|10168,10179|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|10168,10179|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|10181,10185|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|10181,10185|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|10181,10185|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|10181,10185|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|10188,10197|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10188,10197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10188,10197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10188,10197|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10188,10197|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|10188,10207|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|10198,10207|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|10198,10207|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|10198,10207|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10198,10207|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10198,10207|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10209,10216|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|Hospital Course|10209,10226|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|Hospital Course|10209,10226|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|Hospital Course|10217,10226|false|false|false|C1318143|Retention - dental|retention
Event|Event|Hospital Course|10217,10226|false|false|false|||retention
Finding|Cell Function|Hospital Course|10217,10226|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|Hospital Course|10217,10226|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|Hospital Course|10217,10226|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Disorder|Acquired Abnormality|Hospital Course|10228,10237|false|false|false|C0149771|Rectocele|rectocele
Event|Event|Hospital Course|10228,10237|false|false|false|||rectocele
Finding|Mental Process|Discharge Condition|10262,10268|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10262,10275|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10262,10275|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10269,10275|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10269,10275|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10277,10282|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|10277,10282|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|10287,10295|false|false|false|||coherent
Finding|Finding|Discharge Condition|10287,10295|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|10297,10302|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|10297,10319|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|10297,10319|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|10306,10319|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|10306,10319|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|10306,10319|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|10321,10326|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|10321,10326|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|10321,10326|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|10321,10326|false|false|false|||Alert
Finding|Finding|Discharge Condition|10321,10326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|10321,10326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|10321,10326|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|10331,10342|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|10331,10342|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|10344,10352|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|10344,10352|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|10344,10352|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|10353,10359|false|false|false|C5889824||Status
Event|Event|Discharge Condition|10353,10359|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|10353,10359|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10361,10371|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|10361,10371|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|10361,10371|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|10361,10371|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|10361,10371|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|10374,10385|false|false|false|||Independent
Finding|Finding|Discharge Condition|10374,10385|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|10374,10385|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|10414,10418|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|10434,10442|false|false|false|||admitted
Event|Occupational Activity|Discharge Instructions|10461,10468|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Discharge Instructions|10461,10468|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Discharge Instructions|10480,10489|false|false|false|||scheduled
Attribute|Clinical Attribute|Discharge Instructions|10491,10496|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Discharge Instructions|10491,10498|false|false|false|C0441767|Stage level 2|Stage 2
Event|Event|Discharge Instructions|10510,10519|false|false|false|||placement
Procedure|Health Care Activity|Discharge Instructions|10510,10519|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10510,10519|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Disorder|Disease or Syndrome|Discharge Instructions|10524,10533|false|false|false|C0751438|Posterior pituitary disease|posterior
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10524,10546|false|false|false|C0195230;C5574717|Posterior repair of vagina;Repair of rectocele|posterior colporrhaphy
Event|Event|Discharge Instructions|10534,10546|false|false|false|||colporrhaphy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10534,10546|false|false|false|C0009416|Suture of vagina|colporrhaphy
Anatomy|Tissue|Discharge Instructions|10553,10558|false|false|false|C0332835|Transplanted tissue|graft
Drug|Biomedical or Dental Material|Discharge Instructions|10553,10558|false|false|false|C0181074;C1705210|Graft Dosage Form;Graft material|graft
Event|Event|Discharge Instructions|10553,10558|false|false|false|||graft
Finding|Intellectual Product|Discharge Instructions|10553,10558|false|false|false|C1546653|Graft - Specimen Source Codes|graft
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10553,10558|false|false|false|C1961139;C3683798|Graft Procedures on the Head;Grafting procedure|graft
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10563,10570|false|false|false|C0042027|Urinary tract|urinary
Attribute|Clinical Attribute|Discharge Instructions|10563,10580|false|false|false|C5700171|Bladder retention of urine|urinary retention
Finding|Functional Concept|Discharge Instructions|10563,10580|false|false|false|C0080274|Urinary Retention|urinary retention
Attribute|Clinical Attribute|Discharge Instructions|10571,10580|false|false|false|C1318143|Retention - dental|retention
Event|Event|Discharge Instructions|10571,10580|false|false|false|||retention
Finding|Cell Function|Discharge Instructions|10571,10580|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Functional Concept|Discharge Instructions|10571,10580|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Finding|Mental Process|Discharge Instructions|10571,10580|false|false|false|C0035280;C0080274;C0333117;C1753315|Retention (Psychology);Retention of content;Urinary Retention;cellular entity retention|retention
Disorder|Acquired Abnormality|Discharge Instructions|10585,10594|false|false|false|C0149771|Rectocele|rectocele
Event|Event|Discharge Instructions|10585,10594|false|false|false|||rectocele
Disorder|Anatomical Abnormality|Discharge Instructions|10599,10609|false|false|false|C0205792|Enterocele|enterocele
Event|Event|Discharge Instructions|10599,10609|false|false|false|||enterocele
Event|Event|Discharge Instructions|10617,10626|false|false|false|||tolerated
Attribute|Clinical Attribute|Discharge Instructions|10631,10640|false|false|false|C0945766||procedure
Event|Event|Discharge Instructions|10631,10640|false|false|false|||procedure
Event|Occupational Activity|Discharge Instructions|10631,10640|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Discharge Instructions|10631,10640|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10631,10640|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|Discharge Instructions|10641,10645|false|false|false|C5575035|Well (answer to question)|well
Event|Activity|Discharge Instructions|10667,10676|false|false|false|C3241922|Operation Activity|operation
Event|Event|Discharge Instructions|10667,10676|false|false|false|||operation
Procedure|Machine Activity|Discharge Instructions|10667,10676|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10667,10676|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Finding|Finding|Discharge Instructions|10689,10695|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|10689,10695|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Discharge Instructions|10689,10713|false|false|false|C2220378|severe allergic reaction|severe allergic reaction
Finding|Functional Concept|Discharge Instructions|10696,10704|false|false|false|C0700624|Allergic|allergic
Finding|Pathologic Function|Discharge Instructions|10696,10713|false|false|false|C0020517;C1527304|Allergic Reaction;Hypersensitivity|allergic reaction
Event|Event|Discharge Instructions|10705,10713|false|false|false|||reaction
Finding|Functional Concept|Discharge Instructions|10705,10713|false|false|false|C0443286|Reaction|reaction
Anatomy|Body Space or Junction|Discharge Instructions|10736,10739|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|Discharge Instructions|10736,10739|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Event|Activity|Discharge Instructions|10745,10755|false|false|false|C1283169||monitoring
Event|Event|Discharge Instructions|10745,10755|false|false|false|||monitoring
Procedure|Health Care Activity|Discharge Instructions|10745,10755|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Intellectual Product|Discharge Instructions|10763,10767|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Discharge Instructions|10778,10787|false|false|false|||recovered
Finding|Finding|Discharge Instructions|10788,10792|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|10807,10817|false|false|false|||determined
Finding|Intellectual Product|Discharge Instructions|10834,10840|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Discharge Instructions|10841,10850|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|10841,10850|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|10841,10850|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|10841,10850|false|false|false|C1705253|Logical Condition|condition
Event|Event|Discharge Instructions|10855,10864|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|10855,10864|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|10855,10864|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|10855,10864|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|10855,10864|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Discharge Instructions|10874,10878|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|10884,10894|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|10884,10894|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|10884,10894|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|10899,10905|false|false|false|||follow
Event|Activity|Discharge Instructions|10917,10929|false|false|false|C0003629|Appointments|appointments
Event|Event|Discharge Instructions|10917,10929|false|false|false|||appointments
Event|Event|Discharge Instructions|10934,10943|false|false|false|||scheduled
Attribute|Clinical Attribute|Discharge Instructions|10950,10962|false|false|false|C3263700||instructions
Event|Event|Discharge Instructions|10950,10962|false|false|false|||instructions
Finding|Intellectual Product|Discharge Instructions|10950,10962|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Attribute|Clinical Attribute|Discharge Instructions|10978,10989|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|10978,10989|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|10978,10989|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|10978,10989|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|10993,11003|false|false|false|||prescribed
Event|Event|Discharge Instructions|11016,11021|true|false|false|||drive
Drug|Hazardous or Poisonous Substance|Discharge Instructions|11035,11044|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Discharge Instructions|11035,11044|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Discharge Instructions|11035,11044|false|false|false|||narcotics
Finding|Body Substance|Discharge Instructions|11056,11061|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|11056,11070|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|11056,11070|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|11062,11070|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|11079,11085|false|false|false|C0282139|Colace|colace
Drug|Pharmacologic Substance|Discharge Instructions|11079,11085|false|false|false|C0282139|Colace|colace
Event|Event|Discharge Instructions|11079,11085|false|false|false|||colace
Drug|Hazardous or Poisonous Substance|Discharge Instructions|11099,11108|false|false|false|C0027415|Narcotics|narcotics
Drug|Pharmacologic Substance|Discharge Instructions|11099,11108|false|false|false|C0027415|Narcotics|narcotics
Event|Event|Discharge Instructions|11099,11108|false|false|false|||narcotics
Event|Event|Discharge Instructions|11121,11133|true|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|11121,11133|true|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|11144,11151|true|false|false|||combine
Drug|Hazardous or Poisonous Substance|Discharge Instructions|11152,11160|true|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|11152,11160|true|false|false|C0027415|Narcotics|narcotic
Event|Event|Discharge Instructions|11152,11160|true|false|false|||narcotic
Drug|Pharmacologic Substance|Discharge Instructions|11165,11173|true|false|false|C0036557|Sedatives|sedative
Attribute|Clinical Attribute|Discharge Instructions|11174,11185|true|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|11174,11185|true|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|11174,11185|true|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|11174,11185|true|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Discharge Instructions|11189,11196|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|11189,11196|true|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|Discharge Instructions|11189,11196|true|false|false|||alcohol
Finding|Intellectual Product|Discharge Instructions|11189,11196|true|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|Discharge Instructions|11208,11212|true|false|false|||take
Drug|Organic Chemical|Discharge Instructions|11230,11243|true|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Discharge Instructions|11230,11243|true|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Discharge Instructions|11230,11243|true|false|false|||acetaminophen
Procedure|Laboratory Procedure|Discharge Instructions|11230,11243|true|false|false|C0373527|Acetaminophen measurement|acetaminophen
Disorder|Disease or Syndrome|Discharge Instructions|11245,11249|true|false|false|C1970472|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED|APAP
Drug|Organic Chemical|Discharge Instructions|11245,11249|true|false|false|C0000970|acetaminophen|APAP
Drug|Pharmacologic Substance|Discharge Instructions|11245,11249|true|false|false|C0000970|acetaminophen|APAP
Event|Event|Discharge Instructions|11245,11249|true|false|false|||APAP
Disorder|Disease or Syndrome|Discharge Instructions|11257,11260|true|false|false|C0751781|Dentatorubral-Pallidoluysian Atrophy|hrs
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|11257,11260|true|false|false|C1568891|HGS protein, human|hrs
Drug|Biologically Active Substance|Discharge Instructions|11257,11260|true|false|false|C1568891|HGS protein, human|hrs
Event|Event|Discharge Instructions|11257,11260|true|false|false|||hrs
Finding|Gene or Genome|Discharge Instructions|11257,11260|true|false|false|C1366514;C1415473;C1419996;C1708271;C5575450;C5780798|ATN1 wt Allele;HARS1 gene;HARS1 wt Allele;HGS gene;HGS wt Allele;SRSF5 gene|hrs
Finding|Daily or Recreational Activity|Discharge Instructions|11268,11286|true|false|false|C1514989|Strenuous Exercise|strenuous activity
Event|Activity|Discharge Instructions|11278,11286|true|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|11278,11286|true|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|11278,11286|true|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|11278,11286|true|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Activity|Discharge Instructions|11306,11317|true|false|false|C0003629|Appointments|appointment
Event|Event|Discharge Instructions|11306,11317|true|false|false|||appointment
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11337,11343|true|false|false|C0042232;C1519910;C4482396|Mouse Vagina;Pelvis>Vagina;Vagina|vagina
Anatomy|Tissue|Discharge Instructions|11337,11343|true|false|false|C0042232;C1519910;C4482396|Mouse Vagina;Pelvis>Vagina;Vagina|vagina
Disorder|Disease or Syndrome|Discharge Instructions|11337,11343|true|false|false|C0042251;C0154002;C0686277|Benign neoplasm vagina;Carcinoma in situ of vagina;Vaginal Diseases|vagina
Disorder|Neoplastic Process|Discharge Instructions|11337,11343|true|false|false|C0042251;C0154002;C0686277|Benign neoplasm vagina;Carcinoma in situ of vagina;Vaginal Diseases|vagina
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11337,11343|true|false|false|C0869896|Procedure on vagina|vagina
Event|Event|Discharge Instructions|11348,11355|true|false|false|||tampons
Event|Event|Discharge Instructions|11360,11368|true|false|false|||douching
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11360,11368|true|false|false|C2936784|Douching procedure|douching
Attribute|Clinical Attribute|Discharge Instructions|11373,11376|true|false|false|C0804628||sex
Finding|Behavior|Discharge Instructions|11373,11376|true|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|sex
Finding|Finding|Discharge Instructions|11373,11376|true|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|sex
Finding|Gene or Genome|Discharge Instructions|11373,11376|true|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|sex
Finding|Organism Function|Discharge Instructions|11373,11376|true|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|sex
Event|Activity|Discharge Instructions|11402,11409|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|11402,11409|true|false|false|||lifting
Event|Event|Discharge Instructions|11413,11420|true|false|false|||objects
Event|Event|Discharge Instructions|11455,11458|false|false|false|||eat
Finding|Daily or Recreational Activity|Discharge Instructions|11461,11473|false|false|false|C0184625||regular diet
Drug|Food|Discharge Instructions|11469,11473|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Discharge Instructions|11469,11473|false|false|false|||diet
Finding|Functional Concept|Discharge Instructions|11469,11473|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Discharge Instructions|11469,11473|false|false|false|C0012159|Diet therapy|diet
Event|Event|Discharge Instructions|11481,11489|false|false|false|||anything
Anatomy|Body Location or Region|Discharge Instructions|11509,11517|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|Discharge Instructions|11509,11517|false|false|false|C0332803|Surgical wound|Incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11509,11517|false|false|false|C0184898|Surgical incisions|Incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11509,11522|false|false|false|C0150258|Incision care|Incision care
Event|Activity|Discharge Instructions|11518,11522|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|11518,11522|false|false|false|||care
Finding|Finding|Discharge Instructions|11518,11522|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11518,11522|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|11536,11542|false|false|false|||shower
Event|Event|Discharge Instructions|11547,11552|false|false|false|||allow
Drug|Inorganic Chemical|Discharge Instructions|11559,11564|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|Discharge Instructions|11559,11564|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|Discharge Instructions|11559,11564|false|false|false|||water
Finding|Intellectual Product|Discharge Instructions|11559,11564|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11559,11564|false|false|false|C0020311|Hydrotherapy|water
Event|Event|Discharge Instructions|11568,11571|false|false|false|||run
Finding|Daily or Recreational Activity|Discharge Instructions|11568,11571|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Finding|Discharge Instructions|11568,11571|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Functional Concept|Discharge Instructions|11568,11571|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Finding|Intellectual Product|Discharge Instructions|11568,11571|false|false|false|C0035953;C0600140;C1704688;C4722187|Does run (finding);Go Jogging or Running Question;Run action;Running (physical activity)|run
Anatomy|Body Location or Region|Discharge Instructions|11577,11585|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|11577,11585|false|true|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|11577,11585|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11577,11585|false|true|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|Discharge Instructions|11604,11612|true|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|11604,11612|true|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|11604,11612|true|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11604,11612|true|false|false|C0184898|Surgical incisions|incision
Procedure|Health Care Activity|Discharge Instructions|11617,11621|true|false|false|C0150141|Bathing|bath
Event|Event|Discharge Instructions|11622,11626|true|false|false|||tubs
Event|Event|Discharge Instructions|11644,11648|false|false|false|||Call
Event|Event|Discharge Instructions|11654,11660|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|11654,11660|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|11670,11675|false|false|false|||fever
Finding|Finding|Discharge Instructions|11670,11675|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|11670,11675|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Finding|Discharge Instructions|11688,11694|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|11688,11694|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Location or Region|Discharge Instructions|11695,11704|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|Discharge Instructions|11695,11709|false|true|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|Discharge Instructions|11705,11709|false|true|false|C2598155||pain
Event|Event|Discharge Instructions|11705,11709|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|11705,11709|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|11705,11709|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|11714,11724|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Discharge Instructions|11725,11734|false|false|false|||urinating
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11739,11746|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Discharge Instructions|11739,11746|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Discharge Instructions|11739,11746|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Discharge Instructions|11739,11746|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Finding|Discharge Instructions|11739,11755|false|false|false|C0578503;C2979982|Abnormal vaginal bleeding;Vaginal Hemorrhage|vaginal bleeding
Finding|Pathologic Function|Discharge Instructions|11739,11755|false|false|false|C0578503;C2979982|Abnormal vaginal bleeding;Vaginal Hemorrhage|vaginal bleeding
Event|Event|Discharge Instructions|11747,11755|false|false|false|||bleeding
Finding|Pathologic Function|Discharge Instructions|11747,11755|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Discharge Instructions|11756,11765|false|false|false|||requiring
Anatomy|Anatomical Structure|Discharge Instructions|11769,11772|false|false|false|C3669270|Strucure of thick cushion of skin|pad
Disorder|Disease or Syndrome|Discharge Instructions|11769,11772|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Disorder|Neoplastic Process|Discharge Instructions|11769,11772|false|false|false|C0332568;C1704436|Pad Mass;Peripheral Arterial Diseases|pad
Drug|Biomedical or Dental Material|Discharge Instructions|11769,11772|false|false|false|C2347441|Pad Dosage Form|pad
Event|Event|Discharge Instructions|11769,11772|false|false|false|||pad
Finding|Gene or Genome|Discharge Instructions|11769,11772|false|false|false|C1425244;C1425478;C3540603|DHX40 gene;PADI4 gene;PADI4 wt Allele|pad
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11769,11772|false|false|false|C3814046|PAD Regimen|pad
Finding|Finding|Discharge Instructions|11780,11788|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Discharge Instructions|11780,11788|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Finding|Discharge Instructions|11780,11806|false|false|false|C0566986|Abnormal Vaginal Discharge|abnormal vaginal discharge
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11789,11796|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Discharge Instructions|11789,11796|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Discharge Instructions|11789,11796|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Discharge Instructions|11789,11796|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Finding|Discharge Instructions|11789,11806|false|false|false|C0227791;C0438692|Vaginal Discharge;Vaginal discharge symptom|vaginal discharge
Finding|Sign or Symptom|Discharge Instructions|11789,11806|false|false|false|C0227791;C0438692|Vaginal Discharge;Vaginal discharge symptom|vaginal discharge
Event|Event|Discharge Instructions|11797,11806|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|11797,11806|false|true|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|11797,11806|false|true|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|11797,11806|false|true|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|11797,11806|false|true|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Discharge Instructions|11811,11818|false|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|11811,11818|false|false|false|||redness
Finding|Finding|Discharge Instructions|11811,11818|false|false|false|C0332575|Redness|redness
Event|Event|Discharge Instructions|11822,11830|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|11822,11830|false|true|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|11822,11830|false|true|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11822,11830|false|true|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|Discharge Instructions|11836,11844|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|11836,11844|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|11836,11844|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11836,11844|false|false|false|C0184898|Surgical incisions|incision
Attribute|Clinical Attribute|Discharge Instructions|11849,11855|false|false|false|C4255480||nausea
Finding|Sign or Symptom|Discharge Instructions|11849,11855|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|Discharge Instructions|11849,11864|false|false|false|C0027498|Nausea and vomiting|nausea/vomiting
Event|Event|Discharge Instructions|11856,11864|false|false|false|||vomiting
Finding|Sign or Symptom|Discharge Instructions|11856,11864|false|false|false|C0042963|Vomiting|vomiting
Event|Event|Discharge Instructions|11879,11885|false|false|false|||unable
Finding|Finding|Discharge Instructions|11879,11885|false|false|false|C1299582|Unable|unable
Event|Event|Discharge Instructions|11889,11893|false|false|false|||keep
Drug|Substance|Discharge Instructions|11899,11905|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|11899,11905|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|11899,11905|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11899,11905|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Food|Discharge Instructions|11906,11910|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|Discharge Instructions|11906,11910|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|Discharge Instructions|11906,11910|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|Discharge Instructions|11906,11910|false|false|false|||food
Drug|Pharmacologic Substance|Discharge Instructions|11920,11930|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|11920,11930|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|11920,11930|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|11938,11946|false|false|false|||anything
Finding|Functional Concept|Discharge Instructions|11975,11982|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|11975,11982|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|11975,11982|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|11975,11982|false|false|false|C0199168|Medical service|medical
Attribute|Clinical Attribute|Discharge Instructions|11975,11990|false|false|false|C0551625||medical records
Finding|Intellectual Product|Discharge Instructions|11975,11990|false|false|false|C0025102;C1554096|HL7 Committee ID In RIM - Medical records;Medical Records|medical records
Event|Event|Discharge Instructions|11983,11990|false|false|false|||records
Finding|Idea or Concept|Discharge Instructions|11983,11990|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|Discharge Instructions|11983,11990|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|Discharge Instructions|12002,12009|false|false|false|||records
Finding|Idea or Concept|Discharge Instructions|12002,12009|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|Discharge Instructions|12002,12009|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|Discharge Instructions|12021,12036|false|false|false|||hospitalization
Procedure|Health Care Activity|Discharge Instructions|12021,12036|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|Discharge Instructions|12037,12041|false|false|false|||sent
Event|Event|Discharge Instructions|12050,12056|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|12050,12056|false|false|false|C2348314|Doctor - Title|doctor
Finding|Finding|Discharge Instructions|12057,12064|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|12060,12064|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|12060,12064|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|12060,12064|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|12066,12070|false|false|false|||call
Procedure|Health Care Activity|Discharge Instructions|12080,12088|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|12089,12101|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|12089,12101|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|12089,12101|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

