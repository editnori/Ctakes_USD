 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|179,189|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Allergies|179,189|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Allergies|179,189|false|false|false|||omeprazole
Event|Event|Allergies|192,201|false|false|false|||Attending
Finding|Functional Concept|Allergies|192,201|false|false|false|C1999232|Attending (action)|Attending
Disorder|Disease or Syndrome|Chief Complaint|227,236|false|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|Chief Complaint|227,236|false|false|false|||dysphagia
Finding|Classification|Chief Complaint|240,245|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|246,254|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|258,276|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|267,276|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|267,276|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|267,276|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|267,276|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|267,276|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|284,293|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|Chief Complaint|284,293|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|337,344|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|337,344|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|337,344|false|false|false|C0860603|Anxiety symptoms|anxiety
Disorder|Disease or Syndrome|History of Present Illness|366,375|false|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|History of Present Illness|366,375|false|false|false|||dysphagia
Event|Event|History of Present Illness|381,382|false|false|false|||/
Event|Event|History of Present Illness|384,392|false|false|false|||worsened
Finding|Finding|History of Present Illness|384,392|false|false|false|C1457868;C4084902|Got Worse;Worse|worsened
Finding|Intellectual Product|History of Present Illness|384,392|false|false|false|C1457868;C4084902|Got Worse;Worse|worsened
Finding|Idea or Concept|History of Present Illness|394,401|false|false|false|C0376327|International Aspects|foreign
Disorder|Injury or Poisoning|History of Present Illness|394,406|false|false|false|C0016542|Foreign Bodies|foreign body
Finding|Finding|History of Present Illness|394,416|false|false|false|C0423602;C0920171|Foreign body sensation (finding);Foreign body sensation in eyes|foreign body sensation
Anatomy|Anatomical Structure|History of Present Illness|402,406|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|402,406|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|History of Present Illness|402,406|false|false|false|C1551342|Document Body|body
Event|Event|History of Present Illness|407,416|false|false|false|||sensation
Finding|Finding|History of Present Illness|407,416|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|407,416|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|407,416|false|false|false|C2229507|sensory exam|sensation
Event|Event|History of Present Illness|424,433|false|false|false|||describes
Event|Event|History of Present Illness|434,441|false|false|false|||feeling
Drug|Food|History of Present Illness|452,456|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|452,456|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|452,456|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|History of Present Illness|452,456|false|false|false|||food
Event|Event|History of Present Illness|457,461|false|false|false|||gets
Anatomy|Body Location or Region|History of Present Illness|475,479|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|475,479|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|475,479|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|History of Present Illness|490,494|false|false|false|||eats
Drug|Food|History of Present Illness|524,528|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|History of Present Illness|524,528|false|false|false|||diet
Finding|Functional Concept|History of Present Illness|524,528|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|History of Present Illness|524,528|false|false|false|C0012159|Diet therapy|diet
Event|Event|History of Present Illness|532,539|false|false|false|||address
Event|Event|History of Present Illness|545,549|false|false|false|||over
Drug|Food|History of Present Illness|582,586|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|582,586|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|582,586|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Event|Event|History of Present Illness|582,586|false|false|false|||food
Event|Event|History of Present Illness|587,592|false|false|false|||stuck
Anatomy|Body Location or Region|History of Present Illness|600,606|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|600,606|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|History of Present Illness|600,606|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|History of Present Illness|600,606|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|History of Present Illness|600,606|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|History of Present Illness|620,625|false|false|false|||feels
Event|Event|History of Present Illness|647,653|true|false|false|||breath
Finding|Body Substance|History of Present Illness|647,653|true|false|false|C0225386|Breath|breath
Event|Event|History of Present Illness|663,669|true|false|false|||denies
Event|Event|History of Present Illness|670,677|true|false|false|||trouble
Event|Event|History of Present Illness|679,688|true|false|false|||breathing
Finding|Finding|History of Present Illness|702,706|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|702,706|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|702,706|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|730,737|true|false|false|||history
Finding|Conceptual Entity|History of Present Illness|730,737|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|730,737|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|730,737|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|730,740|true|true|false|C0262926|Medical History|history of
Drug|Food|History of Present Illness|742,746|true|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Immunologic Factor|History of Present Illness|742,746|true|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Drug|Pharmacologic Substance|History of Present Illness|742,746|true|false|false|C0016452;C3540798|Food;Food allergenic extracts|food
Disorder|Disease or Syndrome|History of Present Illness|742,756|true|false|false|C0016470|Food Allergy|food allergies
Attribute|Clinical Attribute|History of Present Illness|747,756|true|false|false|C1717415||allergies
Event|Event|History of Present Illness|747,756|true|false|false|||allergies
Finding|Pathologic Function|History of Present Illness|747,756|true|false|false|C0020517|Hypersensitivity|allergies
Anatomy|Body System|History of Present Illness|760,764|true|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|History of Present Illness|760,764|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|History of Present Illness|760,764|true|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|History of Present Illness|760,764|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|History of Present Illness|760,764|true|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Sign or Symptom|History of Present Illness|760,771|true|false|false|C5779628|Skin rash|skin rashes
Event|Event|History of Present Illness|765,771|false|false|false|||rashes
Finding|Sign or Symptom|History of Present Illness|765,771|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Idea or Concept|History of Present Illness|787,794|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|795,801|false|false|false|||vitals
Event|Event|History of Present Illness|835,842|false|false|false|||Imaging
Finding|Finding|History of Present Illness|835,842|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|835,842|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|843,849|false|false|false|||showed
Event|Event|History of Present Illness|851,854|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|851,854|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|855,861|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|874,883|false|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|History of Present Illness|874,883|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|History of Present Illness|874,883|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|History of Present Illness|874,883|false|false|false|||esophagus
Finding|Finding|History of Present Illness|874,883|false|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|874,883|false|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|History of Present Illness|884,892|false|false|false|||Consults
Procedure|Health Care Activity|History of Present Illness|884,892|false|false|false|C0009818|Consultation|Consults
Event|Event|History of Present Illness|901,910|false|false|false|||consulted
Event|Event|History of Present Illness|926,929|false|false|false|||EGD
Procedure|Diagnostic Procedure|History of Present Illness|926,929|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|History of Present Illness|936,942|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|962,971|false|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|History of Present Illness|962,971|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|History of Present Illness|962,971|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|History of Present Illness|962,971|false|false|false|||esophagus
Finding|Finding|History of Present Illness|962,971|false|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|962,971|false|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|History of Present Illness|974,982|false|false|false|||Biopsies
Procedure|Diagnostic Procedure|History of Present Illness|974,982|false|false|false|C0005558|Biopsy|Biopsies
Event|Event|History of Present Illness|988,993|false|false|false|||taken
Event|Event|History of Present Illness|1011,1019|false|false|false|||endorses
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1020,1027|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|1020,1027|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|1020,1027|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|History of Present Illness|1034,1040|false|false|false|||eating
Event|Event|History of Present Illness|1065,1071|false|false|false|||eating
Event|Event|History of Present Illness|1086,1093|false|false|false|||leaving
Event|Event|History of Present Illness|1098,1106|false|false|false|||hospital
Finding|Idea or Concept|History of Present Illness|1098,1106|false|false|false|C1547192|Organization unit type - Hospital|hospital
Disorder|Disease or Syndrome|Past Medical History|1136,1140|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Past Medical History|1136,1140|false|false|false|||GERD
Disorder|Disease or Syndrome|Past Medical History|1146,1166|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|Past Medical History|1146,1166|false|false|false|||Hypercholesterolemia
Finding|Finding|Past Medical History|1146,1166|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1172,1178|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|Past Medical History|1172,1178|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Finding|Sign or Symptom|Past Medical History|1172,1178|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|Past Medical History|1172,1178|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1172,1178|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Disease or Syndrome|Past Medical History|1172,1185|false|false|false|C0392525;C5779632|NEPHROLITHIASIS, CALCIUM OXALATE, 1;Nephrolithiasis|Kidney stones
Finding|Body Substance|Past Medical History|1172,1185|false|false|false|C0022650|Kidney Calculi|Kidney stones
Event|Event|Past Medical History|1179,1185|false|false|false|||stones
Finding|Body Substance|Past Medical History|1179,1185|false|false|false|C0006736|Calculi|stones
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1191,1203|false|false|false|C0026264|Mitral Valve|Mitral valve
Disorder|Disease or Syndrome|Past Medical History|1191,1212|false|false|false|C0026267|Mitral Valve Prolapse Syndrome|Mitral valve prolapse
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1198,1203|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|Past Medical History|1204,1212|false|false|false|C0033377|Ptosis|prolapse
Event|Event|Past Medical History|1204,1212|false|false|false|||prolapse
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1218,1225|false|false|false|C0042149|Uterus|Uterine
Disorder|Neoplastic Process|Past Medical History|1218,1234|false|false|false|C0042133|Uterine Fibroids|Uterine fibroids
Disorder|Neoplastic Process|Past Medical History|1226,1234|false|false|false|C0023267;C0042133|Fibroid Tumor;Uterine Fibroids|fibroids
Event|Event|Past Medical History|1226,1234|false|false|false|||fibroids
Disorder|Disease or Syndrome|Past Medical History|1240,1252|false|false|false|C0029456|Osteoporosis|Osteoporosis
Event|Event|Past Medical History|1240,1252|false|false|false|||Osteoporosis
Finding|Finding|Past Medical History|1240,1252|false|false|false|C2911643|Encounter due to family history of osteoporosis|Osteoporosis
Disorder|Disease or Syndrome|Past Medical History|1258,1266|false|false|false|C0149931|Migraine Disorders|Migraine
Disorder|Disease or Syndrome|Past Medical History|1258,1276|false|false|false|C0149931|Migraine Disorders|Migraine headaches
Event|Event|Past Medical History|1267,1276|false|false|false|||headaches
Finding|Sign or Symptom|Past Medical History|1267,1276|false|false|false|C0018681|Headache|headaches
Disorder|Disease or Syndrome|Family Medical History|1318,1321|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|1318,1321|false|false|false|||HTN
Event|Event|Family Medical History|1324,1330|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|1324,1330|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|1324,1330|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Disorder|Mental or Behavioral Dysfunction|Family Medical History|1335,1343|false|false|false|C0011265;C0497327|Dementia;Presenile dementia|Dementia
Event|Event|Family Medical History|1335,1343|false|false|false|||Dementia
Event|Event|Family Medical History|1346,1352|false|false|false|||father
Finding|Conceptual Entity|Family Medical History|1346,1352|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|1346,1352|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Procedure|Health Care Activity|General Exam|1392,1401|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Body Substance|General Exam|1402,1411|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|1402,1411|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|1402,1411|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|1402,1411|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|1412,1416|false|false|false|||EXAM
Finding|Functional Concept|General Exam|1412,1416|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|1412,1416|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|1471,1474|false|false|false|||GEN
Finding|Classification|General Exam|1471,1474|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|1471,1474|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Mental or Behavioral Dysfunction|General Exam|1481,1488|true|false|false|C0003467|Anxiety|anxious
Event|Event|General Exam|1481,1488|true|false|false|||anxious
Event|Event|General Exam|1496,1501|true|false|false|||lying
Disorder|Disease or Syndrome|General Exam|1505,1508|true|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|1505,1508|true|false|false|C2346952|Bachelor of Education|bed
Finding|Intellectual Product|General Exam|1513,1518|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|1519,1527|true|false|false|||distress
Finding|Finding|General Exam|1519,1527|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|1519,1527|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|1530,1535|true|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|1547,1556|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|1557,1564|false|false|false|||sclerae
Event|Event|General Exam|1566,1570|false|false|false|||NCAT
Event|Event|General Exam|1572,1577|false|false|false|||PERRL
Finding|Finding|General Exam|1572,1577|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|1579,1583|false|false|false|||EOMI
Anatomy|Body Location or Region|General Exam|1586,1590|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|1586,1590|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|1586,1590|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|1592,1598|true|false|false|||Supple
Finding|Functional Concept|General Exam|1592,1598|true|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|1607,1610|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|1607,1610|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|1607,1610|true|false|false|||LAD
Finding|Gene or Genome|General Exam|1607,1610|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|1615,1618|true|false|false|||JVD
Finding|Finding|General Exam|1615,1618|true|false|false|C0425687|Jugular venous engorgement|JVD
Event|Event|General Exam|1621,1625|true|false|false|||PULM
Procedure|Health Care Activity|General Exam|1621,1625|true|false|false|C1315068|Pulmonary ventilator management|PULM
Anatomy|Body Part, Organ, or Organ Component|General Exam|1642,1645|true|false|false|C0018787|Heart|COR
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1642,1645|true|false|false|C0056331|cordycepin|COR
Drug|Pharmacologic Substance|General Exam|1642,1645|true|false|false|C0056331|cordycepin|COR
Anatomy|Body Location or Region|General Exam|1671,1674|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|1671,1674|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|1671,1674|true|false|false|||ABD
Disorder|Disease or Syndrome|General Exam|1676,1680|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|1676,1680|false|false|false|||Soft
Event|Event|General Exam|1717,1720|true|false|false|||HSM
Finding|Gene or Genome|General Exam|1717,1720|true|false|false|C1537594|LRRC4B gene|HSM
Event|Event|General Exam|1731,1735|true|false|false|||Warm
Finding|Finding|General Exam|1731,1735|true|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1731,1735|true|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1737,1741|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1742,1750|true|false|false|||perfused
Attribute|Clinical Attribute|General Exam|1759,1764|true|false|false|C1717255||edema
Event|Event|General Exam|1759,1764|true|false|false|||edema
Finding|Pathologic Function|General Exam|1759,1764|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|1792,1798|false|false|false|||intact
Finding|Finding|General Exam|1792,1798|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|General Exam|1800,1805|false|false|false|C1513492|motor movement|motor
Finding|Finding|General Exam|1800,1814|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|General Exam|1800,1814|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|General Exam|1806,1814|false|false|false|||function
Finding|Finding|General Exam|1806,1814|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|1806,1814|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|1806,1814|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|1806,1814|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|General Exam|1832,1841|false|false|false|||sensation
Finding|Finding|General Exam|1832,1841|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|1832,1841|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|1832,1841|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|1850,1856|false|false|false|||intact
Finding|Finding|General Exam|1850,1856|false|false|false|C1554187|Gender Status - Intact|intact
Procedure|Health Care Activity|General Exam|1894,1903|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|1904,1908|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|1904,1908|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|1936,1941|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|1936,1941|false|false|false|||BLOOD
Finding|Body Substance|General Exam|1936,1941|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|1942,1945|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|1950,1953|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|1950,1953|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|1950,1953|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|1959,1962|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|1959,1962|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|1959,1962|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|1959,1962|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|1968,1971|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|1968,1971|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|1977,1980|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|1977,1980|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|1977,1980|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|1977,1980|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|1977,1980|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|1985,1988|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|1985,1988|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|1985,1988|false|false|false|||MCH
Finding|Gene or Genome|General Exam|1985,1988|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|1985,1988|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|1985,1988|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|1994,1998|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|1994,1998|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|2024,2027|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|2044,2049|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2044,2049|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2044,2049|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2054,2057|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|2054,2057|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|2054,2057|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|2079,2084|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2079,2084|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2079,2084|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|2079,2092|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|2079,2092|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|2079,2092|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|2085,2092|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|2085,2092|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|2085,2092|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|2085,2092|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|2085,2092|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|2085,2092|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|2116,2117|false|false|false|||-
Drug|Inorganic Chemical|General Exam|2135,2139|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|2135,2139|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|2135,2139|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|2164,2169|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2164,2169|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2164,2169|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|2170,2173|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|2170,2173|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|2170,2173|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|2170,2173|false|false|false|||ALT
Finding|Gene or Genome|General Exam|2170,2173|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|2170,2173|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|2170,2173|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|2170,2173|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|2177,2180|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|2177,2180|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2177,2180|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|2177,2180|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|2177,2180|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|2177,2180|false|false|false|||AST
Finding|Gene or Genome|General Exam|2177,2180|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|2187,2190|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|General Exam|2187,2190|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|General Exam|2187,2190|false|false|false|||LDH
Finding|Finding|General Exam|2187,2190|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|General Exam|2187,2190|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|General Exam|2196,2203|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|2196,2203|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|2232,2237|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|2232,2237|false|false|false|||BLOOD
Finding|Body Substance|General Exam|2232,2237|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|2232,2245|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|2238,2245|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|2238,2245|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|2238,2245|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|2238,2245|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|2238,2245|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|2238,2245|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|2238,2245|false|false|false|C0201838|Albumin measurement|Albumin
Event|Event|General Exam|2264,2271|false|false|false|||IMAGING
Finding|Finding|General Exam|2264,2271|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|2264,2271|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|2287,2290|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|2287,2290|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Body Part, Organ, or Organ Component|Impression|2324,2333|true|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|Impression|2324,2333|true|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|Impression|2324,2333|true|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|Impression|2324,2333|true|false|false|||esophagus
Finding|Finding|Impression|2324,2333|true|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|Impression|2324,2333|true|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|Impression|2345,2349|true|false|false|||view
Drug|Inorganic Chemical|Impression|2359,2362|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Impression|2359,2362|true|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Impression|2359,2362|true|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Impression|2359,2362|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Impression|2359,2362|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Impression|2359,2362|true|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Substance|Impression|2363,2368|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Impression|2363,2368|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Impression|2369,2374|true|false|false|||level
Finding|Body Substance|Impression|2387,2394|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|2387,2394|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|2387,2394|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|2397,2404|false|false|false|||history
Finding|Conceptual Entity|Impression|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Impression|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Impression|2397,2404|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Phenomenon|Natural Phenomenon or Process|Impression|2409,2421|false|false|false|C0444708|Radiographic|radiographic
Attribute|Clinical Attribute|Impression|2422,2432|false|false|false|C0550215||appearance
Event|Event|Impression|2422,2432|false|false|false|||appearance
Procedure|Health Care Activity|Impression|2422,2432|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Drug|Element, Ion, or Isotope|Impression|2434,2440|false|false|false|C0004749|barium|barium
Event|Event|Impression|2434,2440|false|false|false|||barium
Event|Event|Impression|2442,2449|false|false|false|||swallow
Finding|Functional Concept|Impression|2442,2449|false|false|false|C1706486;C4521686|Swallow (administration method);Swallow - dosing instruction imperative|swallow
Event|Event|Impression|2453,2462|false|false|false|||indicated
Anatomy|Body Location or Region|Impression|2493,2497|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Impression|2493,2497|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Impression|2493,2497|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Procedure|Diagnostic Procedure|Impression|2493,2503|false|false|false|C0202757;C1963529|Neck X-ray;Radiographic procedure on neck|NECK X-ray
Event|Event|Impression|2498,2503|false|false|false|||X-ray
Finding|Functional Concept|Impression|2498,2503|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-ray
Finding|Intellectual Product|Impression|2498,2503|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|X-ray
Phenomenon|Natural Phenomenon or Process|Impression|2498,2503|false|false|false|C0043309|Roentgen Rays|X-ray
Procedure|Diagnostic Procedure|Impression|2498,2503|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|X-ray
Event|Event|Impression|2537,2547|true|false|false|||limitation
Finding|Functional Concept|Impression|2537,2547|true|false|false|C0443288;C0449295|Limitation;Restricted|limitation
Procedure|Diagnostic Procedure|Impression|2551,2568|true|false|false|C1306645|Plain x-ray|plain radiography
Event|Event|Impression|2557,2568|true|false|false|||radiography
Finding|Functional Concept|Impression|2557,2568|true|false|false|C0034571|roentgenographic|radiography
Procedure|Diagnostic Procedure|Impression|2557,2568|true|false|false|C0043299;C1962945;C4721829|Diagnostic radiologic examination;Radiographic Examination;Radiographic imaging procedure|radiography
Event|Event|Impression|2573,2581|true|false|false|||evidence
Finding|Idea or Concept|Impression|2573,2581|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|2573,2584|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Impression|2599,2603|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Impression|2599,2610|true|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Impression|2599,2610|true|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Disorder|Disease or Syndrome|Impression|2599,2619|true|false|false|C0037580|Soft tissue swelling|soft tissue swelling
Anatomy|Tissue|Impression|2604,2610|true|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Impression|2604,2610|true|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|Impression|2611,2619|true|false|false|||swelling
Finding|Finding|Impression|2611,2619|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Impression|2611,2619|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|Impression|2623,2627|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Impression|2623,2634|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Impression|2623,2634|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Disorder|Anatomical Abnormality|Impression|2623,2639|false|false|false|C0457193|Soft tissue mass|soft tissue mass
Anatomy|Tissue|Impression|2628,2634|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Impression|2628,2634|false|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|Impression|2635,2639|false|false|false|||mass
Finding|Finding|Impression|2635,2639|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Impression|2635,2639|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Impression|2635,2639|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Anatomy|Body Location or Region|Impression|2648,2652|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Impression|2648,2652|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Impression|2648,2652|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|Impression|2658,2661|false|false|false|||EGD
Procedure|Diagnostic Procedure|Impression|2658,2661|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Impression|2668,2678|false|false|false|||Impression
Finding|Intellectual Product|Impression|2668,2678|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Finding|Mental Process|Impression|2668,2678|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|Impression
Disorder|Acquired Abnormality|Impression|2680,2693|false|false|false|C3489393|Hiatal Hernia|Hiatal hernia
Disorder|Anatomical Abnormality|Impression|2687,2693|false|false|false|C0019270|Hernia|hernia
Event|Event|Impression|2687,2693|false|false|false|||hernia
Disorder|Disease or Syndrome|Impression|2694,2706|false|false|false|C0002959|Angiectasis|Angioectasia
Event|Event|Impression|2694,2706|false|false|false|||Angioectasia
Anatomy|Body Part, Organ, or Organ Component|Impression|2714,2721|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Impression|2714,2721|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Impression|2714,2721|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Impression|2714,2721|false|false|false|||stomach
Finding|Finding|Impression|2714,2721|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Impression|2714,2721|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Disease or Syndrome|Impression|2722,2734|false|false|false|C0002959|Angiectasis|Angioectasia
Event|Event|Impression|2722,2734|false|false|false|||Angioectasia
Anatomy|Body Part, Organ, or Organ Component|Impression|2742,2750|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|Impression|2742,2750|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Event|Event|Impression|2753,2759|false|false|false|||biopsy
Finding|Finding|Impression|2753,2759|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Impression|2753,2759|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Impression|2753,2759|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Impression|2753,2759|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Impression|2761,2767|false|false|false|||biopsy
Finding|Finding|Impression|2761,2767|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Impression|2761,2767|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Impression|2761,2767|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Impression|2761,2767|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Impression|2786,2789|false|false|false|||EGD
Procedure|Diagnostic Procedure|Impression|2786,2789|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Impression|2799,2803|false|false|false|||part
Finding|Idea or Concept|Impression|2799,2803|false|false|false|C1552020|Role Class - part|part
Anatomy|Body Part, Organ, or Organ Component|Impression|2811,2819|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|Impression|2811,2819|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Event|Event|Impression|2822,2837|false|false|false|||Recommendations
Finding|Idea or Concept|Impression|2822,2837|false|false|false|C0034866|Recommendation|Recommendations
Event|Event|Impression|2861,2866|true|false|false|||cause
Finding|Conceptual Entity|Impression|2861,2866|true|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Impression|2861,2866|true|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Body Substance|Impression|2875,2882|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Impression|2875,2882|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Impression|2875,2882|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Impression|2886,2894|false|false|false|||symptoms
Finding|Functional Concept|Impression|2886,2894|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Impression|2886,2894|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Impression|2897,2903|true|false|false|||follow
Finding|Functional Concept|Impression|2897,2903|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Impression|2897,2903|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Impression|2897,2906|true|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Impression|2897,2906|true|false|false|C1522577|follow-up|follow-up
Event|Event|Impression|2907,2913|true|false|false|||biopsy
Finding|Finding|Impression|2907,2913|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|Impression|2907,2913|true|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|Impression|2907,2913|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|Impression|2907,2913|true|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Event|Event|Impression|2914,2921|true|false|false|||results
Event|Event|Impression|2925,2929|false|false|false|||rule
Finding|Functional Concept|Impression|2934,2946|true|false|false|C0333930|eosinophilic|eosinophilic
Disorder|Disease or Syndrome|Impression|2934,2958|true|false|false|C0341106|Eosinophilic esophagitis|eosinophilic esophagitis
Finding|Finding|Impression|2934,2958|true|false|false|C4703646|Eosinophilic infiltration of the esophagus|eosinophilic esophagitis
Disorder|Disease or Syndrome|Impression|2947,2958|true|false|false|C0014868|Esophagitis|esophagitis
Event|Event|Impression|2947,2958|true|false|false|||esophagitis
Event|Event|Impression|2961,2967|true|false|false|||follow
Finding|Functional Concept|Impression|2961,2967|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Impression|2961,2967|true|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Impression|2961,2970|true|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Impression|2961,2970|true|false|false|C1522577|follow-up|follow-up
Event|Event|Impression|2968,2970|false|false|false|||up
Event|Event|Impression|2987,2995|false|false|false|||biopsies
Procedure|Diagnostic Procedure|Impression|2987,2995|false|false|false|C0005558|Biopsy|biopsies
Event|Event|Impression|3001,3013|false|false|false|||eosinophilic
Finding|Functional Concept|Impression|3001,3013|false|false|false|C0333930|eosinophilic|eosinophilic
Disorder|Disease or Syndrome|Impression|3015,3026|false|false|false|C0014868|Esophagitis|esophagitis
Event|Event|Impression|3015,3026|false|false|false|||esophagitis
Event|Event|Hospital Course|3076,3083|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|3076,3083|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3076,3083|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|3076,3083|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|3076,3086|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|3087,3091|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Hospital Course|3087,3091|false|false|false|||GERD
Event|Event|Hospital Course|3096,3104|false|false|false|||presents
Event|Event|Hospital Course|3120,3129|false|false|false|||worsening
Finding|Idea or Concept|Hospital Course|3120,3129|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|Hospital Course|3133,3142|false|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|Hospital Course|3133,3142|false|false|false|||dysphagia
Finding|Idea or Concept|Hospital Course|3147,3154|false|false|false|C0376327|International Aspects|foreign
Disorder|Injury or Poisoning|Hospital Course|3147,3159|false|false|false|C0016542|Foreign Bodies|foreign body
Finding|Finding|Hospital Course|3147,3169|false|false|false|C0423602;C0920171|Foreign body sensation (finding);Foreign body sensation in eyes|foreign body sensation
Anatomy|Anatomical Structure|Hospital Course|3155,3159|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3155,3159|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Hospital Course|3155,3159|false|false|false|C1551342|Document Body|body
Event|Event|Hospital Course|3160,3169|false|false|false|||sensation
Finding|Finding|Hospital Course|3160,3169|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Hospital Course|3160,3169|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Hospital Course|3160,3169|false|false|false|C2229507|sensory exam|sensation
Event|Event|Hospital Course|3181,3189|false|false|false|||worsened
Event|Event|Hospital Course|3213,3219|false|false|false|||placed
Event|Event|Hospital Course|3233,3239|false|false|false|||pureed
Drug|Food|Hospital Course|3241,3245|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|3241,3245|false|false|false|||diet
Finding|Functional Concept|Hospital Course|3241,3245|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|3241,3245|false|false|false|C0012159|Diet therapy|diet
Event|Event|Hospital Course|3282,3285|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|3282,3285|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|3292,3298|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3312,3321|false|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|Hospital Course|3312,3321|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|Hospital Course|3312,3321|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|Hospital Course|3312,3321|false|false|false|||esophagus
Finding|Finding|Hospital Course|3312,3321|false|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3312,3321|false|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|Hospital Course|3340,3346|false|false|false|||normal
Event|Event|Hospital Course|3356,3365|false|false|false|||evaluated
Finding|Intellectual Product|Hospital Course|3370,3386|false|false|false|C4050121|Gastrointestinal studies and measurements|Gastroenterology
Event|Event|Hospital Course|3410,3419|false|false|false|||endoscopy
Procedure|Diagnostic Procedure|Hospital Course|3410,3419|false|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|Hospital Course|3434,3440|false|false|false|||showed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3460,3469|false|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|Hospital Course|3460,3469|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|Hospital Course|3460,3469|false|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|Hospital Course|3460,3469|false|false|false|||esophagus
Finding|Finding|Hospital Course|3460,3469|false|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3460,3469|false|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|Hospital Course|3471,3479|false|false|false|||Biopsies
Procedure|Diagnostic Procedure|Hospital Course|3471,3479|false|false|false|C0005558|Biopsy|Biopsies
Event|Event|Hospital Course|3485,3490|false|false|false|||taken
Finding|Idea or Concept|Hospital Course|3494,3506|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|3507,3513|false|false|false|||ISSUES
Event|Event|Hospital Course|3520,3528|false|false|false|||biopsies
Procedure|Diagnostic Procedure|Hospital Course|3520,3528|false|false|false|C0005558|Biopsy|biopsies
Event|Event|Hospital Course|3534,3537|false|false|false|||EGD
Procedure|Diagnostic Procedure|Hospital Course|3534,3537|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|Hospital Course|3542,3549|false|false|false|||results
Finding|Functional Concept|Hospital Course|3555,3567|false|false|false|C0333930|eosinophilic|eosinophilic
Disorder|Disease or Syndrome|Hospital Course|3555,3579|false|false|false|C0341106|Eosinophilic esophagitis|eosinophilic esophagitis
Finding|Finding|Hospital Course|3555,3579|false|false|false|C4703646|Eosinophilic infiltration of the esophagus|eosinophilic esophagitis
Disorder|Disease or Syndrome|Hospital Course|3568,3579|false|false|false|C0014868|Esophagitis|esophagitis
Event|Event|Hospital Course|3568,3579|false|false|false|||esophagitis
Event|Event|Hospital Course|3581,3587|false|false|false|||follow
Event|Event|Hospital Course|3614,3624|false|false|false|||management
Event|Occupational Activity|Hospital Course|3614,3624|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|3614,3624|false|false|false|C0376636|Disease Management|management
Drug|Element, Ion, or Isotope|Hospital Course|3644,3650|false|false|false|C0004749|barium|barium
Event|Event|Hospital Course|3644,3650|false|false|false|||barium
Procedure|Diagnostic Procedure|Hospital Course|3644,3658|false|false|false|C0203065|Barium swallow|barium swallow
Event|Event|Hospital Course|3651,3658|false|false|false|||swallow
Finding|Functional Concept|Hospital Course|3651,3658|false|false|false|C1706486;C4521686|Swallow (administration method);Swallow - dosing instruction imperative|swallow
Event|Event|Hospital Course|3665,3675|false|false|false|||outpatient
Finding|Classification|Hospital Course|3665,3675|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|3665,3675|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|3689,3695|false|false|false|||workup
Disorder|Disease or Syndrome|Hospital Course|3703,3712|false|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|Hospital Course|3703,3712|false|false|false|||dysphagia
Anatomy|Body Location or Region|Hospital Course|3723,3726|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3723,3726|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|Hospital Course|3723,3726|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|Hospital Course|3723,3726|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Event|Event|Hospital Course|3730,3737|false|false|false|||planned
Event|Event|Hospital Course|3739,3743|false|false|false|||Code
Event|Occupational Activity|Hospital Course|3739,3743|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|3739,3743|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|Hospital Course|3751,3759|false|false|false|||presumed
Attribute|Clinical Attribute|Hospital Course|3764,3775|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3764,3775|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|3764,3775|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|3764,3775|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|3764,3788|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|3779,3788|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|3779,3788|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|3807,3817|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|3807,3817|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|3807,3822|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|3818,3822|false|false|false|||list
Finding|Intellectual Product|Hospital Course|3818,3822|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|3826,3834|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|3839,3847|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|3839,3847|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|3839,3847|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|3839,3847|false|false|false|||complete
Finding|Functional Concept|Hospital Course|3839,3847|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|3839,3847|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|3852,3862|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|3852,3862|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3872,3875|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3872,3875|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3872,3875|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|3872,3875|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|3872,3875|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|3880,3889|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3880,3889|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3880,3889|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3880,3889|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3880,3889|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3880,3901|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|3890,3901|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3890,3901|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|3890,3901|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|3890,3901|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|3907,3917|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|3907,3917|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3927,3930|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3927,3930|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3927,3930|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|3927,3930|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|3927,3930|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|3936,3945|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3936,3945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3936,3945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3936,3945|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3936,3945|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|3936,3957|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|3936,3957|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|3946,3957|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|3946,3957|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|3946,3957|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|3959,3963|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|3959,3963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|3959,3963|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|3959,3963|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|3966,3975|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3966,3975|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3966,3975|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3966,3975|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3966,3975|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3966,3985|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|3976,3985|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|3976,3985|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|3976,3985|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|3976,3985|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|3976,3985|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|4007,4016|false|false|false|C0011168|Deglutition Disorders|dysphagia
Event|Event|Principle Diagnosis|4007,4016|false|false|false|||dysphagia
Finding|Idea or Concept|Principle Diagnosis|4021,4028|false|false|false|C0376327|International Aspects|foreign
Disorder|Injury or Poisoning|Principle Diagnosis|4021,4033|false|false|false|C0016542|Foreign Bodies|foreign body
Finding|Finding|Principle Diagnosis|4021,4043|false|false|false|C0423602;C0920171|Foreign body sensation (finding);Foreign body sensation in eyes|foreign body sensation
Anatomy|Anatomical Structure|Principle Diagnosis|4029,4033|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Principle Diagnosis|4029,4033|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Principle Diagnosis|4029,4033|false|false|false|C1551342|Document Body|body
Event|Event|Principle Diagnosis|4034,4043|false|false|false|||sensation
Finding|Finding|Principle Diagnosis|4034,4043|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Principle Diagnosis|4034,4043|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Principle Diagnosis|4034,4043|false|false|false|C2229507|sensory exam|sensation
Disorder|Neoplastic Process|Principle Diagnosis|4045,4054|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Event|Event|Principle Diagnosis|4045,4054|false|false|false|||SECONDARY
Finding|Functional Concept|Principle Diagnosis|4045,4054|false|false|false|C1522484|metastatic qualifier|SECONDARY
Attribute|Clinical Attribute|Principle Diagnosis|4045,4064|false|false|false|C4255018||SECONDARY DIAGNOSIS
Finding|Finding|Principle Diagnosis|4045,4064|false|false|false|C0332138|Secondary diagnosis|SECONDARY DIAGNOSIS
Attribute|Clinical Attribute|Principle Diagnosis|4055,4064|false|false|false|C0945731||DIAGNOSIS
Finding|Classification|Principle Diagnosis|4055,4064|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Finding|Functional Concept|Principle Diagnosis|4055,4064|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|DIAGNOSIS
Procedure|Diagnostic Procedure|Principle Diagnosis|4055,4064|false|false|false|C0011900|Diagnosis|DIAGNOSIS
Disorder|Disease or Syndrome|Principle Diagnosis|4067,4071|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|Principle Diagnosis|4067,4071|false|false|false|||GERD
Finding|Mental Process|Discharge Condition|4097,4103|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|4097,4110|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|4097,4110|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|4104,4110|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|4104,4110|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|4112,4117|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|4112,4117|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|4122,4130|false|false|false|||coherent
Finding|Finding|Discharge Condition|4122,4130|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|4132,4137|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|4132,4154|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|4132,4154|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|4141,4154|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|4141,4154|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|4141,4154|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|4156,4161|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|4156,4161|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|4156,4161|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|4156,4161|false|false|false|||Alert
Finding|Finding|Discharge Condition|4156,4161|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|4156,4161|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|4156,4161|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|4166,4177|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|4166,4177|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|4179,4187|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|4179,4187|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|4179,4187|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|4188,4194|false|false|false|C5889824||Status
Event|Event|Discharge Condition|4188,4194|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|4188,4194|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|4196,4206|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|4196,4206|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|4196,4206|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|4196,4206|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|4196,4206|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|4209,4220|false|false|false|||Independent
Finding|Finding|Discharge Condition|4209,4220|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|4209,4220|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|4249,4253|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|4273,4285|false|false|false|||hospitalized
Event|Event|Discharge Instructions|4299,4303|false|false|false|||came
Event|Event|Discharge Instructions|4314,4324|false|false|false|||difficulty
Finding|Finding|Discharge Instructions|4314,4324|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Discharge Instructions|4325,4335|false|false|false|||swallowing
Event|Event|Discharge Instructions|4348,4357|true|false|false|||endoscopy
Procedure|Diagnostic Procedure|Discharge Instructions|4348,4357|true|false|false|C0014245;C0079278|Endoscopy (procedure);Endoscopy, Gastrointestinal|endoscopy
Event|Event|Discharge Instructions|4362,4366|true|false|false|||look
Disorder|Congenital Abnormality|Discharge Instructions|4375,4388|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Discharge Instructions|4375,4388|true|false|false|||abnormalities
Finding|Functional Concept|Discharge Instructions|4375,4388|true|false|false|C0000769|teratologic|abnormalities
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4396,4405|true|false|false|C0014876;C4266613|Chest>Esophagus;Esophagus|esophagus
Disorder|Disease or Syndrome|Discharge Instructions|4396,4405|true|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Disorder|Neoplastic Process|Discharge Instructions|4396,4405|true|false|false|C0014852;C0153942;C0154059|Benign neoplasm of esophagus;Carcinoma in situ of esophagus;Esophageal Diseases|esophagus
Event|Event|Discharge Instructions|4396,4405|true|false|false|||esophagus
Finding|Finding|Discharge Instructions|4396,4405|true|false|false|C0812418|Esophagus problem|esophagus
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4396,4405|true|false|false|C0872395|Procedures on the esophagus|esophagus
Event|Event|Discharge Instructions|4429,4435|false|false|false|||normal
Event|Event|Discharge Instructions|4447,4455|false|false|false|||biopsies
Procedure|Diagnostic Procedure|Discharge Instructions|4447,4455|false|false|false|C0005558|Biopsy|biopsies
Event|Event|Discharge Instructions|4473,4479|false|false|false|||called
Event|Event|Discharge Instructions|4490,4497|false|false|false|||results
Anatomy|Body Location or Region|Discharge Instructions|4517,4521|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Discharge Instructions|4517,4521|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|4517,4521|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|4517,4521|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|4517,4521|false|false|false|C0022885|Laboratory Procedures|test
Event|Event|Discharge Instructions|4522,4528|false|false|false|||called
Drug|Element, Ion, or Isotope|Discharge Instructions|4531,4537|false|false|false|C0004749|barium|barium
Procedure|Diagnostic Procedure|Discharge Instructions|4531,4545|false|false|false|C0203065|Barium swallow|barium swallow
Event|Event|Discharge Instructions|4538,4545|false|false|false|||swallow
Finding|Functional Concept|Discharge Instructions|4538,4545|false|false|false|C1706486;C4521686|Swallow (administration method);Swallow - dosing instruction imperative|swallow
Event|Event|Discharge Instructions|4553,4563|false|false|false|||outpatient
Finding|Classification|Discharge Instructions|4553,4563|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|4553,4563|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Discharge Instructions|4586,4590|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|4586,4590|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|4586,4590|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Procedure|Health Care Activity|Discharge Instructions|4610,4618|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|4619,4631|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|4619,4631|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|4619,4631|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

