CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|Iodine, Homeopathic preparation|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodine
null|iodine|Drug|false|false||Iodinenull|Iodides|Drug|false|false||Iodidenull|Containing (qualifier value)|Finding|false|false||Containingnull|Contain (action)|Event|false|false||Containingnull|Hallucinogens|Drug|false|false||hallucinogens
null|Hallucinogens|Drug|false|false||hallucinogensnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Pain of left hip joint|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|Left hip painnull|Left hip region structure|Anatomy|false|false|C2598155;C1292890;C0019559;C4551516;C2141922;C1430701;C0529134;C1505163;C1654726;C1552822;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725;C1549543;C0030193;C1716793|Left hipnull|Table Cell Horizontal Align - left|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Hip joint pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip pain
null|Hip pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip painnull|null|Attribute|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip painnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|hipnull|RPL29 wt Allele|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0524471;C0022122;C0228391;C0019552;C4299095|hipnull|Lower extremity>Hip|Anatomy|false|false|C0019559;C4551516;C1549543;C0030193;C1292890;C1430701;C0529134;C1505163;C1654726;C1552822;C1716793;C2141922;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Hip structure|Anatomy|false|false|C0019559;C4551516;C1549543;C0030193;C1292890;C1430701;C0529134;C1505163;C1654726;C1552822;C1716793;C2141922;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Structure of habenulopeduncular tract|Anatomy|false|false|C0019559;C4551516;C1549543;C0030193;C1292890;C1430701;C0529134;C1505163;C1654726;C1552822;C1716793;C2141922;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Bone structure of ischium|Anatomy|false|false|C0019559;C4551516;C1549543;C0030193;C1292890;C1430701;C0529134;C1505163;C1654726;C1552822;C1716793;C2141922;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hipnull|Administration Method - Pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|pain
null|Pain|Finding|false|false|C0022122;C0228391;C0019552;C4299095;C0524471|painnull|null|Attribute|false|false|C0524471|painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Indication of (contextual qualifier)|Finding|false|false||REASON FORnull|Indication of (contextual qualifier)|Finding|false|false||REASONnull|Consultation|Procedure|false|false||CONSULTnull|Femoral Fractures|Disorder|false|false|C4299098;C0015811|Femur fracturenull|Lower extremity>Femur|Anatomy|false|false|C0015802;C0016658|Femur
null|Femur|Anatomy|false|false|C0015802;C0016658|Femurnull|Fracture|Disorder|false|false|C4299098;C0015811|fracturenull|Proline dehydrogenase deficiency|Disorder|false|false||HPInull|History of present illness (finding)|Finding|false|false||HPI
null|allene oxide synthase activity|Finding|false|false||HPInull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Fracture|Disorder|false|false||fracturenull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Morning|Time|false|false||morningnull|Dog antigen|Drug|false|false||dognull|allergy testing dog|Procedure|false|false||dognull|Dog family|Entity|false|false||dog
null|Canis familiaris|Entity|false|false||dognull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Movement|Finding|false|false||movementnull|Problems with head|Disorder|false|false|C0018670;C0152336|Headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|Headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076|Head
null|Head|Anatomy|false|false|C0876917;C0362076|Headnull|Head Device|Device|false|false||Headnull|Strikes, Employee|Event|false|false||strikenull|Location|Modifier|false|false||LOCnull|Anticoagulants|Drug|true|false||blood thinnersnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Thinners|Drug|false|false||thinnersnull|Numbness|Finding|true|false|C0278454;C0015385|numbness
null|Hypesthesia|Finding|true|false|C0278454;C0015385|numbnessnull|Weakness|Finding|true|false|C0278454;C0015385|weakness
null|Asthenia|Finding|true|false|C0278454;C0015385|weaknessnull|All extremities|Anatomy|false|false|C3714552;C0004093;C0028643;C0020580|extremities
null|Limb structure|Anatomy|false|false|C3714552;C0004093;C0028643;C0020580|extremitiesnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|NEPHROLITHIASIS, CALCIUM OXALATE, 1|Disorder|false|false|C0227665;C0022646|Kidney stones
null|Nephrolithiasis|Disorder|false|false|C0227665;C0022646|Kidney stonesnull|Kidney Calculi|Finding|false|false|C0227665;C0022646|Kidney stonesnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|Kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|Kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|Kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|Kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|Kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0006736;C0022650;C0392525;C5779632;C0812426|Kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0006736;C0022650;C0392525;C5779632;C0812426|Kidneynull|Calculi|Finding|false|false|C0227665;C0022646|stonesnull|stones - unit|LabModifier|false|false||stonesnull|Mitral Valve Prolapse Syndrome|Disorder|false|false|C1186983;C0026264|Mitral valve prolapsenull|Mitral Valve|Anatomy|false|false|C0026267;C0033377|Mitral valvenull|mitral|Modifier|false|false||Mitralnull|Anatomical valve|Anatomy|false|false|C0026267;C0033377|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Ptosis|Disorder|false|false|C1186983;C0026264|prolapsenull|Uterine Fibroids|Disorder|false|false|C0042149|Uterine fibroidsnull|Uterus|Anatomy|false|false|C0023267;C0042133;C0042133|Uterinenull|Uterine Fibroids|Disorder|false|false|C0042149|fibroids
null|Fibroid Tumor|Disorder|false|false|C0042149|fibroidsnull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Migraine Disorders|Disorder|false|false||Migraine headachesnull|Migraine Disorders|Disorder|false|false||Migrainenull|Headache|Finding|false|false||headachesnull|Hypertensive disease|Disorder|false|false||HTNnull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Left lower extremity|Anatomy|false|false|C1552822;C2003888|Left Lower extremitynull|Table Cell Horizontal Align - left|Finding|false|false|C0230416;C0023216;C1548802|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Lower Extremity|Anatomy|false|false|C1552822|Lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888;C1552822|Lowernull|Lower (action)|Event|false|false|C1548802;C0230416|Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Limb structure|Anatomy|false|false||extremitynull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1554187;C1546781;C0444099|Skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1554187;C1546781;C0444099|Skinnull|Gender Status - Intact|Finding|false|false|C1123023;C4520765|intactnull|Intact|Modifier|false|false||intactnull|Deformity|Disorder|true|false||deformity
null|Congenital Abnormality|Disorder|true|false||deformitynull|null|Finding|true|false||deformitynull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Ecchymosis|Finding|true|false||ecchymosis
null|Skin Bruise|Finding|true|false||ecchymosisnull|Erythema|Disorder|false|false||erythemanull|Induration|Finding|false|false||indurationnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Full|Modifier|false|false||Fullnull|Painless|Finding|false|false||painlessnull|Rupture of Membranes|Finding|false|false|C1963703;C0022742;C4299094;C0022745|ROM
null|ROM1 gene|Finding|false|false|C1963703;C0022742;C4299094;C0022745|ROMnull|Range of motion technique (procedure)|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C1419600;C0948106;C0562271;C1562926|knee
null|Knee|Anatomy|false|false|C1419600;C0948106;C0562271;C1562926|knee
null|Lower extremity>Knee|Anatomy|false|false|C1419600;C0948106;C0562271;C1562926|knee
null|Knee joint|Anatomy|false|false|C1419600;C0948106;C0562271;C1562926|kneenull|Lower extremity>Ankle|Anatomy|false|false||ankle
null|Ankle|Anatomy|false|false||ankle
null|Ankle joint structure|Anatomy|false|false||anklenull|Febrile infection related epilepsy syndrome|Disorder|false|false||Firesnull|Fire (physical force)|Phenomenon|false|false||Firesnull|fire disaster|Event|false|false||Firesnull|Spatial Distribution|Modifier|false|false||distributionsnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Accident and Emergency department|Device|false|false||emergency departmentnull|Accident and Emergency department|Entity|false|false||emergency department
null|interventional services emergency department|Entity|false|false||emergency departmentnull|Certification patient type - Emergency|Finding|false|false||emergency
null|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Department - No suggested values defined|Finding|false|false||department
null|Organization Unit Type - Department|Finding|false|false||department
null|Department - Charge type|Finding|false|false||departmentnull|Department|Entity|false|false||departmentnull|Patient location type - Department|Modifier|false|false||department
null|Department - Person location type|Modifier|false|false||departmentnull|Orthopedic Rehabilitation Surgery|Procedure|false|false||orthopedic surgery
null|Orthopedic Surgical Procedures|Procedure|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Team|Subject|false|false||teamnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Valgus deformity|Disorder|false|false|C0015815|valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Femoral Neck Fractures|Disorder|false|false|C0015811;C0027530;C3159206;C0015815|femoral neck fracturenull|Structure of neck of femur|Anatomy|false|false|C0262414;C0016658;C0015806;C0042282;C0812434;C0684335|femoral necknull|Femur|Anatomy|false|false|C0015806;C0262414;C0016658;C0812434;C0684335|femoralnull|Fracture of cervical spine|Disorder|false|false|C0015815;C0015811;C0027530;C3159206|neck fracturenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0015811;C0015815|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0015811;C0015815|necknull|dendritic spine neck|Anatomy|false|false|C0016658;C0262414;C0015806;C0812434;C0684335|neck
null|Neck|Anatomy|false|false|C0016658;C0262414;C0015806;C0812434;C0684335|necknull|Fracture|Disorder|false|false|C0027530;C3159206;C0015811;C0015815|fracturenull|Orthopedic Rehabilitation Surgery|Procedure|false|false||orthopedic surgery
null|Orthopedic Surgical Procedures|Procedure|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Reduced|Finding|false|false||reductionnull|Reduction procedure|Procedure|false|false||reduction
null|Surgical reduction|Procedure|false|false||reductionnull|Reduction (chemical)|Phenomenon|false|false||reductionnull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Intramedullary Nailing|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|pinningnull|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP protein, human|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|heme iron polypeptide|Drug|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|RPL29 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|REG3A gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|RPL29 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|ST13 gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP gene|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|HHIP wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hip
null|REG3A wt Allele|Finding|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|Procedure on hip|Procedure|false|false|C0022122;C0228391;C0019552;C4299095|hipnull|Structure of habenulopeduncular tract|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0021885;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Hip structure|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0021885;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Lower extremity>Hip|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0021885;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hip
null|Bone structure of ischium|Anatomy|false|false|C1430701;C0529134;C1505163;C1654726;C0021885;C1292890;C1704840;C1337104;C1538823;C1423009;C1335638;C3538851;C1709823;C4284725|hipnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Full|Modifier|false|false||fullnull|Details|Modifier|false|false||detailsnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Operative report|Finding|false|false||operative reportnull|Operative|Time|false|false||operativenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Satisfactory - Patient Condition Code|Finding|false|false||satisfactorynull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Anesthesia substance|Drug|false|false||anesthesianull|null|Finding|false|false||anesthesia
null|Absence of sensation|Finding|false|false||anesthesianull|Anesthesia procedures|Procedure|false|false||anesthesia
null|Dental anesthesia|Procedure|false|false||anesthesianull|null|Attribute|false|false||anesthesianull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Initially|Time|false|false||initiallynull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C4284232;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false|C0226896|medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Patient's home|Device|false|false||patient's homenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Hospitalization|Procedure|false|false||hospitalizationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Discharge to home|Procedure|false|false||discharge to homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Home with services|Finding|false|false||home with servicesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|Appropriate|Modifier|false|false||appropriatenull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|null|Modifier|false|false||unremarkablenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919;C4284232|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false|C0226896|medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Surgical incisions|Procedure|false|false||incisionsnull|Cleaning (activity)|Event|false|false||cleannull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Urination|Finding|false|false|C0021853|voiding
null|Voids|Finding|false|false|C0021853|voidingnull|Moving|Finding|false|false|C0021853|movingnull|Intestines|Anatomy|false|false|C0560560;C0042034;C4067975|bowelsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Weight-Bearing state|Subject|false|false||weightbearingnull|Left lower extremity|Anatomy|false|false|C1552822;C2003888|left lower extremitynull|Table Cell Horizontal Align - left|Finding|false|false|C0230416;C0023216|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower Extremity|Anatomy|false|false|C2003888;C1552822|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802;C0023216;C0230416|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|DVT prophylaxis|Procedure|false|false|C5239664|DVT prophylaxisnull|Deep thrombophlebitis|Disorder|false|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|false|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0199176;C2926618;C0149871;C0151950;C0853245|DVTnull|null|Attribute|false|false|C5239664|DVTnull|Prophylactic treatment|Procedure|false|false|C5239664|prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Extended Priority Codes - Routine|Finding|false|false||routine
null|Report priority - Routine|Finding|false|false||routine
null|Admission Type - Routine|Finding|false|false||routine
null|Level of Care - Routine|Finding|false|false||routine
null|Processing priority - Routine|Finding|false|false||routine
null|Referral priority - Routine|Finding|false|false||routinenull|Routine coag|Procedure|false|false||routinenull|Priority - Routine|Time|false|false||routinenull|Routine|Modifier|false|false||routinenull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Course|Time|false|false||coursenull|Indication of (contextual qualifier)|Finding|false|false||reasonsnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Appropriate|Modifier|false|false||appropriatenull|Follow-Up Care|Procedure|false|false||follow-up carenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Ready for discharge|Finding|false|false||readiness for dischargenull|Readiness for discharge|Attribute|false|false||readiness for dischargenull|Readiness|Finding|false|false||readinessnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Lactaid|Drug|false|false||Lactaid
null|Lactaid|Drug|false|false||Lactaid
null|Lactaid|Drug|false|false||Lactaidnull|Lactaid Pharmaceuticals|Entity|false|false||Lactaidnull|lactase|Drug|false|false||lactase
null|GLB1 protein, human|Drug|false|false||lactase
null|GLB1 protein, human|Drug|false|false||lactase
null|lactase|Drug|false|false||lactase
null|lactase|Drug|false|false||lactasenull|LCT gene|Finding|false|false||lactasenull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|calcium citrate|Drug|false|false||Calcium Citrate
null|calcium citrate|Drug|false|false||Calcium Citratenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|citrate|Drug|false|false||Citrate
null|citrate|Drug|false|false||Citrate
null|Citrates|Drug|false|false||Citratenull|Citrate measurement|Procedure|false|false||Citratenull|calcium citrate|Drug|false|false||calcium citrate
null|calcium citrate|Drug|false|false||calcium citratenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|citrate|Drug|false|false||citrate
null|citrate|Drug|false|false||citrate
null|Citrates|Drug|false|false||citratenull|Citrate measurement|Procedure|false|false||citratenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Once a day, at bedtime|Time|false|false||QHSnull|enoxaparin|Drug|false|false||enoxaparin
null|enoxaparin|Drug|false|false||enoxaparinnull|Syringes|Device|false|false||Syringenull|Syringe (unit of presentation)|LabModifier|false|false||Syringe
null|Syringe Dosing Unit|LabModifier|false|false||Syringenull|refill|Finding|false|false||Refillsnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1422467;C1527415|mouth
null|Oral region|Anatomy|false|false|C1422467;C1527415|mouthnull|CIAO3 gene|Finding|false|false|C0230028;C0226896|PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|calcium citrate|Drug|false|false||Calcium Citrate
null|calcium citrate|Drug|false|false||Calcium Citratenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|citrate|Drug|false|false||Citrate
null|citrate|Drug|false|false||Citrate
null|Citrates|Drug|false|false||Citratenull|Citrate measurement|Procedure|false|false||Citratenull|calcium citrate|Drug|false|false||calcium citrate
null|calcium citrate|Drug|false|false||calcium citratenull|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|calcium|Drug|false|false||calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||calcium
null|Calcium, Dietary|Drug|false|false||calcium
null|Calcium [EPC]|Drug|false|false||calcium
null|Calcium Drug Class|Drug|false|false||calciumnull|Calcium metabolic function|Finding|false|false||calciumnull|Calcium measurement|Procedure|false|false||calciumnull|citrate|Drug|false|false||citrate
null|citrate|Drug|false|false||citrate
null|Citrates|Drug|false|false||citratenull|Citrate measurement|Procedure|false|false||citratenull|vitamin D3|Drug|false|false||vitamin D3
null|vitamin D3|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3
null|cholecalciferol|Drug|false|false||vitamin D3null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|Lactaid|Drug|false|false||Lactaid
null|Lactaid|Drug|false|false||Lactaid
null|Lactaid|Drug|false|false||Lactaidnull|Lactaid Pharmaceuticals|Entity|false|false||Lactaidnull|lactase|Drug|false|false||lactase
null|GLB1 protein, human|Drug|false|false||lactase
null|GLB1 protein, human|Drug|false|false||lactase
null|lactase|Drug|false|false||lactase
null|lactase|Drug|false|false||lactasenull|LCT gene|Finding|false|false||lactasenull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin preparation|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitamins
null|Multivitamin Drug Class|Drug|false|false||Multivitaminsnull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Valgus deformity|Disorder|false|false|C0015815|valgusnull|Valgus <Valginae>|Entity|false|false||valgusnull|Valgus position|Modifier|false|false||valgusnull|Impacted tooth|Disorder|false|false|C0015815|impactednull|Impacted|Finding|false|false|C0015815|impactednull|Femoral Neck Fractures|Disorder|false|false|C0015815;C0027530;C3159206;C0015811|femoral neck fracturenull|Structure of neck of femur|Anatomy|false|false|C0262414;C0015806;C0333125;C0042282;C0812434;C0684335;C0016658;C0040456|femoral necknull|Femur|Anatomy|false|false|C0015806|femoralnull|Fracture of cervical spine|Disorder|false|false|C0015815;C0027530;C3159206|neck fracturenull|Passive joint movement of neck (finding)|Finding|false|false|C0015815;C0027530;C3159206|neck
null|Neck problem|Finding|false|false|C0015815;C0027530;C3159206|necknull|dendritic spine neck|Anatomy|false|false|C0262414;C0015806;C0812434;C0684335;C0016658|neck
null|Neck|Anatomy|false|false|C0262414;C0015806;C0812434;C0684335;C0016658|necknull|Fracture|Disorder|false|false|C0015815;C0027530;C3159206|fracturenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Surgical wound|Disorder|false|false|C2338258|Incisionnull|Surgical incisions|Procedure|false|false|C2338258|Incisionnull|Cranial incision point|Anatomy|false|false|C5575035;C0332803;C0184898|Incisionnull|Well (answer to question)|Finding|false|false|C2338258|wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Dressing Dosage Form|Drug|false|false||Dressingnull|null|Finding|false|false||Dressing
null|Ability to dress|Finding|false|false||Dressingnull|Dressing patient (procedure)|Procedure|false|false||Dressing
null|Dressing of skin or wound|Procedure|false|false||Dressingnull|Medical dressing|Device|false|false||Dressing
null|Dress (garment)|Device|false|false||Dressing
null|Wound Dressings (device)|Device|false|false||Dressingnull|Dressing (unit of presentation)|LabModifier|false|false||Dressingnull|Cleaning (activity)|Event|false|false||cleannull|Febrile infection related epilepsy syndrome|Disorder|false|false||Firesnull|Fire (physical force)|Phenomenon|false|false||Firesnull|fire disaster|Event|false|false||Firesnull|Ceramide Glucosyltransferase, human|Drug|false|false||GCS
null|GCLC protein, human|Drug|false|false||GCS
null|GCLC protein, human|Drug|false|false||GCS
null|Ceramide Glucosyltransferase, human|Drug|false|false||GCSnull|GCLC wt Allele|Finding|false|false||GCS
null|UGCG gene|Finding|false|false||GCS
null|GCLC gene|Finding|false|false||GCS
null|UGCG wt Allele|Finding|false|false||GCSnull|Spatial Distribution|Modifier|false|false||distributionsnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Instructions|Finding|false|false||INSTRUCTIONS
null|Instruction [Publication Type]|Finding|false|false||INSTRUCTIONSnull|null|Attribute|false|false||INSTRUCTIONSnull|Orthopedic Surgical Procedures|Procedure|false|false||ORTHOPAEDIC SURGERYnull|Orthopedics|Title|false|false||ORTHOPAEDICnull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Orthopedic Rehabilitation Surgery|Procedure|false|false||orthopedic surgery
null|Orthopedic Surgical Procedures|Procedure|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedic surgerynull|Orthopedics|Title|false|false||orthopedicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Feel Tired question|Finding|false|false||feel tired
null|Feeling tired|Finding|false|false||feel tirednull|Feelings|Finding|false|false||feelnull|Feel Tired question|Finding|false|false||tired
null|Fatigue|Finding|false|false||tired
null|Feeling tired|Finding|false|false||tirednull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Feelings|Finding|false|false||feelingnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|day|Time|false|false||daysnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Resume - Remote control command|Finding|false|false||Resume
null|Curriculum Vitae|Finding|false|false||Resume
null|resume - DataOperation|Finding|false|false||Resumenull|Regular|Modifier|false|false||regularnull|activities (history)|Finding|false|false||activitiesnull|Activities|Event|false|false||activitiesnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Precaution|Finding|false|false||precautionsnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Activity (animal life circumstance)|Finding|false|false||ACTIVITY
null|Physical activity|Finding|false|false||ACTIVITYnull|Activities|Event|false|false||ACTIVITYnull|null|Modifier|false|false||ACTIVITYnull|Weight-Bearing state|Subject|false|false||WEIGHT BEARINGnull|infant weight for previous delivery (history)|Finding|false|false||WEIGHT
null|Weight symptom (finding)|Finding|false|false||WEIGHTnull|Weighing patient|Procedure|false|false||WEIGHTnull|null|Attribute|false|false||WEIGHTnull|Body Weight|Subject|false|false||WEIGHTnull|Importance Weight|Modifier|false|false||WEIGHTnull|Weight|LabModifier|false|false||WEIGHTnull|Bearing Device|Device|false|false||BEARINGnull|Weight-Bearing state|Subject|false|false||Weightbearingnull|Left lower extremity|Anatomy|false|false|C1552822|left lower extremitynull|Table Cell Horizontal Align - left|Finding|false|false|C0023216;C0230416|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower Extremity|Anatomy|false|false|C1552822|lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Around the Clock|Time|false|false||around the clocknull|CLOCK protein, human|Drug|false|false||clock
null|CLOCK protein, human|Drug|false|false||clocknull|CLOCK gene|Finding|false|false||clocknull|Clock Device|Device|false|false||clocknull|Drugs, Non-Prescription|Drug|false|false||over the counternull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Weaning|Finding|false|false||weannull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|1 Week|Time|false|false||1 weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Example|Finding|false|false||examplenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|3 Hours|Time|false|false||3 hoursnull|Hour|Time|false|false||hoursnull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|4 Hours|Time|false|false||4 hoursnull|Hour|Time|false|false||hoursnull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|12 hours (qualifier value)|Time|false|false||12 hoursnull|Hour|Time|false|false||hoursnull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|Before Bedtime|Time|false|false||before bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|1 Day|Time|false|false||1 daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Then - dosing instruction fragment|Finding|false|false||Thennull|Then|Time|false|false||Thennull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Regulation|Event|false|false||regulationsnull|regulatory|Entity|false|false||regulationsnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|More|LabModifier|false|false||morenull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Appointments|Event|false|false||appointmentnull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Authorization Mode - Phone|Finding|false|false||phone
null|Visit User Code - Phone|Finding|false|false||phone
null|Telephone Number|Finding|false|false||phone
null|MDFAttributeType - Phone|Finding|false|false||phonenull|Telephone|Device|false|false||phonenull|Person location type - Phone|Modifier|false|false||phonenull|Narcotics|Drug|false|false||Narcotic
null|Narcotics|Drug|false|false||Narcoticnull|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relieversnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Constipation|Finding|false|false||constipationnull|Eyeglasses|Device|false|false||glassesnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Daily|Time|false|false||dailynull|Bowel Regimen|Procedure|false|false|C0021853|bowel regimennull|Intestines|Anatomy|false|false|C5979615|bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Prescription list|Finding|false|false||prescription listnull|null|Attribute|false|false||prescription listnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Disorder|false|false||medsnull|Medications|Finding|false|false||medsnull|sennosides, USP|Drug|false|false||senna
null|sennosides, USP|Drug|false|false||sennanull|Senna alexandrina|Entity|false|false||senna
null|Senna Plant|Entity|false|false||sennanull|Colace|Drug|false|false||colace
null|Colace|Drug|false|false||colacenull|Miralax|Drug|false|false||miralax
null|Miralax|Drug|false|false||miralaxnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Motor Vehicles|Device|false|false||motor vehiclenull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Drug vehicle|Drug|false|false||vehiclenull|Vehicle (transportation)|Device|false|false||vehiclenull|operate|Finding|false|false||operatenull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Pain Relieve brand of acetaminophen|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relievers
null|Analgesics|Drug|false|false||pain relieversnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Physicians|Subject|false|false||physiciansnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|ANTICOAGULATION (finding)|Finding|false|false||ANTICOAGULATION
null|Anticoagulation function|Finding|false|false||ANTICOAGULATION
null|Decreased Coagulation Activity [PE]|Finding|false|false||ANTICOAGULATIONnull|Anticoagulation Therapy|Procedure|false|false||ANTICOAGULATIONnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|Daily|Time|false|false||dailynull|4 Weeks|Time|false|false||4 weeksnull|week|Time|false|false||weeksnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions