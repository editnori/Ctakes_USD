 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|156,164|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|179,186|false|false|false|C0009214|codeine|Codeine
Event|Event|Allergies|189,198|false|false|false|||Attending
Finding|Functional Concept|Allergies|189,198|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|223,233|false|false|false|||Difficulty
Finding|Finding|Chief Complaint|223,233|false|false|false|C1299586|Has difficulty doing (qualifier value)|Difficulty
Finding|Organism Function|Chief Complaint|234,246|false|false|false|C0004048|Inspiration (function)|in breathing
Attribute|Clinical Attribute|Chief Complaint|237,246|false|false|false|C5885990||breathing
Event|Event|Chief Complaint|237,246|false|false|false|||breathing
Finding|Finding|Chief Complaint|237,246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Chief Complaint|237,246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Chief Complaint|237,246|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Chief Complaint|237,246|false|false|false|C1160636|respiratory system process|breathing
Finding|Classification|Chief Complaint|249,254|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|255,263|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|255,263|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|267,285|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|276,285|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|276,285|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|276,285|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|276,285|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|276,285|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Body Substance|History of Present Illness|327,334|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|327,334|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|327,334|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|344,348|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|344,348|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|349,352|false|false|false|||old
Event|Event|History of Present Illness|367,374|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|367,374|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|367,377|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|History of Present Illness|378,383|false|false|false|C0007131||NSCLC
Event|Event|History of Present Illness|378,383|false|false|false|||NSCLC
Attribute|Clinical Attribute|History of Present Illness|386,391|false|false|false|C1300072|Tumor stage|stage
Event|Event|History of Present Illness|400,408|false|false|false|||presents
Event|Event|History of Present Illness|414,423|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|414,433|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|414,433|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|427,433|false|false|false|C0225386|Breath|breath
Finding|Body Substance|History of Present Illness|441,448|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|441,448|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|441,448|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|466,471|false|false|false|||state
Finding|Functional Concept|History of Present Illness|466,471|false|false|false|C1442792|State|state
Finding|Finding|History of Present Illness|466,481|false|false|false|C0683314|personal health|state of health
Event|Event|History of Present Illness|475,481|false|false|false|||health
Finding|Idea or Concept|History of Present Illness|475,481|false|false|false|C0018684|Health|health
Event|Event|History of Present Illness|508,517|false|false|false|||admission
Procedure|Health Care Activity|History of Present Illness|508,517|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|History of Present Illness|527,532|false|false|false|||began
Event|Event|History of Present Illness|536,540|false|false|false|||feel
Finding|Finding|History of Present Illness|541,549|false|false|false|C2984079|Somewhat|somewhat
Event|Event|History of Present Illness|550,555|false|false|false|||short
Event|Event|History of Present Illness|560,566|false|false|false|||breath
Finding|Body Substance|History of Present Illness|560,566|false|false|false|C0225386|Breath|breath
Finding|Idea or Concept|History of Present Illness|573,577|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|History of Present Illness|592,601|false|false|false|||sensation
Finding|Finding|History of Present Illness|592,601|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|592,601|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|592,601|false|false|false|C2229507|sensory exam|sensation
Event|Event|History of Present Illness|602,611|false|false|false|||persisted
Event|Event|History of Present Illness|621,627|false|false|false|||became
Event|Event|History of Present Illness|628,637|false|false|false|||concerned
Event|Event|History of Present Illness|649,656|false|false|false|||reports
Finding|Idea or Concept|History of Present Illness|663,666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|663,666|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|History of Present Illness|667,674|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|667,674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|667,674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|667,674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|667,677|false|false|false|C0262926|Medical History|history of
Drug|Organic Chemical|History of Present Illness|696,701|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|696,701|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|696,701|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|696,701|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|704,710|false|false|false|||Denies
Finding|Sign or Symptom|History of Present Illness|711,715|true|false|false|C0221423|Illness (finding)|sick
Event|Event|History of Present Illness|716,724|true|false|false|||contacts
Procedure|Health Care Activity|History of Present Illness|716,724|true|false|false|C4036459|Contacts|contacts
Event|Event|History of Present Illness|733,739|true|false|false|||travel
Finding|Daily or Recreational Activity|History of Present Illness|733,739|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|733,739|true|false|false|C1555670|travel charge|travel
Finding|Finding|History of Present Illness|744,753|false|false|false|C1532253|Sedentary lifestyle|sedentary
Finding|Finding|History of Present Illness|744,763|false|false|false|C1532253|Sedentary lifestyle|sedentary lifestyle
Event|Event|History of Present Illness|754,763|false|false|false|||lifestyle
Finding|Social Behavior|History of Present Illness|754,763|false|false|false|C0023676|Life Style|lifestyle
Event|Event|History of Present Illness|770,776|false|false|false|||denied
Anatomy|Body Location or Region|History of Present Illness|777,782|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|777,782|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|777,787|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|777,787|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|783,787|true|false|false|C2598155||pain
Event|Event|History of Present Illness|783,787|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|783,787|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|783,787|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|789,794|true|false|false|||fever
Finding|Finding|History of Present Illness|789,794|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|789,794|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|796,802|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|796,802|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|805,814|false|false|false|||dizziness
Finding|Sign or Symptom|History of Present Illness|805,814|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Event|Event|History of Present Illness|816,831|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|816,831|false|false|false|C0220870|Lightheadedness|lightheadedness
Event|Event|History of Present Illness|835,842|false|false|false|||syncope
Finding|Sign or Symptom|History of Present Illness|835,842|false|false|false|C0039070|Syncope|syncope
Event|Event|History of Present Illness|849,858|false|false|false|||presented
Event|Event|History of Present Illness|884,889|false|false|false|||found
Event|Event|History of Present Illness|896,903|false|false|false|||hypoxic
Finding|Pathologic Function|History of Present Illness|896,903|false|false|false|C0242184|Hypoxia|hypoxic
Finding|Finding|History of Present Illness|915,926|false|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|History of Present Illness|918,926|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|History of Present Illness|923,926|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|History of Present Illness|923,926|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|History of Present Illness|923,926|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|History of Present Illness|923,926|false|false|false|||air
Finding|Finding|History of Present Illness|923,926|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|History of Present Illness|923,926|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|History of Present Illness|923,926|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|History of Present Illness|951,957|false|false|false|||placed
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|983,987|false|false|false|C0312448|short-acting thyroid stimulator|sats
Drug|Hormone|History of Present Illness|983,987|false|false|false|C0312448|short-acting thyroid stimulator|sats
Event|Event|History of Present Illness|983,987|false|false|false|||sats
Finding|Finding|History of Present Illness|999,1003|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|History of Present Illness|999,1003|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|History of Present Illness|999,1003|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|History of Present Illness|1011,1019|false|false|false|||Attempts
Event|Event|History of Present Illness|1033,1037|false|false|false|||wean
Event|Event|History of Present Illness|1063,1075|false|false|false|||unsuccessful
Event|Event|History of Present Illness|1088,1095|false|false|false|||satting
Event|Event|History of Present Illness|1106,1108|false|false|false|||NC
Event|Event|History of Present Illness|1116,1124|false|false|false|||remained
Event|Event|History of Present Illness|1125,1133|false|false|false|||afebrile
Finding|Finding|History of Present Illness|1125,1133|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|History of Present Illness|1152,1157|false|false|false|||found
Anatomy|Cell|History of Present Illness|1166,1169|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|1166,1169|false|false|false|||WBC
Drug|Antibiotic|History of Present Illness|1204,1216|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|History of Present Illness|1204,1216|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|History of Present Illness|1204,1216|false|false|false|||levofloxacin
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1221,1231|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|History of Present Illness|1221,1231|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|History of Present Illness|1221,1231|false|false|false|||vancomycin
Procedure|Laboratory Procedure|History of Present Illness|1221,1231|false|false|false|C0489941|Vancomycin measurement|vancomycin
Disorder|Disease or Syndrome|History of Present Illness|1234,1239|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|History of Present Illness|1234,1239|false|false|false|||Blood
Finding|Body Substance|History of Present Illness|1234,1239|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|History of Present Illness|1241,1249|false|false|false|||cultures
Finding|Idea or Concept|History of Present Illness|1241,1249|false|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|History of Present Illness|1255,1260|false|false|false|||drawn
Drug|Antibiotic|History of Present Illness|1270,1280|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1270,1295|false|false|false|C0199779|Injection of antibiotic|antibiotic administration
Event|Event|History of Present Illness|1281,1295|false|false|false|||administration
Event|Occupational Activity|History of Present Illness|1281,1295|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1281,1295|false|false|false|C1533734|Administration (procedure)|administration
Event|Event|History of Present Illness|1298,1301|true|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1298,1301|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1311,1315|true|false|false|||show
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|1316,1319|true|true|false|C0600500|Peptide Nucleic Acids|PNA
Event|Event|History of Present Illness|1316,1319|true|false|false|||PNA
Event|Event|History of Present Illness|1325,1337|false|false|false|||demonstrated
Event|Event|History of Present Illness|1338,1349|false|false|false|||progression
Finding|Functional Concept|History of Present Illness|1338,1349|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|History of Present Illness|1338,1349|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Anatomy|Body Location or Region|History of Present Illness|1359,1363|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1359,1363|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|History of Present Illness|1359,1363|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|History of Present Illness|1359,1363|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|History of Present Illness|1359,1370|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|History of Present Illness|1364,1370|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|History of Present Illness|1364,1370|false|false|false|||cancer
Attribute|Clinical Attribute|History of Present Illness|1390,1397|true|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|History of Present Illness|1390,1397|true|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|History of Present Illness|1393,1397|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1393,1397|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1393,1397|true|false|false|C0362076|Problems with head|head
Event|Event|History of Present Illness|1393,1397|true|false|false|||head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1393,1397|true|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|1401,1405|false|false|false|||rule
Disorder|Neoplastic Process|History of Present Illness|1410,1420|true|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastases
Event|Event|History of Present Illness|1410,1420|true|false|false|||metastases
Finding|Finding|History of Present Illness|1410,1420|true|false|false|C1513183|Metastatic Lesion|metastases
Event|Event|History of Present Illness|1433,1441|false|false|false|||negative
Finding|Classification|History of Present Illness|1433,1441|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1433,1441|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1433,1441|false|false|false|C5237010|Expression Negative|negative
Event|Event|History of Present Illness|1447,1455|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1447,1455|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1447,1455|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1447,1455|false|false|false|C4706767|Transfer (immobility management)|transfer
Procedure|Health Care Activity|History of Present Illness|1447,1464|false|false|false|C0030704|Patient Transfer|transfer, patient
Event|Event|History of Present Illness|1457,1464|false|false|false|||patient
Finding|Body Substance|History of Present Illness|1457,1464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1457,1464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1457,1464|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1469,1477|false|false|false|||afebrile
Finding|Finding|History of Present Illness|1469,1477|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|History of Present Illness|1529,1532|false|false|false|||NRB
Event|Event|History of Present Illness|1540,1548|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1540,1548|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1540,1548|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1540,1548|false|false|false|C4706767|Transfer (immobility management)|transfer
Anatomy|Body Space or Junction|History of Present Illness|1556,1559|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Finding|Intellectual Product|History of Present Illness|1556,1559|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Finding|Body Substance|History of Present Illness|1565,1572|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1565,1572|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1565,1572|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1577,1583|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1577,1583|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|History of Present Illness|1588,1599|false|false|false|||comfortable
Finding|Finding|History of Present Illness|1588,1599|false|false|false|C5546696|Feeling comfortable|comfortable
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1603,1607|false|false|false|C0312448|short-acting thyroid stimulator|Sats
Drug|Hormone|History of Present Illness|1603,1607|false|false|false|C0312448|short-acting thyroid stimulator|Sats
Event|Event|History of Present Illness|1603,1607|false|false|false|||Sats
Event|Event|History of Present Illness|1623,1625|false|false|false|||NC
Finding|Finding|History of Present Illness|1634,1638|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|History of Present Illness|1634,1638|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|History of Present Illness|1634,1638|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|History of Present Illness|1639,1643|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1639,1643|false|false|false|C0806140|Flow|flow
Anatomy|Body Location or Region|History of Present Illness|1651,1655|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|History of Present Illness|1651,1655|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|History of Present Illness|1651,1655|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Space or Junction|History of Present Illness|1668,1671|false|false|false|C0262327|rostral sulcus|ROS
Drug|Biologically Active Substance|History of Present Illness|1668,1671|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Element, Ion, or Isotope|History of Present Illness|1668,1671|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Organic Chemical|History of Present Illness|1668,1671|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Drug|Pharmacologic Substance|History of Present Illness|1668,1671|false|false|false|C0162772;C0289313|Reactive Oxygen Species;rosiglitazone|ROS
Event|Event|History of Present Illness|1668,1671|false|false|false|||ROS
Finding|Gene or Genome|History of Present Illness|1668,1671|false|false|false|C0812281;C1709820|ROS1 gene;ROS1 wt Allele|ROS
Procedure|Health Care Activity|History of Present Illness|1668,1671|false|false|false|C0489633|Review of systems (procedure)|ROS
Finding|Body Substance|History of Present Illness|1677,1684|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1677,1684|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1677,1684|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1685,1691|true|false|false|||denies
Event|Event|History of Present Illness|1696,1702|true|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|1696,1702|true|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|1704,1710|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1704,1710|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|1712,1718|true|false|false|C0944911||weight
Event|Event|History of Present Illness|1712,1718|true|false|false|||weight
Finding|Finding|History of Present Illness|1712,1718|true|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|1712,1718|true|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|1712,1718|true|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|1712,1725|true|false|false|C0005911|Body Weight Changes|weight change
Event|Event|History of Present Illness|1719,1725|true|false|false|||change
Finding|Functional Concept|History of Present Illness|1719,1725|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1719,1725|true|false|false|C4319952|Change - procedure|change
Attribute|Clinical Attribute|History of Present Illness|1728,1734|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1728,1734|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1728,1734|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1736,1744|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1736,1744|false|false|false|C0042963|Vomiting|vomiting
Anatomy|Body Location or Region|History of Present Illness|1746,1755|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1746,1760|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1756,1760|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1756,1760|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1756,1760|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1756,1760|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1762,1770|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|1762,1770|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1762,1770|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|1772,1784|false|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|1772,1784|false|false|false|C0009806|Constipation|constipation
Event|Event|History of Present Illness|1787,1793|false|false|false|||melena
Finding|Pathologic Function|History of Present Illness|1787,1793|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|History of Present Illness|1795,1807|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|History of Present Illness|1795,1807|false|false|false|||hematochezia
Finding|Sign or Symptom|History of Present Illness|1795,1807|false|false|false|C1321898|Blood in stool|hematochezia
Anatomy|Body Location or Region|History of Present Illness|1809,1814|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1809,1814|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1809,1819|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1809,1819|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1815,1819|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1815,1819|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1815,1819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1815,1819|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1821,1830|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|1821,1830|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1821,1830|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|History of Present Illness|1832,1835|false|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Event|Event|History of Present Illness|1832,1835|false|false|false|||PND
Finding|Gene or Genome|History of Present Illness|1832,1835|false|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Anatomy|Body Location or Region|History of Present Illness|1837,1842|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|1837,1842|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1844,1853|false|false|false|C0015385|Limb structure|extremity
Finding|Pathologic Function|History of Present Illness|1844,1859|false|false|false|C0085649|Peripheral edema|extremity edema
Attribute|Clinical Attribute|History of Present Illness|1854,1859|false|false|false|C1717255||edema
Event|Event|History of Present Illness|1854,1859|false|false|false|||edema
Finding|Pathologic Function|History of Present Illness|1854,1859|false|false|false|C0013604|Edema|edema
Drug|Organic Chemical|History of Present Illness|1861,1866|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1861,1866|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1861,1866|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1861,1866|false|false|false|C0010200|Coughing|cough
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1868,1875|false|false|false|C0042027|Urinary tract|urinary
Finding|Finding|History of Present Illness|1868,1885|false|false|false|C0042023|Increased frequency of micturition|urinary frequency
Event|Event|History of Present Illness|1876,1885|false|false|false|||frequency
Finding|Intellectual Product|History of Present Illness|1876,1885|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|History of Present Illness|1887,1894|false|false|false|||urgency
Event|Event|History of Present Illness|1896,1903|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|1896,1903|false|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|1906,1921|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|1906,1921|false|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Finding|History of Present Illness|1923,1927|false|false|false|C0016928|Gait|gait
Event|Event|History of Present Illness|1928,1940|false|false|false|||unsteadiness
Finding|Finding|History of Present Illness|1928,1940|false|false|false|C0427108|General unsteadiness|unsteadiness
Event|Event|History of Present Illness|1948,1956|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1948,1956|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Attribute|Clinical Attribute|History of Present Illness|1958,1964|false|false|false|C2707266||vision
Event|Event|History of Present Illness|1958,1964|false|false|false|||vision
Finding|Organism Function|History of Present Illness|1958,1964|false|false|false|C0042789|Vision|vision
Event|Event|History of Present Illness|1966,1973|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|1966,1973|false|false|false|C0392747|Changing|changes
Event|Event|History of Present Illness|1975,1983|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|1975,1983|false|false|false|C0018681|Headache|headache
Disorder|Disease or Syndrome|History of Present Illness|1985,1989|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|History of Present Illness|1985,1989|false|false|false|||rash
Finding|Pathologic Function|History of Present Illness|1985,1989|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|1985,1989|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Anatomy|Body System|History of Present Illness|1993,1997|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|History of Present Illness|1993,1997|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|History of Present Illness|1993,1997|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|History of Present Illness|1993,1997|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|History of Present Illness|1993,1997|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|History of Present Illness|1993,2005|false|false|false|C0421292|Skin symptom change|skin changes
Event|Event|History of Present Illness|1998,2005|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|1998,2005|false|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|Past Medical History|2038,2041|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2038,2041|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|2038,2041|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Past Medical History|2038,2041|false|false|false|||CAD
Finding|Gene or Genome|Past Medical History|2038,2041|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|2038,2041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|2038,2041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2038,2041|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Past Medical History|2057,2061|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2057,2061|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Disorder|Disease or Syndrome|Past Medical History|2066,2078|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|2066,2078|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Past Medical History|2079,2091|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Event|Event|Past Medical History|2079,2091|false|false|false|||Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|2092,2095|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|2092,2095|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|Past Medical History|2092,2095|false|false|false|||CVA
Finding|Functional Concept|Past Medical History|2103,2107|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|Past Medical History|2108,2117|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|Past Medical History|2126,2133|false|false|false|||infarct
Finding|Pathologic Function|Past Medical History|2126,2133|false|false|false|C0021308|Infarction|infarct
Disorder|Disease or Syndrome|Past Medical History|2141,2161|false|false|false|C0024437;C0242383|Age related macular degeneration;Macular degeneration|Macular Degeneration
Event|Event|Past Medical History|2149,2161|false|false|false|||Degeneration
Finding|Functional Concept|Past Medical History|2149,2161|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degeneration
Finding|Pathologic Function|Past Medical History|2149,2161|false|false|false|C0011164;C1880269|Abnormal degeneration;biologic degeneration|Degeneration
Disorder|Neoplastic Process|Past Medical History|2162,2167|false|false|false|C0007131||NSCLC
Event|Event|Past Medical History|2162,2167|false|false|false|||NSCLC
Attribute|Clinical Attribute|Past Medical History|2169,2174|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|2169,2177|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Neoplastic Process|Past Medical History|2179,2187|false|false|false|C0027651|Neoplasms|oncology
Procedure|Health Care Activity|Past Medical History|2179,2187|false|false|false|C1555459|oncology services|oncology
Event|Event|Past Medical History|2188,2195|false|false|false|||history
Finding|Conceptual Entity|Past Medical History|2188,2195|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Past Medical History|2188,2195|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Past Medical History|2188,2195|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|Past Medical History|2212,2221|false|false|false|||presented
Finding|Functional Concept|Past Medical History|2242,2247|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2254,2263|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Past Medical History|2254,2263|false|false|false|C2707265||pulmonary
Finding|Finding|Past Medical History|2254,2263|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Past Medical History|2265,2275|false|false|false|||infiltrate
Finding|Functional Concept|Past Medical History|2265,2275|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Past Medical History|2265,2275|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Past Medical History|2265,2275|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Finding|Past Medical History|2283,2292|false|false|false|C0445356|Unrelated (finding)|unrelated
Anatomy|Tissue|Past Medical History|2293,2303|false|false|false|C0027061|Myocardium|myocardial
Attribute|Clinical Attribute|Past Medical History|2293,2314|false|false|false|C2926063||myocardial infarction
Disorder|Disease or Syndrome|Past Medical History|2293,2314|false|false|false|C0027051|Myocardial Infarction|myocardial infarction
Event|Event|Past Medical History|2304,2314|false|false|false|||infarction
Finding|Pathologic Function|Past Medical History|2304,2314|false|false|false|C0021308|Infarction|infarction
Event|Event|Past Medical History|2338,2347|false|false|false|||confirmed
Disorder|Neoplastic Process|Past Medical History|2348,2362|false|false|false|C0001418;C5551397|Adenocarcinoma;Malignant adenomatous neoplasm|adenocarcinoma
Event|Event|Past Medical History|2348,2362|false|false|false|||adenocarcinoma
Event|Event|Past Medical History|2371,2378|false|false|false|||pattern
Event|Event|Past Medical History|2382,2397|false|false|false|||stainpositivity
Event|Event|Past Medical History|2398,2408|false|false|false|||consistent
Finding|Idea or Concept|Past Medical History|2398,2408|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Past Medical History|2398,2413|false|false|false|C0332290|Consistent with|consistent with
Anatomy|Body Location or Region|Past Medical History|2414,2418|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2414,2418|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Past Medical History|2414,2418|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Past Medical History|2414,2418|false|false|false|C0740941|Lung Problem|lung
Event|Event|Past Medical History|2419,2425|false|false|false|||origin
Finding|Classification|Past Medical History|2419,2425|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Intellectual Product|Past Medical History|2419,2425|false|false|false|C0079946;C1550512|National origin;Participation Type - origin|origin
Finding|Gene or Genome|Past Medical History|2427,2430|false|false|false|C1416745;C3272782|KRT7 gene;KRT7 wt Allele|CK7
Event|Event|Past Medical History|2436,2439|false|false|false|||TTF
Finding|Gene or Genome|Past Medical History|2436,2439|false|false|false|C1332112;C1705840|RHOH gene;RHOH wt Allele|TTF
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2436,2439|false|false|false|C4087167|Tumour treating fields therapy|TTF
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2436,2441|false|false|false|C0084785;C1452466;C1610981|NKX2-1 protein, human;TTF1 protein, human;thyroid transcription factor 1|TTF-1
Drug|Biologically Active Substance|Past Medical History|2436,2441|false|false|false|C0084785;C1452466;C1610981|NKX2-1 protein, human;TTF1 protein, human;thyroid transcription factor 1|TTF-1
Finding|Gene or Genome|Past Medical History|2436,2441|false|false|false|C1384616;C2347318;C3811254|NKX2-1 gene;NKX2-1 wt Allele;TTF1 wt Allele|TTF-1
Disorder|Cell or Molecular Dysfunction|Past Medical History|2442,2450|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Past Medical History|2442,2450|false|false|false|||positive
Finding|Classification|Past Medical History|2442,2450|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Past Medical History|2442,2450|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Attribute|Clinical Attribute|Past Medical History|2461,2466|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|2461,2469|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Neoplastic Process|Past Medical History|2461,2495|false|false|false|C0278987|Metastatic non-small cell lung cancer|stage IV nonsmall cell lung cancer
Anatomy|Cell|Past Medical History|2479,2483|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Past Medical History|2479,2483|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Past Medical History|2484,2488|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2484,2488|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Past Medical History|2484,2488|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Past Medical History|2484,2488|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Past Medical History|2484,2495|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Past Medical History|2489,2495|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|2489,2495|false|false|false|||cancer
Event|Event|Past Medical History|2498,2503|false|false|false|||based
Finding|Functional Concept|Past Medical History|2520,2534|false|false|false|C1522224|Intrapulmonary Route of Administration|intrapulmonary
Event|Event|Past Medical History|2535,2542|false|false|false|||lesions
Finding|Finding|Past Medical History|2535,2542|false|false|false|C0221198|Lesion|lesions
Event|Event|Past Medical History|2556,2564|true|false|false|||evidence
Finding|Idea or Concept|Past Medical History|2556,2564|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Past Medical History|2556,2567|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Past Medical History|2568,2581|true|false|false|||extrathoracic
Drug|Pharmacologic Substance|Past Medical History|2585,2592|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Drug|Vitamin|Past Medical History|2585,2592|true|false|false|C0719205|Central brand of multivitamin with minerals|central
Event|Event|Past Medical History|2585,2592|true|false|false|||central
Procedure|Laboratory Procedure|Past Medical History|2585,2592|true|false|false|C1879652|Central Minus|central
Anatomy|Body System|Past Medical History|2585,2607|true|false|false|C3714787|Central Nervous System|central nervous system
Drug|Indicator, Reagent, or Diagnostic Aid|Past Medical History|2585,2607|true|false|false|C3540014|CENTRAL NERVOUS SYSTEM DIAGNOSTIC RADIOPHARMACEUTICALS|central nervous system
Finding|Finding|Past Medical History|2585,2619|true|false|false|C4050309|Central Nervous System Involvement|central nervous system involvement
Finding|Functional Concept|Past Medical History|2593,2600|true|false|false|C0027769;C0599851|Nervous - anatomy qualifier;Nervousness|nervous
Finding|Sign or Symptom|Past Medical History|2593,2600|true|false|false|C0027769;C0599851|Nervous - anatomy qualifier;Nervousness|nervous
Anatomy|Body System|Past Medical History|2593,2607|true|false|false|C0027763|Nervous system structure|nervous system
Drug|Pharmacologic Substance|Past Medical History|2593,2607|true|false|false|C3542961|NERVOUS SYSTEM DRUGS|nervous system
Drug|Biomedical or Dental Material|Past Medical History|2601,2607|false|false|false|C5671121|System (basic dose form)|system
Finding|Functional Concept|Past Medical History|2601,2607|false|false|false|C0449913;C5441654|System;System, LOINC Axis 4|system
Event|Event|Past Medical History|2608,2619|false|false|false|||involvement
Finding|Functional Concept|Past Medical History|2608,2619|false|false|false|C1314939|Involvement with|involvement
Disorder|Neoplastic Process|Past Medical History|2626,2636|false|false|false|C0027627;C2939419|Metastatic malignant neoplasm;Neoplasm Metastasis|metastasis
Event|Event|Past Medical History|2626,2636|false|false|false|||metastasis
Finding|Finding|Past Medical History|2626,2636|false|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Finding|Pathologic Function|Past Medical History|2626,2636|false|false|false|C1513183;C4255448|Metastasis;Metastatic Lesion|metastasis
Attribute|Clinical Attribute|Past Medical History|2646,2652|false|false|false|C5889824||Status
Event|Event|Past Medical History|2646,2652|false|false|false|||Status
Finding|Idea or Concept|Past Medical History|2646,2652|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Past Medical History|2660,2666|false|false|false|||cycles
Drug|Organic Chemical|Past Medical History|2670,2680|false|false|false|C0210657|pemetrexed|pemetrexed
Drug|Pharmacologic Substance|Past Medical History|2670,2680|false|false|false|C0210657|pemetrexed|pemetrexed
Event|Event|Past Medical History|2670,2680|false|false|false|||pemetrexed
Event|Event|Past Medical History|2740,2751|false|false|false|||complicated
Disorder|Disease or Syndrome|Past Medical History|2756,2766|false|false|false|C5779593|Cytopenia|cytopenias
Event|Event|Past Medical History|2756,2766|false|false|false|||cytopenias
Finding|Finding|Past Medical History|2756,2766|false|false|false|C0010828|Cytopenia (finding)|cytopenias
Event|Event|Past Medical History|2771,2782|false|false|false|||development
Finding|Functional Concept|Past Medical History|2771,2782|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|Past Medical History|2771,2782|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Finding|Past Medical History|2786,2806|false|false|false|C0151578;C0700225|Creatinine increased;Serum creatinine raised|increased creatinine
Drug|Biologically Active Substance|Past Medical History|2796,2806|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Past Medical History|2796,2806|false|false|false|C0010294|creatinine|creatinine
Event|Event|Past Medical History|2796,2806|false|false|false|||creatinine
Finding|Physiologic Function|Past Medical History|2796,2806|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Past Medical History|2796,2806|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Finding|Past Medical History|2796,2813|false|false|false|C0428279|Finding of creatinine level|creatinine levels
Event|Event|Past Medical History|2807,2813|false|false|false|||levels
Anatomy|Body Location or Region|Past Medical History|2823,2828|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|2823,2828|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|Past Medical History|2823,2831|false|false|false|C0202823|Chest CT|Chest CT
Event|Event|Past Medical History|2829,2831|false|false|false|||CT
Event|Event|Past Medical History|2832,2838|false|false|false|||showed
Finding|Idea or Concept|Past Medical History|2839,2846|false|false|false|C1550516|Target Awareness - partial|partial
Finding|Classification|Past Medical History|2839,2855|false|false|false|C1521726;C4723835;C5202624;C5202892;C5575501|IMWG Partial Response;ITMIG MRECIST Partial Response;RECIL PR;irPR (Immune-Related Response Criteria);partial response|partial response
Finding|Finding|Past Medical History|2839,2855|false|false|false|C1521726;C4723835;C5202624;C5202892;C5575501|IMWG Partial Response;ITMIG MRECIST Partial Response;RECIL PR;irPR (Immune-Related Response Criteria);partial response|partial response
Event|Event|Past Medical History|2847,2855|false|false|false|||response
Finding|Finding|Past Medical History|2847,2855|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Past Medical History|2847,2855|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Past Medical History|2847,2855|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Event|Event|Past Medical History|2861,2869|false|false|false|||interval
Finding|Intellectual Product|Past Medical History|2861,2869|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|Past Medical History|2871,2882|false|false|false|||improvement
Finding|Conceptual Entity|Past Medical History|2871,2882|false|false|false|C2986411|Improvement|improvement
Disorder|Disease or Syndrome|Past Medical History|2890,2903|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Past Medical History|2890,2903|false|false|false|||consolidation
Finding|Functional Concept|Past Medical History|2936,2941|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2936,2952|false|false|false|C1261075|Structure of right lower lobe of lung|right lower lobe
Anatomy|Body Location or Region|Past Medical History|2942,2947|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Past Medical History|2942,2947|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2942,2952|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2948,2952|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Past Medical History|2948,2952|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Past Medical History|2965,2974|false|false|false|||densities
Finding|Functional Concept|Past Medical History|2982,2986|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2982,2997|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|Past Medical History|2987,2992|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Past Medical History|2987,2992|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2987,2997|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2993,2997|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Past Medical History|2993,2997|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|Past Medical History|3001,3006|false|false|false|C1410088|Still|Still
Event|Event|Past Medical History|3014,3026|false|false|false|||disseminated
Anatomy|Cell Component|Past Medical History|3027,3030|false|false|false|C1621493|polyhedral organelle|BAC
Disorder|Neoplastic Process|Past Medical History|3027,3030|false|false|false|C0007120|Bronchioloalveolar Adenocarcinoma|BAC
Drug|Amino Acid, Peptide, or Protein|Past Medical History|3027,3030|false|false|false|C0004599|bacitracin|BAC
Drug|Antibiotic|Past Medical History|3027,3030|false|false|false|C0004599|bacitracin|BAC
Event|Event|Past Medical History|3027,3030|false|false|false|||BAC
Finding|Finding|Past Medical History|3027,3030|false|false|false|C0684262|Blood alcohol concentration|BAC
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3027,3030|false|false|false|C4553150|BAC Regimen|BAC
Attribute|Clinical Attribute|Past Medical History|3040,3048|false|false|false|C0881858||CT Chest
Procedure|Diagnostic Procedure|Past Medical History|3040,3048|false|false|false|C0202823|Chest CT|CT Chest
Anatomy|Body Location or Region|Past Medical History|3043,3048|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|3043,3048|false|false|false|C0741025|Chest problem|Chest
Event|Event|Past Medical History|3055,3064|false|false|false|||increased
Finding|Finding|Past Medical History|3055,3072|false|false|false|C0029053;C5779786|Decreased translucency;Density above reference range|increased density
Event|Event|Past Medical History|3065,3072|false|false|false|||density
Finding|Functional Concept|Past Medical History|3076,3081|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3076,3092|false|false|false|C1261075|Structure of right lower lobe of lung|right lower lobe
Anatomy|Body Location or Region|Past Medical History|3082,3087|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Past Medical History|3082,3087|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3082,3092|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3088,3092|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Past Medical History|3088,3092|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|Past Medical History|3093,3106|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Past Medical History|3093,3106|false|false|false|||consolidation
Event|Event|Past Medical History|3111,3119|false|false|false|||worsened
Disorder|Disease or Syndrome|Past Medical History|3143,3148|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|Past Medical History|3143,3148|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|Past Medical History|3143,3148|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|Past Medical History|3143,3148|false|false|false|C0025611|methamphetamine|glass
Event|Event|Past Medical History|3143,3148|false|false|false|||glass
Event|Event|Past Medical History|3150,3159|false|false|false|||opacities
Finding|Finding|Past Medical History|3150,3159|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|Past Medical History|3150,3159|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3167,3174|false|false|false|C0225740;C0228475;C1561517|Lingula;Lingula of cerebellum;Lingula of left lung|lingula
Event|Event|Past Medical History|3184,3194|false|false|false|||consistent
Finding|Idea or Concept|Past Medical History|3184,3194|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Past Medical History|3184,3199|false|false|false|C0332290|Consistent with|consistent with
Event|Event|Past Medical History|3200,3209|false|false|false|||worsening
Finding|Idea or Concept|Past Medical History|3200,3209|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Event|Event|Past Medical History|3220,3232|false|false|false|||disseminated
Anatomy|Cell|Past Medical History|3243,3247|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Past Medical History|3243,3247|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Past Medical History|3248,3252|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3248,3252|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Past Medical History|3248,3252|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Past Medical History|3248,3252|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Past Medical History|3248,3259|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Past Medical History|3253,3259|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|3253,3259|false|false|false|||cancer
Finding|Finding|Past Medical History|3261,3265|false|false|false|C4281574|Much|much
Finding|Finding|Past Medical History|3271,3277|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Past Medical History|3271,3277|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Past Medical History|3285,3294|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Past Medical History|3285,3294|false|false|false|||infection
Finding|Pathologic Function|Past Medical History|3285,3294|false|false|false|C3714514|Infection|infection
Anatomy|Body Location or Region|Past Medical History|3304,3309|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|3304,3309|false|false|false|C0741025|Chest problem|Chest
Procedure|Diagnostic Procedure|Past Medical History|3304,3312|false|false|false|C0202823|Chest CT|Chest CT
Finding|Finding|Past Medical History|3314,3320|false|false|false|C5202796|Intensity and Distress 1|slight
Event|Event|Past Medical History|3321,3329|true|false|false|||interval
Finding|Intellectual Product|Past Medical History|3321,3329|true|false|false|C1552654|Parameterized Data Type - Interval|interval
Event|Event|Past Medical History|3330,3341|true|false|false|||progression
Finding|Functional Concept|Past Medical History|3330,3341|true|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Past Medical History|3330,3341|true|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Past Medical History|3352,3359|true|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|3352,3359|true|false|false|||disease
Finding|Finding|Past Medical History|3364,3367|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Past Medical History|3364,3367|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|Past Medical History|3368,3373|true|false|false|||sites
Finding|Conceptual Entity|Family Medical History|3418,3424|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|Family Medical History|3418,3424|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|Family Medical History|3425,3429|false|false|false|||died
Disorder|Disease or Syndrome|Family Medical History|3437,3440|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3437,3440|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|3437,3440|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Family Medical History|3437,3440|false|false|false|||CAD
Finding|Gene or Genome|Family Medical History|3437,3440|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|3437,3440|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|3437,3440|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3437,3440|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|Family Medical History|3444,3447|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|3444,3447|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|3444,3447|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Family Medical History|3444,3447|false|false|false|||age
Finding|Idea or Concept|Family Medical History|3457,3463|false|false|false|C1546508|Relationship - Mother|mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3468,3475|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Family Medical History|3468,3475|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Family Medical History|3468,3475|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|Family Medical History|3468,3475|false|false|false|||stomach
Finding|Finding|Family Medical History|3468,3475|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3468,3475|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|Family Medical History|3477,3483|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3477,3483|false|false|false|||cancer
Disorder|Neoplastic Process|Family Medical History|3488,3500|false|false|false|C0029463;C0585442|Osteosarcoma;Osteosarcoma of bone|osteosarcoma
Event|Event|Family Medical History|3488,3500|false|false|false|||osteosarcoma
Finding|Gene or Genome|Family Medical History|3488,3500|false|false|false|C0694889|RB1 gene|osteosarcoma
Event|Event|Family Medical History|3505,3512|true|false|false|||history
Finding|Conceptual Entity|Family Medical History|3505,3512|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3505,3512|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|3505,3512|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|3505,3515|true|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Family Medical History|3516,3520|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3516,3520|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|3516,3520|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|3516,3520|true|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Family Medical History|3516,3527|true|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Family Medical History|3521,3527|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3521,3527|true|false|false|||cancer
Disorder|Neoplastic Process|Family Medical History|3521,3534|true|false|false|C0007102|Malignant tumor of colon|cancer, colon
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3529,3534|true|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|3529,3534|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|3529,3534|true|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|3529,3534|true|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|3529,3541|true|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|Family Medical History|3535,3541|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3535,3541|true|false|false|||cancer
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3546,3552|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Family Medical History|3546,3552|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Event|Event|Family Medical History|3546,3552|false|false|false|||breast
Finding|Finding|Family Medical History|3546,3552|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3546,3552|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|Family Medical History|3546,3559|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|Family Medical History|3553,3559|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3553,3559|false|false|false|||cancer
Event|Event|General Exam|3581,3590|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|3581,3590|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Anatomy|Body Location or Region|General Exam|3656,3660|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|General Exam|3656,3660|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|General Exam|3656,3660|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|General Exam|3668,3671|false|false|false|||GEN
Finding|Classification|General Exam|3668,3671|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|General Exam|3668,3671|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Finding|General Exam|3673,3677|true|false|false|C5575035|Well (answer to question)|Well
Event|Event|General Exam|3678,3687|true|false|false|||appearing
Finding|Finding|General Exam|3695,3715|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|3701,3706|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3707,3715|true|false|false|||distress
Finding|Finding|General Exam|3707,3715|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3707,3715|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3718,3723|true|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3725,3729|false|false|false|||EOMI
Event|Event|General Exam|3731,3736|false|false|false|||PERRL
Finding|Finding|General Exam|3731,3736|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Part, Organ, or Organ Component|General Exam|3738,3744|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|General Exam|3738,3744|false|false|false|C0036412|Scleral Diseases|sclera
Event|Event|General Exam|3738,3744|false|false|false|||sclera
Procedure|Health Care Activity|General Exam|3738,3744|false|false|false|C2228481|examination of sclera|sclera
Event|Event|General Exam|3745,3754|false|false|false|||anicteric
Finding|Finding|General Exam|3745,3754|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3756,3759|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3756,3759|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3764,3769|false|false|false|||Clear
Finding|Idea or Concept|General Exam|3764,3769|false|false|false|C1550016|Remote control command - Clear|Clear
Anatomy|Body Location or Region|General Exam|3772,3776|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3772,3776|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3772,3776|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|3781,3784|true|false|false|||JVD
Finding|Finding|General Exam|3781,3784|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|General Exam|3789,3797|true|false|false|C0027530|Neck|cervical
Disorder|Disease or Syndrome|General Exam|3789,3813|true|false|false|C0235592|Cervical lymphadenopathy|cervical lymphadenopathy
Finding|Finding|General Exam|3789,3813|true|false|false|C4551446|Swollen lymph nodes in the neck|cervical lymphadenopathy
Disorder|Disease or Syndrome|General Exam|3798,3813|true|false|false|C0497156|Lymphadenopathy|lymphadenopathy
Event|Event|General Exam|3798,3813|true|false|false|||lymphadenopathy
Finding|Sign or Symptom|General Exam|3798,3813|true|false|false|C4282165|Swollen Lymph Node|lymphadenopathy
Anatomy|Body Part, Organ, or Organ Component|General Exam|3815,3822|true|false|false|C0040578;C4299086|Neck+Chest>Trachea;Trachea|trachea
Disorder|Disease or Syndrome|General Exam|3815,3822|true|false|false|C0040580;C0153953;C0154070|Benign neoplasm of trachea;Carcinoma in situ of trachea;Tracheal Diseases|trachea
Disorder|Neoplastic Process|General Exam|3815,3822|true|false|false|C0040580;C0153953;C0154070|Benign neoplasm of trachea;Carcinoma in situ of trachea;Tracheal Diseases|trachea
Event|Event|General Exam|3815,3822|true|false|false|||trachea
Finding|Finding|General Exam|3815,3822|true|false|false|C5848218|trachea findings|trachea
Procedure|Therapeutic or Preventive Procedure|General Exam|3815,3822|true|false|false|C0872391|Procedure on trachea|trachea
Anatomy|Cell Component|General Exam|3823,3830|true|false|false|C1660780|midline cell component|midline
Anatomy|Body Part, Organ, or Organ Component|General Exam|3833,3836|true|false|false|C0018787|Heart|COR
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3833,3836|true|false|false|C0056331|cordycepin|COR
Drug|Pharmacologic Substance|General Exam|3833,3836|true|false|false|C0056331|cordycepin|COR
Event|Activity|General Exam|3846,3850|true|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3846,3850|true|false|false|||rate
Finding|Idea or Concept|General Exam|3846,3850|true|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|3855,3861|true|false|false|||rhythm
Finding|Finding|General Exam|3855,3861|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3855,3861|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|3873,3879|true|false|false|||normal
Event|Event|General Exam|3886,3890|false|false|false|||PULM
Procedure|Health Care Activity|General Exam|3886,3890|false|false|false|C1315068|Pulmonary ventilator management|PULM
Finding|Finding|General Exam|3892,3915|false|false|false|C0238844|Decreased breath sounds|Decreased breath sounds
Finding|Body Substance|General Exam|3902,3908|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|General Exam|3902,3915|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Event|Event|General Exam|3909,3915|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3909,3915|false|false|false|C0037709||sounds
Event|Event|General Exam|3939,3944|false|false|false|||faint
Finding|Finding|General Exam|3939,3944|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Finding|Sign or Symptom|General Exam|3939,3944|false|false|false|C0039070;C4554554|Faint - appearance;Syncope|faint
Event|Event|General Exam|3956,3964|false|false|false|||crackles
Finding|Finding|General Exam|3956,3964|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Idea or Concept|General Exam|3967,3971|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Event|Event|General Exam|3972,3978|false|false|false|||effort
Finding|Organism Function|General Exam|3972,3978|false|false|false|C0015264|Exertion|effort
Anatomy|Body Location or Region|General Exam|3984,3987|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3984,3987|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|3984,3987|false|false|false|||ABD
Disorder|Disease or Syndrome|General Exam|3989,3993|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|3989,3993|false|false|false|||Soft
Event|Event|General Exam|3995,3997|true|false|false|||NT
Event|Event|General Exam|4011,4014|true|false|false|||HSM
Finding|Gene or Genome|General Exam|4011,4014|true|false|false|C1537594|LRRC4B gene|HSM
Disorder|Congenital Abnormality|General Exam|4016,4019|true|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|4016,4019|true|false|false|||EXT
Finding|Gene or Genome|General Exam|4016,4019|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Attribute|Clinical Attribute|General Exam|4039,4044|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|4039,4044|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|4039,4044|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|4039,4044|false|false|false|||alert
Finding|Finding|General Exam|4039,4044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|4039,4044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|4039,4044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|4046,4054|false|false|false|||oriented
Finding|Finding|General Exam|4046,4054|false|false|false|C1961028|Oriented to place|oriented
Finding|Finding|General Exam|4046,4064|false|false|false|C1961030|Oriented to person|oriented to person
Attribute|Clinical Attribute|General Exam|4058,4064|false|false|false|C5890614||person
Event|Event|General Exam|4058,4064|false|false|false|||person
Finding|Intellectual Product|General Exam|4058,4064|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|4066,4071|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|4066,4071|false|false|false|||place
Finding|Functional Concept|General Exam|4066,4071|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|4066,4071|false|false|false|C1533810||place
Finding|Finding|General Exam|4077,4081|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|General Exam|4077,4081|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|General Exam|4077,4081|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|General Exam|4104,4110|false|false|false|||intact
Finding|Finding|General Exam|4104,4110|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|4112,4117|false|false|false|||Moves
Anatomy|Body Part, Organ, or Organ Component|General Exam|4124,4135|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Anatomy|Body System|General Exam|4139,4143|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|4139,4143|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|4139,4143|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|General Exam|4139,4143|false|false|false|||SKIN
Finding|Body Substance|General Exam|4139,4143|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|4139,4143|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|General Exam|4148,4156|true|false|false|||jaundice
Finding|Finding|General Exam|4148,4156|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|General Exam|4148,4156|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|General Exam|4158,4166|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|4158,4166|true|false|false|C0010520|Cyanosis|cyanosis
Disorder|Disease or Syndrome|General Exam|4177,4187|true|false|false|C0011603|Dermatitis|dermatitis
Event|Event|General Exam|4177,4187|true|false|false|||dermatitis
Event|Event|General Exam|4192,4202|true|false|false|||ecchymoses
Finding|Pathologic Function|General Exam|4192,4202|true|false|false|C0013491|Ecchymosis|ecchymoses
Anatomy|Cell|General Exam|4247,4250|false|false|false|C0023516|Leukocytes|WBC
Event|Event|General Exam|4247,4250|false|false|false|||WBC
Anatomy|Cell|General Exam|4258,4261|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4258,4261|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4258,4261|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4269,4272|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|General Exam|4269,4272|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|General Exam|4269,4272|false|false|false|||HGB
Finding|Gene or Genome|General Exam|4269,4272|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|General Exam|4269,4272|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|General Exam|4278,4281|false|false|false|||HCT
Procedure|Laboratory Procedure|General Exam|4278,4281|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|General Exam|4278,4281|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|General Exam|4289,4292|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4289,4292|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4289,4292|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4289,4292|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4289,4292|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4297,4300|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4297,4300|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4297,4300|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4297,4300|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4297,4300|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4297,4300|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4307,4311|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|4317,4320|false|false|false|||RDW
Event|Event|General Exam|4341,4344|false|false|false|||PLT
Procedure|Laboratory Procedure|General Exam|4341,4344|false|false|false|C0201617|Primed lymphocyte test|PLT
Event|Event|General Exam|4369,4374|false|false|false|||NEUTS
Finding|Body Substance|General Exam|4388,4394|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|General Exam|4398,4403|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|General Exam|4398,4403|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|General Exam|4398,4403|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|General Exam|4406,4409|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|General Exam|4406,4409|false|false|false|||EOS
Finding|Gene or Genome|General Exam|4406,4409|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Finding|Body Substance|General Exam|4540,4548|false|false|false|C0039409|Tears (substance)|TEARDROP
Disorder|Neoplastic Process|General Exam|4582,4585|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4582,4585|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4582,4585|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|General Exam|4609,4616|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|4609,4616|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|4609,4616|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|4609,4616|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|4609,4616|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|4609,4616|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|General Exam|4622,4626|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|General Exam|4622,4626|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|General Exam|4622,4626|false|false|false|C0041942|urea|UREA
Event|Event|General Exam|4622,4626|false|false|false|||UREA
Procedure|Laboratory Procedure|General Exam|4622,4626|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|General Exam|4644,4650|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|General Exam|4644,4650|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|General Exam|4644,4650|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|General Exam|4644,4650|false|false|false|||SODIUM
Finding|Physiologic Function|General Exam|4644,4650|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|General Exam|4644,4650|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|General Exam|4656,4665|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4656,4665|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|General Exam|4656,4665|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|General Exam|4656,4665|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|General Exam|4656,4665|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|General Exam|4656,4665|false|false|false|||POTASSIUM
Finding|Physiologic Function|General Exam|4656,4665|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|General Exam|4656,4665|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|General Exam|4670,4678|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|General Exam|4670,4678|false|false|false|||CHLORIDE
Finding|Physiologic Function|General Exam|4670,4678|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|General Exam|4670,4678|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|General Exam|4688,4691|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|General Exam|4688,4691|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|General Exam|4688,4691|false|false|false|||CO2
Finding|Finding|General Exam|4688,4691|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|General Exam|4688,4691|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|General Exam|4695,4700|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|General Exam|4695,4704|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|General Exam|4695,4704|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|General Exam|4695,4704|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|General Exam|4701,4704|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|General Exam|4701,4704|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|General Exam|4701,4704|false|false|false|||GAP
Finding|Gene or Genome|General Exam|4701,4704|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Organic Chemical|General Exam|4722,4729|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Drug|Pharmacologic Substance|General Exam|4722,4729|false|false|false|C0022924;C0376261|Lactates;lactate|LACTATE
Event|Event|General Exam|4722,4729|false|false|false|||LACTATE
Procedure|Laboratory Procedure|General Exam|4722,4729|false|false|false|C0202115|Lactic acid measurement|LACTATE
Finding|Body Substance|General Exam|4775,4780|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4775,4780|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4775,4780|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|4775,4787|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|General Exam|4782,4787|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4782,4787|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|General Exam|4782,4787|false|false|false|||COLOR
Drug|Organic Chemical|General Exam|4788,4793|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|General Exam|4801,4806|false|false|false|||Clear
Finding|Idea or Concept|General Exam|4801,4806|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|4826,4831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|4826,4831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|4826,4831|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|4826,4838|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|General Exam|4833,4838|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4833,4838|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4833,4838|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4839,4842|false|false|false|||NEG
Finding|Finding|General Exam|4839,4842|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|4843,4850|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|General Exam|4843,4850|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|General Exam|4843,4850|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Finding|Finding|General Exam|4851,4854|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|4855,4862|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|General Exam|4855,4862|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|General Exam|4855,4862|false|false|false|||PROTEIN
Finding|Conceptual Entity|General Exam|4855,4862|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|General Exam|4855,4862|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|General Exam|4863,4866|false|false|false|||NEG
Finding|Finding|General Exam|4863,4866|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|4868,4875|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|General Exam|4868,4875|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|General Exam|4868,4875|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|General Exam|4868,4875|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|General Exam|4868,4875|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|General Exam|4868,4875|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|General Exam|4876,4879|false|false|false|||NEG
Finding|Finding|General Exam|4876,4879|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|4880,4886|false|false|false|C0022634|Ketones|KETONE
Event|Event|General Exam|4887,4890|false|false|false|||NEG
Finding|Finding|General Exam|4887,4890|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|4891,4900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|General Exam|4891,4900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|General Exam|4891,4900|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|General Exam|4891,4900|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|General Exam|4901,4904|false|false|false|||NEG
Finding|Finding|General Exam|4901,4904|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|4915,4918|false|false|false|||NEG
Finding|Finding|General Exam|4915,4918|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|4932,4935|false|false|false|||NEG
Finding|Finding|General Exam|4932,4935|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|4938,4943|false|false|false|||Micro
Finding|Conceptual Entity|General Exam|4938,4943|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Finding|Intellectual Product|General Exam|4938,4943|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|Micro
Procedure|Laboratory Procedure|General Exam|4938,4943|false|false|false|C0085672|Microbiology procedure|Micro
Procedure|Laboratory Procedure|General Exam|4945,4971|false|false|false|C2721555|Legionella urinary antigen|Legionella Urinary Antigen
Anatomy|Body Part, Organ, or Organ Component|General Exam|4956,4963|false|false|false|C0042027|Urinary tract|Urinary
Drug|Immunologic Factor|General Exam|4964,4971|false|false|false|C0003320|Antigens|Antigen
Event|Event|General Exam|4964,4971|false|false|false|||Antigen
Finding|Idea or Concept|General Exam|4974,4979|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|4992,5000|false|false|false|||NEGATIVE
Finding|Classification|General Exam|4992,5000|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|General Exam|4992,5000|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|General Exam|4992,5000|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Finding|General Exam|4992,5004|false|false|false|C0205160|Negative|NEGATIVE FOR
Finding|Intellectual Product|General Exam|5016,5025|true|false|false|C0449543|Serogroup|SEROGROUP
Drug|Immunologic Factor|General Exam|5028,5035|true|false|false|C0003320|Antigens|ANTIGEN
Event|Event|General Exam|5028,5035|true|false|false|||ANTIGEN
Finding|Body Substance|General Exam|5038,5043|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|General Exam|5038,5043|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|General Exam|5038,5043|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Body Substance|General Exam|5050,5055|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|5050,5055|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|5050,5055|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|General Exam|5050,5063|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|General Exam|5056,5063|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|General Exam|5056,5063|false|false|false|||CULTURE
Finding|Functional Concept|General Exam|5056,5063|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|5056,5063|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|5056,5063|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|General Exam|5065,5070|false|false|false|||Final
Finding|Idea or Concept|General Exam|5065,5070|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|General Exam|5082,5088|true|false|false|||GROWTH
Finding|Finding|General Exam|5082,5088|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|5082,5088|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|5082,5088|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|5082,5088|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|5082,5088|true|false|false|C2911660|Growth action|GROWTH
Disorder|Disease or Syndrome|General Exam|5091,5096|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|General Exam|5091,5096|false|false|false|||Blood
Finding|Body Substance|General Exam|5091,5096|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|5108,5115|false|false|false|||Studies
Procedure|Research Activity|General Exam|5108,5115|false|false|false|C0947630|Scientific Study|Studies
Event|Event|General Exam|5116,5123|false|false|false|||Imaging
Finding|Finding|General Exam|5116,5123|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|General Exam|5116,5123|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|General Exam|5127,5130|false|false|false|||EKG
Finding|Intellectual Product|General Exam|5127,5130|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|5127,5130|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|General Exam|5136,5141|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|General Exam|5136,5141|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|General Exam|5136,5141|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|General Exam|5136,5141|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|General Exam|5136,5148|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|General Exam|5142,5148|false|false|false|||rhythm
Finding|Finding|General Exam|5142,5148|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|5142,5148|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|5155,5158|false|false|false|||bpm
Procedure|Therapeutic or Preventive Procedure|General Exam|5155,5158|false|false|false|C1706504|Bilateral Prophylactic Mastectomy|bpm
Anatomy|Body Part, Organ, or Organ Component|General Exam|5167,5171|false|false|false|C0004457|Axis vertebra|axis
Disorder|Injury or Poisoning|General Exam|5167,5171|false|false|false|C0349013|Fracture of second cervical vertebra|axis
Event|Event|General Exam|5180,5189|false|false|false|||intervals
Event|Event|General Exam|5191,5195|false|false|false|||poor
Finding|Intellectual Product|General Exam|5191,5195|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Gene or Genome|General Exam|5199,5203|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|General Exam|5199,5203|false|false|false|C0678544||wave
Event|Event|General Exam|5204,5214|false|false|false|||progresion
Disorder|Mental or Behavioral Dysfunction|General Exam|5219,5230|false|false|false|C0011570|Mental Depression|depressions
Event|Event|General Exam|5219,5230|false|false|false|||depressions
Event|Event|General Exam|5243,5246|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5243,5246|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|General Exam|5252,5258|false|false|false|||SINGLE
Finding|Finding|General Exam|5252,5258|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|SINGLE
Event|Event|General Exam|5262,5266|false|false|false|||VIEW
Anatomy|Body Location or Region|General Exam|5274,5279|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|General Exam|5274,5279|false|false|false|C0741025|Chest problem|CHEST
Finding|Body Substance|General Exam|5281,5288|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|5281,5288|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|5281,5288|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|General Exam|5292,5298|false|false|false|C5889824||status
Event|Event|General Exam|5292,5298|false|false|false|||status
Finding|Idea or Concept|General Exam|5292,5298|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|5312,5322|false|false|false|||sternotomy
Procedure|Therapeutic or Preventive Procedure|General Exam|5312,5322|false|false|false|C0185792|Sternotomy (procedure)|sternotomy
Anatomy|Body Part, Organ, or Organ Component|General Exam|5329,5336|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|General Exam|5329,5336|false|false|false|C1314974|Cardiac attachment|cardiac
Anatomy|Body Location or Region|General Exam|5338,5349|false|false|false|C0025066|Mediastinum|mediastinal
Event|Event|General Exam|5360,5368|false|false|false|||contours
Event|Event|General Exam|5373,5382|false|false|false|||unchanged
Finding|Finding|General Exam|5373,5382|false|false|false|C0442739||unchanged
Event|Event|General Exam|5391,5400|false|false|false|||continues
Event|Event|General Exam|5407,5418|false|false|false|||progression
Finding|Functional Concept|General Exam|5407,5418|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|General Exam|5407,5418|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|General Exam|5422,5429|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5422,5429|false|false|false|||disease
Finding|Finding|General Exam|5435,5444|false|false|true|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|General Exam|5435,5444|false|false|true|C0442805;C5236002|Increase;Increased (finding)|increased
Event|Event|General Exam|5445,5451|false|false|false|||extent
Event|Event|General Exam|5470,5477|false|false|false|||opacity
Finding|Finding|General Exam|5470,5477|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|General Exam|5470,5477|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Functional Concept|General Exam|5489,5494|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5489,5499|false|false|false|C0225706|Right lung|right lung
Anatomy|Body Location or Region|General Exam|5489,5504|false|false|false|C0225708|Structure of base of right lung|right lung base
Anatomy|Body Location or Region|General Exam|5495,5499|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|5495,5499|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|5495,5499|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|5495,5499|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|5495,5504|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|General Exam|5500,5504|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|5500,5504|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|5500,5504|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|5500,5504|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|5500,5504|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|5500,5504|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Sign or Symptom|General Exam|5506,5509|false|false|false|C0231218|Malaise|Ill
Event|Event|General Exam|5510,5517|false|false|false|||defined
Event|Event|General Exam|5519,5528|false|false|false|||opacities
Finding|Finding|General Exam|5519,5528|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|General Exam|5519,5528|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Anatomy|Body Part, Organ, or Organ Component|General Exam|5540,5547|false|false|false|C0225740;C0228475;C1561517|Lingula;Lingula of cerebellum;Lingula of left lung|lingula
Finding|Functional Concept|General Exam|5552,5556|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5552,5567|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|General Exam|5557,5562|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5557,5562|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5557,5567|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|General Exam|5563,5567|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|General Exam|5563,5567|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|General Exam|5572,5579|false|false|false|||similar
Finding|Functional Concept|General Exam|5597,5602|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Tissue|General Exam|5603,5610|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|5603,5610|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Body Substance|General Exam|5603,5619|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Finding|General Exam|5603,5619|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Finding|Pathologic Function|General Exam|5603,5619|false|false|false|C0032227;C1253943;C2073625|Pleural effusion (disorder);Pleural effusion fluid|pleural effusion
Event|Event|General Exam|5611,5619|false|false|false|||effusion
Finding|Body Substance|General Exam|5611,5619|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|5611,5619|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|5611,5619|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|General Exam|5623,5630|false|false|false|||present
Finding|Finding|General Exam|5623,5630|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|5623,5630|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Disease or Syndrome|General Exam|5645,5657|true|false|false|C0032326|Pneumothorax|pneumothorax
Event|Event|General Exam|5645,5657|true|false|false|||pneumothorax
Disorder|Anatomical Abnormality|General Exam|5668,5682|false|false|false|C0020449|Hyperdistention|hyperinflation
Event|Event|General Exam|5668,5682|false|false|false|||hyperinflation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5690,5695|false|false|false|C0024109|Lung|lungs
Event|Event|General Exam|5698,5708|false|false|false|||IMPRESSION
Finding|Intellectual Product|General Exam|5698,5708|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|5698,5708|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|General Exam|5710,5718|false|false|false|||Evidence
Finding|Idea or Concept|General Exam|5710,5718|false|false|false|C3887511|Evidence|Evidence
Finding|Functional Concept|General Exam|5710,5721|false|false|false|C0332120|Evidence of (contextual qualifier)|Evidence of
Disorder|Disease or Syndrome|General Exam|5722,5729|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|5722,5729|false|false|false|||disease
Finding|Pathologic Function|General Exam|5722,5741|false|false|false|C0242656|Disease Progression|disease progression
Event|Event|General Exam|5730,5741|false|false|false|||progression
Finding|Functional Concept|General Exam|5730,5741|true|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|General Exam|5730,5741|true|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Attribute|Clinical Attribute|General Exam|5746,5753|false|false|false|C0881943||CT Head
Procedure|Diagnostic Procedure|General Exam|5746,5753|false|false|false|C0202691|CAT scan of head|CT Head
Anatomy|Body Location or Region|General Exam|5749,5753|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|General Exam|5749,5753|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|General Exam|5749,5753|false|false|false|C0362076|Problems with head|Head
Event|Event|General Exam|5749,5753|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|General Exam|5749,5753|false|false|false|C0876917|Procedure on head|Head
Event|Event|Findings|5781,5789|true|false|false|||evidence
Finding|Idea or Concept|Findings|5781,5789|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|5781,5792|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|Findings|5793,5798|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Findings|5793,5809|true|false|false|C0333276|Acute hemorrhage|acute hemorrhage
Event|Event|Findings|5799,5809|true|false|false|||hemorrhage
Finding|Pathologic Function|Findings|5799,5809|true|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|Findings|5811,5816|true|false|false|C1717255||edema
Event|Event|Findings|5811,5816|true|false|false|||edema
Finding|Pathologic Function|Findings|5811,5816|true|false|false|C0013604|Edema|edema
Event|Event|Findings|5818,5822|false|false|false|||mass
Finding|Finding|Findings|5818,5822|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|5818,5822|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|5818,5822|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Findings|5824,5830|false|false|false|||effect
Event|Event|Findings|5842,5852|false|false|false|||infarction
Finding|Pathologic Function|Findings|5842,5852|false|false|false|C0021308|Infarction|infarction
Event|Governmental or Regulatory Activity|Findings|5857,5861|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Disease or Syndrome|Findings|5865,5881|false|false|false|C0014068|Encephalomalacia|encephalomalacia
Event|Event|Findings|5865,5881|false|false|false|||encephalomalacia
Finding|Functional Concept|Findings|5889,5893|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Findings|5895,5907|false|false|false|C0016733|frontal lobe|frontal lobe
Disorder|Neoplastic Process|Findings|5895,5907|false|false|false|C0153635|malignant neoplasm of frontal lobe|frontal lobe
Anatomy|Body Part, Organ, or Organ Component|Findings|5903,5907|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Findings|5903,5907|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Findings|5910,5920|false|false|false|||compatible
Finding|Idea or Concept|Findings|5910,5920|false|false|false|C0332290|Consistent with|compatible
Finding|Idea or Concept|Findings|5910,5925|false|false|false|C0332290|Consistent with|compatible with
Event|Event|Findings|5926,5933|false|false|false|||chronic
Finding|Intellectual Product|Findings|5926,5933|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Findings|5926,5933|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Event|Event|Findings|5934,5941|false|false|false|||infarct
Finding|Pathologic Function|Findings|5934,5941|false|false|false|C0021308|Infarction|infarct
Event|Event|Findings|5945,5954|false|false|false|||unchanged
Finding|Finding|Findings|5945,5954|false|false|false|C0442739||unchanged
Event|Event|Findings|5956,5966|false|false|false|||Prominence
Anatomy|Body Part, Organ, or Organ Component|Findings|5975,5985|false|false|false|C0018827|Heart Ventricle|ventricles
Event|Event|Findings|5997,6005|false|false|false|||reflects
Event|Event|Findings|6018,6025|false|false|false|||atrophy
Finding|Pathologic Function|Findings|6018,6025|false|false|false|C0333641|Atrophic|atrophy
Event|Event|Findings|6064,6070|false|false|false|||spaces
Anatomy|Body Location or Region|Findings|6101,6112|false|false|false|C0815275|Subcortical|subcortical
Anatomy|Tissue|Findings|6114,6126|false|false|false|C0682708|White matter|white matter
Finding|Finding|Findings|6139,6145|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Findings|6139,6145|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Findings|6146,6153|false|false|false|||reflect
Event|Event|Findings|6154,6161|false|false|false|||sequela
Finding|Pathologic Function|Findings|6154,6161|false|true|false|C0543419|Sequela of disorder|sequela
Event|Event|Findings|6165,6172|false|false|false|||chronic
Finding|Intellectual Product|Findings|6165,6172|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Findings|6165,6172|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Location or Region|Findings|6180,6186|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Findings|6180,6186|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Finding|Functional Concept|Findings|6187,6195|false|false|false|C0475224|Ischemic|ischemic
Disorder|Disease or Syndrome|Findings|6196,6203|false|false|false|C0012634|Disease|disease
Event|Event|Findings|6196,6203|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|Findings|6219,6226|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Anatomy|Tissue|Findings|6219,6226|true|false|false|C0262950;C4520924|Bone Tissue, Human;Skeletal bone|osseous
Event|Event|Findings|6227,6233|true|false|false|||lesion
Finding|Finding|Findings|6227,6233|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Findings|6227,6233|true|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|Findings|6237,6241|true|false|false|||seen
Event|Event|Findings|6254,6268|false|false|false|||calcifications
Finding|Finding|Findings|6254,6268|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|Findings|6254,6268|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|Findings|6286,6293|false|false|false|C0007272|Carotid Arteries|carotid
Event|Event|Findings|6294,6301|false|false|false|||siphons
Event|Event|Findings|6308,6318|false|false|false|||visualized
Anatomy|Body Space or Junction|Findings|6319,6336|false|false|false|C0030471|Nasal sinus|paranasal sinuses
Anatomy|Body Space or Junction|Findings|6329,6336|false|false|false|C0030471;C4071871|Head>Sinuses;Nasal sinus|sinuses
Disorder|Anatomical Abnormality|Findings|6329,6336|false|false|false|C0016169|pathologic fistula|sinuses
Event|Event|Findings|6329,6336|false|false|false|||sinuses
Event|Event|Findings|6349,6361|false|false|false|||unremarkable
Event|Event|Findings|6364,6374|false|false|false|||IMPRESSION
Finding|Intellectual Product|Findings|6364,6374|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|6364,6374|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|Findings|6379,6387|true|false|false|||evidence
Finding|Idea or Concept|Findings|6379,6387|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|6379,6390|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|Findings|6391,6396|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Findings|6397,6409|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Findings|6397,6409|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|Findings|6410,6417|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Findings|6410,6417|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Findings|6410,6417|true|false|false|||process
Finding|Functional Concept|Findings|6410,6417|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Findings|6410,6417|true|false|false|C1522240|Process|process
Event|Event|Findings|6421,6425|true|false|false|||mass
Finding|Finding|Findings|6421,6425|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Findings|6421,6425|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Findings|6421,6425|true|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|Findings|6448,6458|false|false|false|||IMPRESSION
Finding|Intellectual Product|Findings|6448,6458|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Findings|6448,6458|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|Findings|6463,6471|true|false|false|||evidence
Finding|Idea or Concept|Findings|6463,6471|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Findings|6463,6474|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Location or Region|Findings|6475,6478|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Findings|6475,6478|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Findings|6475,6478|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Findings|6475,6478|true|false|false|||DVT
Attribute|Clinical Attribute|Findings|6483,6491|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|Findings|6483,6491|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|Findings|6486,6491|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Findings|6486,6491|false|false|false|C0741025|Chest problem|chest
Finding|Intellectual Product|Impression|6513,6521|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Event|Event|Impression|6522,6531|false|false|false|||worsening
Finding|Idea or Concept|Impression|6522,6531|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|Impression|6560,6565|false|false|false|C2676739|Chromosome 2q32-Q33 Deletion Syndrome|glass
Drug|Hazardous or Poisonous Substance|Impression|6560,6565|false|false|false|C0025611|methamphetamine|glass
Drug|Organic Chemical|Impression|6560,6565|false|false|false|C0025611|methamphetamine|glass
Drug|Pharmacologic Substance|Impression|6560,6565|false|false|false|C0025611|methamphetamine|glass
Event|Event|Impression|6560,6565|false|false|false|||glass
Event|Event|Impression|6567,6576|false|false|false|||opacities
Finding|Finding|Impression|6567,6576|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Finding|Pathologic Function|Impression|6567,6576|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacities
Anatomy|Body Part, Organ, or Organ Component|Impression|6579,6590|false|false|false|C0006270|Bronchioles|bronchiolar
Event|Event|Impression|6591,6598|false|false|false|||nodules
Disorder|Disease or Syndrome|Impression|6609,6622|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Impression|6609,6622|false|false|false|||consolidation
Anatomy|Body Part, Organ, or Organ Component|Impression|6634,6641|false|false|false|C0225740;C0228475;C1561517|Lingula;Lingula of cerebellum;Lingula of left lung|lingula
Finding|Functional Concept|Impression|6647,6652|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Intellectual Product|Impression|6654,6660|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|Impression|6654,6665|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|6661,6665|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|6661,6665|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Event|Event|Impression|6673,6679|false|false|false|||review
Finding|Idea or Concept|Impression|6673,6679|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|Impression|6673,6679|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|Impression|6673,6682|false|false|false|C0699752|Review of|review of
Anatomy|Body Location or Region|Impression|6705,6710|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|6705,6710|false|false|false|C0741025|Chest problem|chest
Drug|Pharmacologic Substance|Impression|6711,6717|false|false|false|C0885876|X-rays, Homeopathic Preparations|x-rays
Event|Event|Impression|6711,6717|false|false|false|||x-rays
Phenomenon|Natural Phenomenon or Process|Impression|6711,6717|false|false|false|C0043309|Roentgen Rays|x-rays
Procedure|Diagnostic Procedure|Impression|6711,6717|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|x-rays
Disorder|Disease or Syndrome|Impression|6723,6726|false|false|false|C0007286|Carpal Tunnel Syndrome|CTs
Drug|Amino Acid, Peptide, or Protein|Impression|6723,6726|false|false|false|C3813556|Cancer/Testis Antigen|CTs
Event|Event|Impression|6723,6726|false|false|false|||CTs
Finding|Gene or Genome|Impression|6723,6726|false|false|false|C1421224;C2699876|TTR gene;TTR wt Allele|CTs
Procedure|Molecular Biology Research Technique|Impression|6723,6726|false|false|false|C5891069|Concatenated Tag Sequencing|CTs
Attribute|Clinical Attribute|Impression|6734,6742|false|false|false|C2926606||findings
Event|Event|Impression|6734,6742|false|false|false|||findings
Finding|Functional Concept|Impression|6734,6742|false|false|false|C2607943|findings aspects|findings
Event|Event|Impression|6754,6763|false|false|false|||explained
Event|Event|Impression|6767,6776|false|false|false|||worsening
Finding|Idea or Concept|Impression|6767,6776|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Neoplastic Process|Impression|6778,6804|true|false|false|C0007120|Bronchioloalveolar Adenocarcinoma|bronchioalveolar carcinoma
Disorder|Neoplastic Process|Impression|6795,6804|true|false|false|C0007097|Carcinoma|carcinoma
Event|Event|Impression|6795,6804|true|false|false|||carcinoma
Disorder|Anatomical Abnormality|Impression|6816,6823|true|false|false|C1689985|Absence (morphologic abnormality)|absence
Event|Event|Impression|6816,6823|true|false|false|||absence
Finding|Functional Concept|Impression|6816,6823|true|false|false|C0332197|Absent|absence
Finding|Functional Concept|Impression|6816,6826|true|false|false|C0332197|Absent|absence of
Event|Event|Impression|6831,6837|true|false|false|||change
Finding|Functional Concept|Impression|6831,6837|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Impression|6831,6837|true|false|false|C4319952|Change - procedure|change
Event|Event|Impression|6855,6862|true|false|false|||suggest
Disorder|Disease or Syndrome|Impression|6863,6872|true|true|false|C0032285|Pneumonia|pneumonia
Event|Event|Impression|6863,6872|true|false|false|||pneumonia
Disorder|Disease or Syndrome|Impression|6884,6893|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Impression|6884,6893|false|false|false|||pneumonia
Event|Event|Impression|6904,6911|false|false|false|||present
Finding|Finding|Impression|6904,6911|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Impression|6904,6911|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|Impression|6916,6928|false|false|false|||unrecognized
Event|Event|Impression|6934,6943|false|false|false|||treatment
Finding|Conceptual Entity|Impression|6934,6943|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Impression|6934,6943|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Impression|6934,6943|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Impression|6934,6943|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Impression|6954,6958|false|false|false|||made
Drug|Pharmacologic Substance|Impression|6967,6972|false|false|false|C1874451|Basis|basis
Event|Event|Impression|6967,6972|false|false|false|||basis
Finding|Functional Concept|Impression|6967,6972|false|false|false|C1527178|Basis - conceptual entity|basis
Finding|Intellectual Product|Impression|6976,6984|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Finding|Sign or Symptom|Impression|6976,6993|false|false|false|C0037088|Signs and Symptoms|clinical findings
Attribute|Clinical Attribute|Impression|6985,6993|false|false|false|C2926606||findings
Event|Event|Impression|6985,6993|false|false|false|||findings
Finding|Functional Concept|Impression|6985,6993|false|false|false|C2607943|findings aspects|findings
Event|Event|Impression|6999,7005|false|false|false|||Stable
Finding|Intellectual Product|Impression|6999,7005|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Intellectual Product|Impression|7006,7010|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|Impression|7011,7023|false|false|false|||cardiomegaly
Finding|Finding|Impression|7011,7023|false|false|false|C0018800|Cardiomegaly|cardiomegaly
Finding|Finding|Impression|7029,7037|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Impression|7029,7037|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Disorder|Disease or Syndrome|Impression|7038,7047|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|Impression|7038,7047|false|false|false|||emphysema
Finding|Pathologic Function|Impression|7038,7047|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Disorder|Disease or Syndrome|Impression|7053,7067|true|false|false|C0008350|Cholelithiasis|Cholelithiasis
Event|Event|Impression|7053,7067|true|false|false|||Cholelithiasis
Event|Event|Impression|7076,7084|true|false|false|||evidence
Finding|Idea or Concept|Impression|7076,7084|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|7076,7087|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Impression|7088,7101|true|false|false|C0008325|Cholecystitis|cholecystitis
Event|Event|Impression|7088,7101|true|false|false|||cholecystitis
Disorder|Neoplastic Process|Hospital Course|7146,7151|false|false|false|C0007131||NSCLC
Attribute|Clinical Attribute|Hospital Course|7152,7157|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|7152,7160|false|false|false|C0441772|Stage level 4|stage IV
Event|Event|Hospital Course|7161,7169|false|false|false|||presents
Event|Event|Hospital Course|7175,7182|false|false|false|||hypoxia
Finding|Finding|Hospital Course|7175,7182|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|Hospital Course|7175,7182|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|Hospital Course|7189,7196|false|false|false|||Hypoxia
Finding|Finding|Hospital Course|7189,7196|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Finding|Pathologic Function|Hospital Course|7189,7196|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|Hypoxia
Event|Event|Hospital Course|7201,7210|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7201,7210|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|7211,7218|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7211,7218|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7211,7218|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|7230,7240|false|false|false|||complaints
Finding|Finding|Hospital Course|7230,7240|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Functional Concept|Hospital Course|7245,7256|false|false|false|C0205329|Progressive|progressive
Event|Event|Hospital Course|7257,7266|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|7257,7276|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|7257,7276|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|7270,7276|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|7296,7301|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|7296,7301|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|7296,7301|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|7296,7301|false|false|false|C0010200|Coughing|cough
Finding|Idea or Concept|Hospital Course|7307,7311|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7307,7311|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7307,7311|true|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|7307,7318|true|false|false|C0421203|Home oxygen supply|home oxygen
Drug|Biologically Active Substance|Hospital Course|7312,7318|true|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|7312,7318|true|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|7312,7318|true|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|7312,7318|true|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7312,7318|true|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|7319,7330|true|false|false|||requirement
Finding|Functional Concept|Hospital Course|7319,7330|true|false|false|C1514873|Requirement|requirement
Drug|Biomedical or Dental Material|Hospital Course|7334,7342|true|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|7334,7342|true|false|false|||baseline
Finding|Idea or Concept|Hospital Course|7334,7342|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|7347,7356|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|7347,7356|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|7365,7371|false|false|false|||placed
Event|Event|Hospital Course|7376,7379|false|false|false|||NRB
Event|Event|Hospital Course|7384,7393|false|false|false|||treatment
Finding|Conceptual Entity|Hospital Course|7384,7393|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|7384,7393|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|7384,7393|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7384,7393|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Hospital Course|7400,7411|false|false|false|||saturations
Phenomenon|Natural Phenomenon or Process|Hospital Course|7400,7411|false|false|false|C0522534|Saturated|saturations
Event|Event|Hospital Course|7419,7430|false|false|false|||saturations
Phenomenon|Natural Phenomenon or Process|Hospital Course|7419,7430|false|false|false|C0522534|Saturated|saturations
Procedure|Health Care Activity|Hospital Course|7445,7454|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Hospital Course|7455,7458|true|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|7455,7458|true|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|Hospital Course|7476,7486|true|false|false|||infiltrate
Finding|Functional Concept|Hospital Course|7476,7486|true|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Hospital Course|7476,7486|true|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Hospital Course|7476,7486|true|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|Hospital Course|7495,7502|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|7495,7502|false|false|false|C2699424|Concern|concern
Event|Event|Hospital Course|7508,7519|false|false|false|||progression
Finding|Functional Concept|Hospital Course|7508,7519|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|7508,7519|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Anatomy|Body Location or Region|Hospital Course|7533,7537|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7533,7537|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|7533,7537|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|7533,7537|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Hospital Course|7533,7545|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Hospital Course|7538,7545|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|7538,7545|false|false|false|||disease
Finding|Mental Process|Hospital Course|7550,7557|false|false|false|C0542559|contextual factors|setting
Anatomy|Cell|Hospital Course|7571,7574|false|false|false|C0023516|Leukocytes|WBC
Event|Event|Hospital Course|7576,7583|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|7576,7583|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|7588,7598|false|false|false|C0009450|Communicable Diseases|infectious
Event|Event|Hospital Course|7588,7598|false|false|false|||infectious
Finding|Pathologic Function|Hospital Course|7588,7606|false|false|false|C0745283|INFECTIOUS PROCESS|infectious process
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7599,7606|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|7599,7606|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|Hospital Course|7599,7606|false|false|false|||process
Finding|Functional Concept|Hospital Course|7599,7606|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|7599,7606|false|false|false|C1522240|Process|process
Event|Event|Hospital Course|7624,7631|false|false|false|||treated
Drug|Antibiotic|Hospital Course|7637,7649|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|7637,7649|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|7637,7649|false|false|false|||levofloxacin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7654,7664|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|Hospital Course|7654,7664|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|Hospital Course|7654,7664|false|false|false|||vancomycin
Procedure|Laboratory Procedure|Hospital Course|7654,7664|false|false|false|C0489941|Vancomycin measurement|vancomycin
Event|Event|Hospital Course|7693,7704|false|false|false|||monotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7693,7704|false|false|false|C4763675|Single Agent Therapy|monotherapy
Drug|Antibiotic|Hospital Course|7710,7722|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|7710,7722|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|7710,7722|false|false|false|||levofloxacin
Drug|Antibiotic|Hospital Course|7734,7745|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|7734,7745|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|7734,7745|false|false|false|||ceftriaxone
Event|Event|Hospital Course|7757,7762|false|false|false|||added
Event|Event|Hospital Course|7771,7774|false|false|false|||CXR
Procedure|Diagnostic Procedure|Hospital Course|7771,7774|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Finding|Hospital Course|7795,7798|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|7795,7798|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Functional Concept|Hospital Course|7799,7803|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Hospital Course|7804,7809|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|7804,7809|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7811,7815|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|7811,7815|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Disorder|Disease or Syndrome|Hospital Course|7816,7829|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|Hospital Course|7816,7829|false|false|false|||consolidation
Finding|Functional Concept|Hospital Course|7831,7841|false|false|false|C1524062|Additional|Additional
Finding|Finding|Hospital Course|7842,7849|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|Hospital Course|7842,7849|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|Hospital Course|7850,7854|false|false|false|||work
Event|Occupational Activity|Hospital Course|7850,7854|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|7850,7857|false|false|false|C0750430|Work-up|work-up
Finding|Classification|Hospital Course|7871,7879|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7871,7879|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7871,7879|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|Hospital Course|7880,7890|true|false|false|C0005516|Biological Markers|biomarkers
Event|Event|Hospital Course|7880,7890|false|false|false|||biomarkers
Finding|Classification|Hospital Course|7892,7900|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7892,7900|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7892,7900|false|false|false|C5237010|Expression Negative|negative
Event|Event|Hospital Course|7908,7914|false|false|false|||unable
Finding|Finding|Hospital Course|7908,7914|false|false|false|C1299582|Unable|unable
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7926,7929|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|7926,7929|false|false|false|||CTA
Finding|Gene or Genome|Hospital Course|7926,7929|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|7926,7929|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|Hospital Course|7930,7933|false|false|false|||due
Finding|Functional Concept|Hospital Course|7930,7933|false|false|false|C0678226;C3146286|Due;Due to|due
Finding|Idea or Concept|Hospital Course|7930,7933|false|false|false|C0678226;C3146286|Due;Due to|due
Event|Event|Hospital Course|7938,7945|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|7938,7945|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|7938,7945|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|7938,7960|false|false|false|C1561643|Chronic Kidney Diseases|chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7946,7952|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|7946,7952|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|7946,7952|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|7946,7952|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7946,7952|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|7946,7960|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|7953,7960|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|7953,7960|false|false|false|||disease
Drug|Biologically Active Substance|Hospital Course|7965,7975|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|7965,7975|false|false|false|C0010294|creatinine|creatinine
Event|Event|Hospital Course|7965,7975|false|false|false|||creatinine
Finding|Physiologic Function|Hospital Course|7965,7975|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|7965,7975|false|false|false|C0201975|Creatinine measurement|creatinine
Finding|Body Substance|Hospital Course|7981,7988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7981,7988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7981,7988|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|7993,7997|false|false|false|||able
Finding|Finding|Hospital Course|7993,7997|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|8005,8011|false|false|false|||weaned
Drug|Inorganic Chemical|Hospital Course|8020,8028|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|Hospital Course|8025,8028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|8025,8028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|8025,8028|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|Hospital Course|8025,8028|false|false|false|||air
Finding|Finding|Hospital Course|8025,8028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|8025,8028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|8025,8028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8036,8039|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|8036,8039|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|Hospital Course|8036,8039|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|8036,8039|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Event|Event|Hospital Course|8052,8056|false|false|false|||stay
Event|Event|Hospital Course|8067,8078|false|false|false|||transferred
Finding|Functional Concept|Hospital Course|8086,8093|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|8086,8093|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|8086,8093|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|8086,8093|false|false|false|C0199168|Medical service|medical
Anatomy|Anatomical Structure|Hospital Course|8094,8099|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|8119,8131|false|false|false|||demonstrated
Finding|Sign or Symptom|Hospital Course|8132,8142|false|false|false|C0239313|exercise induced|exertional
Event|Event|Hospital Course|8143,8150|false|false|false|||hypoxia
Finding|Finding|Hospital Course|8143,8150|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|Hospital Course|8143,8150|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Finding|Hospital Course|8152,8159|false|false|false|C3888388|Usually|usually
Finding|Finding|Hospital Course|8152,8172|false|false|false|C1866557|Usually asymptomatic|usually asymptomatic
Event|Event|Hospital Course|8160,8172|false|false|false|||asymptomatic
Finding|Finding|Hospital Course|8160,8172|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Idea or Concept|Hospital Course|8174,8178|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8174,8178|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8174,8178|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|8187,8195|false|false|false|||arranged
Disorder|Disease or Syndrome|Hospital Course|8218,8227|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|8218,8227|false|false|false|||pneumonia
Disorder|Disease or Syndrome|Hospital Course|8229,8242|false|false|false|C0521530|Lung consolidation|Consolidation
Event|Event|Hospital Course|8229,8242|false|false|false|||Consolidation
Finding|Functional Concept|Hospital Course|8246,8250|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8246,8261|false|false|false|C1261077|Structure of left lower lobe of lung|left lower lobe
Anatomy|Body Location or Region|Hospital Course|8251,8256|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|8251,8256|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8251,8261|false|false|false|C0225758|Structure of lower lobe of lung|lower lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8257,8261|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|8257,8261|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Finding|Finding|Hospital Course|8278,8284|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8278,8284|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|Hospital Course|8285,8294|false|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|8285,8294|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|8285,8294|false|true|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|Hospital Course|8298,8307|false|true|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|8298,8307|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|8298,8307|false|true|false|C3714514|Infection|infection
Event|Event|Hospital Course|8321,8332|false|false|false|||progression
Finding|Functional Concept|Hospital Course|8321,8332|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|8321,8332|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Hospital Course|8336,8343|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|8336,8343|false|false|false|||disease
Finding|Finding|Hospital Course|8357,8361|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|8357,8361|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|8357,8361|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|8362,8368|false|false|false|||course
Event|Event|Hospital Course|8372,8382|false|false|false|||infiltrate
Finding|Functional Concept|Hospital Course|8372,8382|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Intellectual Product|Hospital Course|8372,8382|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Finding|Pathologic Function|Hospital Course|8372,8382|false|false|false|C0332448;C1546677;C1549537|Administration Method - Infiltrate;Infiltration|infiltrate
Event|Event|Hospital Course|8384,8395|false|false|false|||development
Finding|Functional Concept|Hospital Course|8384,8395|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|Hospital Course|8384,8395|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Procedure|Diagnostic Procedure|Hospital Course|8409,8416|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|8412,8416|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|8412,8416|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|8429,8440|false|false|false|||radiologist
Finding|Intellectual Product|Hospital Course|8429,8440|false|false|false|C1549438|Procedure Practitioner Identifier Code Type - Radiologist|radiologist
Event|Event|Hospital Course|8442,8451|false|false|false|||concluded
Event|Event|Hospital Course|8471,8478|false|false|false|||changes
Finding|Functional Concept|Hospital Course|8471,8478|false|false|false|C0392747|Changing|changes
Event|Event|Hospital Course|8479,8483|false|false|false|||seen
Finding|Finding|Hospital Course|8489,8495|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|8489,8495|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|8496,8502|false|false|false|||caused
Disorder|Neoplastic Process|Hospital Course|8511,8516|false|false|false|C0007131||NSCLC
Event|Event|Hospital Course|8511,8516|false|false|false|||NSCLC
Disorder|Disease or Syndrome|Hospital Course|8525,8534|true|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|8525,8534|true|false|false|||pneumonia
Event|Event|Hospital Course|8559,8564|true|false|false|||ruled
Event|Event|Hospital Course|8582,8588|false|false|false|||course
Drug|Antibiotic|Hospital Course|8592,8603|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|Hospital Course|8592,8603|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|Hospital Course|8592,8603|false|false|false|||ceftriaxone
Drug|Antibiotic|Hospital Course|8605,8617|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|8605,8617|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|8605,8617|false|false|false|||levofloxacin
Event|Event|Hospital Course|8641,8649|false|false|false|||narrowed
Drug|Antibiotic|Hospital Course|8653,8665|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|8653,8665|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|8653,8665|false|false|false|||levofloxacin
Finding|Finding|Hospital Course|8666,8671|false|false|false|C0439044|Living Alone|alone
Disorder|Disease or Syndrome|Hospital Course|8673,8678|true|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|Hospital Course|8673,8678|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|Hospital Course|8673,8687|true|false|false|C0200949|Blood culture|Blood cultures
Event|Event|Hospital Course|8679,8687|true|false|false|||cultures
Finding|Idea or Concept|Hospital Course|8679,8687|true|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|Hospital Course|8692,8698|true|false|false|||growth
Finding|Finding|Hospital Course|8692,8698|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organ or Tissue Function|Hospital Course|8692,8698|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Organism Function|Hospital Course|8692,8698|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Finding|Physiologic Function|Hospital Course|8692,8698|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|growth
Phenomenon|Phenomenon or Process|Hospital Course|8692,8698|true|false|false|C2911660|Growth action|growth
Finding|Body Substance|Hospital Course|8717,8723|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|8717,8723|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Event|Event|Hospital Course|8724,8732|false|false|false|||cultures
Finding|Idea or Concept|Hospital Course|8724,8732|false|true|false|C0010453|Culture (Anthropological)|cultures
Event|Event|Hospital Course|8757,8769|false|false|false|||contaminated
Anatomy|Body Space or Junction|Hospital Course|8775,8779|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8775,8779|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8775,8779|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8775,8779|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|8780,8785|false|false|false|||flora
Finding|Body Substance|Hospital Course|8787,8792|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|Hospital Course|8787,8792|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|Hospital Course|8787,8792|true|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Event|Event|Hospital Course|8793,8803|false|false|false|||legionella
Event|Event|Hospital Course|8804,8812|false|false|false|||negative
Finding|Classification|Hospital Course|8804,8812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|8804,8812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|8804,8812|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|Hospital Course|8814,8821|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8814,8821|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8814,8821|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|8827,8834|false|false|false|||improve
Drug|Antibiotic|Hospital Course|8851,8862|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|8851,8862|false|false|false|||antibiotics
Drug|Organic Chemical|Hospital Course|8878,8886|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|8878,8886|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|8878,8886|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|8878,8886|false|false|false|||complete
Finding|Functional Concept|Hospital Course|8878,8886|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8878,8886|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8894,8897|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8894,8897|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|8898,8904|false|false|false|||course
Drug|Antibiotic|Hospital Course|8908,8920|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|8908,8920|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|8908,8920|false|false|false|||levofloxacin
Disorder|Neoplastic Process|Hospital Course|8927,8932|false|false|false|C0007131||NSCLC
Attribute|Clinical Attribute|Hospital Course|8934,8939|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|8934,8942|false|false|false|C0441772|Stage level 4|stage IV
Event|Event|Hospital Course|8940,8942|false|false|false|||IV
Event|Event|Hospital Course|8968,8980|true|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|8968,8980|true|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8968,8980|true|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Classification|Hospital Course|8984,8994|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|8984,8994|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Event|Event|Hospital Course|9017,9025|false|false|false|||planning
Event|Event|Hospital Course|9029,9038|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|9029,9038|false|false|false|C0549178|Continuous|continued
Event|Event|Hospital Course|9040,9052|false|false|false|||surveillance
Event|Occupational Activity|Hospital Course|9040,9052|false|false|false|C0684245|legal surveillance|surveillance
Finding|Functional Concept|Hospital Course|9040,9052|false|false|false|C0220920|surveillance aspects|surveillance
Procedure|Health Care Activity|Hospital Course|9040,9052|false|false|false|C0733511|Medical Surveillance|surveillance
Disorder|Disease or Syndrome|Hospital Course|9058,9062|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|Hospital Course|9058,9062|false|false|false|||plan
Finding|Functional Concept|Hospital Course|9058,9062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|9058,9062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|9058,9062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Finding|Hospital Course|9067,9075|false|false|false|C0332149|Possible|possible
Event|Event|Hospital Course|9095,9103|false|false|false|||systemic
Finding|Functional Concept|Hospital Course|9095,9103|false|true|false|C0205373;C5849094|Systemic;Systemic Route of Administration|systemic
Event|Event|Hospital Course|9105,9117|false|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|9105,9117|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9105,9117|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Finding|Functional Concept|Hospital Course|9121,9132|false|false|false|C0231220|Symptomatic|symptomatic
Event|Event|Hospital Course|9133,9144|false|false|false|||progression
Finding|Functional Concept|Hospital Course|9133,9144|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|9133,9144|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Hospital Course|9148,9159|false|false|false|C0017925|Glycogen Storage Disease Type VI|her disease
Disorder|Disease or Syndrome|Hospital Course|9152,9159|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|9152,9159|false|false|false|||disease
Event|Event|Hospital Course|9163,9168|false|false|false|||noted
Procedure|Diagnostic Procedure|Hospital Course|9171,9178|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|9174,9178|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|9174,9178|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|9183,9193|false|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|9183,9193|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|9183,9193|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Disorder|Disease or Syndrome|Hospital Course|9197,9204|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|9197,9204|false|false|false|||disease
Finding|Pathologic Function|Hospital Course|9197,9216|false|false|false|C0242656|Disease Progression|disease progression
Event|Event|Hospital Course|9205,9216|false|false|false|||progression
Finding|Functional Concept|Hospital Course|9205,9216|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|9205,9216|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Event|Event|Hospital Course|9221,9229|false|false|false|||obtained
Event|Event|Hospital Course|9239,9243|false|false|false|||show
Event|Event|Hospital Course|9252,9263|false|false|false|||progression
Finding|Functional Concept|Hospital Course|9252,9263|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|9252,9263|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Event|Event|Hospital Course|9273,9278|false|false|false|||plans
Event|Event|Hospital Course|9282,9287|false|false|false|||weigh
Event|Event|Hospital Course|9292,9297|false|false|false|||risks
Finding|Idea or Concept|Hospital Course|9292,9297|false|false|false|C0035647|Risk|risks
Event|Event|Hospital Course|9303,9311|false|false|false|||benefits
Finding|Functional Concept|Hospital Course|9315,9325|false|false|false|C1524062|Additional|additional
Event|Event|Hospital Course|9326,9338|false|false|false|||chemotherapy
Finding|Functional Concept|Hospital Course|9326,9338|false|false|true|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9326,9338|false|false|true|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Hospital Course|9355,9366|false|false|false|||complicated
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9374,9380|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|9374,9380|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|9374,9380|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|9374,9380|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9374,9380|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Finding|Pathologic Function|Hospital Course|9374,9392|false|false|false|C0151746|Abnormal renal function|kidney dysfunction
Disorder|Disease or Syndrome|Hospital Course|9381,9392|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Hospital Course|9381,9392|false|false|false|||dysfunction
Finding|Conceptual Entity|Hospital Course|9381,9392|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Hospital Course|9381,9392|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Hospital Course|9381,9392|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|Hospital Course|9403,9416|false|false|false|||comorbidities
Finding|Finding|Hospital Course|9403,9416|false|false|false|C0009488|Comorbidity|comorbidities
Event|Event|Hospital Course|9422,9427|false|false|false|||plans
Event|Event|Hospital Course|9431,9437|false|false|false|||repeat
Procedure|Diagnostic Procedure|Hospital Course|9442,9449|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Hospital Course|9445,9449|false|false|false|||scan
Procedure|Diagnostic Procedure|Hospital Course|9445,9449|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Hospital Course|9459,9468|false|false|false|||completes
Drug|Antibiotic|Hospital Course|9474,9485|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Hospital Course|9474,9485|false|false|false|||antibiotics
Event|Event|Hospital Course|9497,9505|false|false|false|||evaluate
Event|Activity|Hospital Course|9510,9514|false|false|false|C0871208|Rating (action)|rate
Event|Event|Hospital Course|9510,9514|false|false|false|||rate
Finding|Idea or Concept|Hospital Course|9510,9514|false|false|false|C1549480|Amount type - Rate|rate
Disorder|Disease or Syndrome|Hospital Course|9518,9525|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|9518,9525|false|false|false|||disease
Finding|Pathologic Function|Hospital Course|9518,9537|false|false|false|C0242656|Disease Progression|disease progression
Event|Event|Hospital Course|9526,9537|false|false|false|||progression
Finding|Functional Concept|Hospital Course|9526,9537|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Hospital Course|9526,9537|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Hospital Course|9548,9551|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9548,9551|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|9548,9551|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|9548,9551|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|9548,9551|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|9548,9551|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|9548,9551|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9548,9551|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|9560,9567|true|false|false|||Patient
Finding|Body Substance|Hospital Course|9560,9567|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9560,9567|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9560,9567|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Anatomy|Body Location or Region|Hospital Course|9576,9581|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|9576,9581|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|9576,9586|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|9576,9586|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|9582,9586|true|true|false|C2598155||pain
Event|Event|Hospital Course|9582,9586|true|false|false|||pain
Finding|Functional Concept|Hospital Course|9582,9586|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9582,9586|true|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|9597,9600|false|false|false|||EKG
Finding|Intellectual Product|Hospital Course|9597,9600|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|9597,9600|false|false|false|C1623258|Electrocardiography|EKG
Finding|Finding|Hospital Course|9606,9609|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|9606,9609|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9614,9625|false|false|false|C0011570|Mental Depression|depressions
Event|Event|Hospital Course|9614,9625|false|false|false|||depressions
Attribute|Clinical Attribute|Hospital Course|9627,9637|false|false|false|C0005516|Biological Markers|Biomarkers
Event|Event|Hospital Course|9638,9644|false|false|false|||cycled
Event|Event|Hospital Course|9649,9657|false|false|false|||negative
Finding|Classification|Hospital Course|9649,9657|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9649,9657|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9649,9657|false|false|false|C5237010|Expression Negative|negative
Finding|Body Substance|Hospital Course|9662,9669|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9662,9669|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9662,9669|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|9671,9680|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|9684,9688|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|9684,9688|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|9684,9688|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|9689,9693|false|false|false|||beta
Finding|Intellectual Product|Hospital Course|9689,9693|false|false|false|C0439096|Greek letter beta|beta
Drug|Pharmacologic Substance|Hospital Course|9689,9701|false|false|false|C0001645|Adrenergic beta-Antagonists|beta-blocker
Event|Event|Hospital Course|9694,9701|false|false|false|||blocker
Finding|Finding|Hospital Course|9707,9716|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Event|Event|Hospital Course|9717,9721|false|false|false|||dose
Attribute|Clinical Attribute|Hospital Course|9730,9738|false|false|false|C3172260||relative
Finding|Idea or Concept|Hospital Course|9730,9738|false|false|false|C1546849|Living Arrangement - Relative|relative
Event|Event|Hospital Course|9739,9750|false|false|false|||hypotension
Finding|Finding|Hospital Course|9739,9750|false|false|false|C0020649|Hypotension|hypotension
Event|Event|Hospital Course|9760,9770|false|false|false|||maintained
Drug|Organic Chemical|Hospital Course|9774,9781|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|9774,9781|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|9774,9781|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|9783,9789|false|false|false|C0633084|Plavix|plavix
Drug|Pharmacologic Substance|Hospital Course|9783,9789|false|false|false|C0633084|Plavix|plavix
Event|Event|Hospital Course|9783,9789|false|false|false|||plavix
Drug|Organic Chemical|Hospital Course|9796,9802|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Hospital Course|9796,9802|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|Hospital Course|9796,9802|false|false|false|||statin
Finding|Gene or Genome|Hospital Course|9796,9802|false|false|false|C1414273|EEF1A2 gene|statin
Event|Event|Hospital Course|9808,9815|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|9808,9815|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|9808,9815|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|9808,9828|false|false|false|C1135194|Chronic systolic heart failure|chronic systolic CHF
Finding|Organ or Tissue Function|Hospital Course|9816,9824|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Hospital Course|9816,9828|false|false|false|C2039715|systolic congestive heart failure|systolic CHF
Anatomy|Body Space or Junction|Hospital Course|9825,9828|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|9825,9828|false|false|false|C0018802|Congestive heart failure|CHF
Attribute|Clinical Attribute|Hospital Course|9830,9834|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Procedure|Diagnostic Procedure|Hospital Course|9830,9834|false|false|false|C3837267|LVEF (procedure)|LVEF
Procedure|Diagnostic Procedure|Hospital Course|9842,9845|false|false|false|C0430462|Transthoracic echocardiography|TTE
Finding|Finding|Hospital Course|9852,9856|false|false|false|C5575035|Well (answer to question)|Well
Event|Event|Hospital Course|9857,9868|false|false|false|||compensated
Event|Event|Hospital Course|9873,9882|false|false|false|||described
Drug|Organic Chemical|Hospital Course|9890,9895|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9890,9895|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|9890,9895|false|false|false|||lasix
Event|Event|Hospital Course|9900,9904|false|false|false|||held
Event|Event|Hospital Course|9912,9919|false|false|false|||blocker
Anatomy|Body Location or Region|Hospital Course|9935,9940|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|9935,9940|false|false|false|C2003888|Lower (action)|lower
Attribute|Clinical Attribute|Hospital Course|9952,9960|false|false|false|C3172260||relative
Finding|Idea or Concept|Hospital Course|9952,9960|false|false|false|C1546849|Living Arrangement - Relative|relative
Event|Event|Hospital Course|9961,9972|false|false|false|||hypotension
Finding|Finding|Hospital Course|9961,9972|false|false|false|C0020649|Hypotension|hypotension
Finding|Sign or Symptom|Hospital Course|9978,9988|false|false|false|C0239313|exercise induced|exertional
Finding|Finding|Hospital Course|9978,10000|false|false|false|C0241324|Exertional tachycardia|exertional tachycardia
Event|Event|Hospital Course|9989,10000|false|false|false|||tachycardia
Finding|Finding|Hospital Course|9989,10000|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Disorder|Disease or Syndrome|Hospital Course|10007,10010|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Hospital Course|10011,10016|false|false|false|C1300072|Tumor stage|stage
Drug|Biologically Active Substance|Hospital Course|10022,10032|false|false|false|C0010294|creatinine|Creatinine
Drug|Organic Chemical|Hospital Course|10022,10032|false|false|false|C0010294|creatinine|Creatinine
Event|Event|Hospital Course|10022,10032|false|false|false|||Creatinine
Finding|Physiologic Function|Hospital Course|10022,10032|false|false|false|C4551889|Creatinine metabolic function|Creatinine
Procedure|Laboratory Procedure|Hospital Course|10022,10032|false|false|false|C0201975|Creatinine measurement|Creatinine
Event|Event|Hospital Course|10036,10045|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|10036,10045|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Hospital Course|10071,10075|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|10071,10075|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|10071,10075|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|10079,10088|false|false|false|||discharge
Finding|Body Substance|Hospital Course|10079,10088|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10079,10088|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10079,10088|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10079,10088|false|false|false|C0030685|Patient Discharge|discharge
Drug|Substance|Hospital Course|10115,10121|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Hospital Course|10115,10121|false|false|false|||fluids
Finding|Body Substance|Hospital Course|10115,10121|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10115,10121|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Body Space or Junction|Hospital Course|10130,10133|false|false|false|C0228479|Structure of intraculminate fissure|ICU
Event|Event|Hospital Course|10130,10133|false|false|false|||ICU
Finding|Intellectual Product|Hospital Course|10130,10133|false|false|false|C4554035|Inventory of Callous-Unemotional Traits|ICU
Drug|Organic Chemical|Hospital Course|10142,10147|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|10142,10147|false|false|false|C0699992|Lasix|lasix
Event|Event|Hospital Course|10142,10147|false|false|false|||lasix
Event|Event|Hospital Course|10152,10156|false|false|false|||held
Finding|Body Substance|Hospital Course|10175,10182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10175,10182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10175,10182|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|Hospital Course|10197,10202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|10197,10202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|10197,10202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Attribute|Clinical Attribute|Hospital Course|10197,10209|false|false|false|C0232856;C0489132||urine output
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10197,10209|false|false|false|C2094175|monitoring of urine output for fluid balance|urine output
Event|Event|Hospital Course|10203,10209|false|false|false|||output
Finding|Conceptual Entity|Hospital Course|10203,10209|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|10203,10209|false|false|false|C3251815|Measurement of fluid output|output
Finding|Finding|Hospital Course|10217,10227|false|false|false|C0302870|microcytic|Microcytic
Disorder|Disease or Syndrome|Hospital Course|10217,10234|false|false|false|C5194182|Microcytic anemia|Microcytic anemia
Disorder|Disease or Syndrome|Hospital Course|10228,10234|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|10228,10234|false|false|false|||anemia
Event|Event|Hospital Course|10239,10251|false|false|false|||presentation
Finding|Idea or Concept|Hospital Course|10239,10251|false|false|false|C0449450|Presentation|presentation
Finding|Body Substance|Hospital Course|10253,10260|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10253,10260|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10253,10260|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Laboratory Procedure|Hospital Course|10263,10266|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10263,10266|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Finding|Finding|Hospital Course|10267,10273|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10267,10273|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|10275,10291|false|false|false|||hemoconcentrated
Event|Event|Hospital Course|10293,10299|false|false|false|||Follow
Event|Event|Hospital Course|10303,10306|false|false|false|||Hct
Procedure|Laboratory Procedure|Hospital Course|10303,10306|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10303,10306|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Event|Event|Hospital Course|10307,10312|false|false|false|||found
Event|Event|Hospital Course|10326,10331|true|false|false|||signs
Finding|Finding|Hospital Course|10326,10331|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|10326,10331|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|Hospital Course|10336,10344|true|false|false|||bleeding
Finding|Pathologic Function|Hospital Course|10336,10344|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|10348,10352|true|false|false|||exam
Finding|Functional Concept|Hospital Course|10348,10352|true|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|10348,10352|true|false|false|C0582103|Medical Examination|exam
Finding|Body Substance|Hospital Course|10354,10361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10354,10361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10354,10361|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|10362,10372|false|false|false|||transfused
Event|Event|Hospital Course|10373,10379|false|false|false|||2units
Event|Event|Hospital Course|10383,10387|false|false|false|||pRBC
Event|Event|Hospital Course|10396,10403|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|10396,10403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|10396,10403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|10396,10403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|10396,10406|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|10407,10410|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10407,10410|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|10407,10410|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|10407,10410|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|10407,10410|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|10407,10410|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|10407,10410|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10407,10410|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|10428,10437|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10428,10437|false|false|false|C0439775|Elevation procedure|elevation
Attribute|Clinical Attribute|Hospital Course|10441,10451|false|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|Hospital Course|10441,10451|false|false|false|||hematocrit
Finding|Finding|Hospital Course|10441,10451|false|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|Hospital Course|10441,10451|false|false|false|C0018935|Hematocrit Measurement|hematocrit
Attribute|Clinical Attribute|Hospital Course|10458,10468|false|false|false|C1542366|hematocrit attribute|hematocrit
Event|Event|Hospital Course|10458,10468|false|false|false|||hematocrit
Finding|Finding|Hospital Course|10458,10468|false|false|false|C0518014|Hematocrit level|hematocrit
Procedure|Laboratory Procedure|Hospital Course|10458,10468|false|false|false|C0018935|Hematocrit Measurement|hematocrit
Event|Event|Hospital Course|10473,10479|false|false|false|||remain
Event|Event|Hospital Course|10499,10505|false|false|false|||course
Event|Event|Hospital Course|10506,10515|false|false|false|||following
Event|Event|Hospital Course|10517,10527|false|false|false|||tranfusion
Event|Event|Hospital Course|10541,10549|false|false|false|||transfer
Finding|Functional Concept|Hospital Course|10541,10549|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|Hospital Course|10541,10549|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|Hospital Course|10541,10549|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Body Substance|Hospital Course|10564,10571|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10564,10571|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10564,10571|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|10574,10579|false|false|false|||stool
Finding|Body Substance|Hospital Course|10574,10579|false|false|false|C0015733|Feces|stool
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|10581,10587|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|Hospital Course|10581,10587|false|false|false|C0018302|guaiac|guaiac
Event|Event|Hospital Course|10581,10587|false|false|false|||guaiac
Disorder|Cell or Molecular Dysfunction|Hospital Course|10592,10600|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|Hospital Course|10592,10600|false|false|false|||positive
Finding|Classification|Hospital Course|10592,10600|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|10592,10600|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Event|Event|Hospital Course|10612,10616|false|false|false|||call
Event|Event|Hospital Course|10629,10633|false|false|false|||work
Event|Occupational Activity|Hospital Course|10629,10633|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|10629,10636|false|false|false|C0750430|Work-up|work-up
Finding|Body Substance|Hospital Course|10643,10650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10643,10650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10643,10650|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|10653,10659|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|10653,10659|false|false|false|||anemia
Finding|Idea or Concept|Hospital Course|10663,10674|false|false|false|C0750501|most likely|most likely
Finding|Finding|Hospital Course|10668,10674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10668,10674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|Hospital Course|10675,10684|false|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Hospital Course|10675,10684|false|false|false|||secondary
Finding|Functional Concept|Hospital Course|10675,10684|false|true|false|C1522484|metastatic qualifier|secondary
Finding|Intellectual Product|Hospital Course|10688,10693|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|Hospital Course|10688,10706|false|true|false|C0333361|Acute inflammation|acute inflammation
Event|Event|Hospital Course|10694,10706|false|false|false|||inflammation
Finding|Pathologic Function|Hospital Course|10694,10706|false|false|false|C0021368|Inflammation|inflammation
Finding|Mental Process|Hospital Course|10715,10722|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|10726,10736|false|false|false|C4722602|Underlying|underlying
Finding|Intellectual Product|Hospital Course|10737,10744|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|10737,10744|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|10737,10752|false|false|false|C0008679|Chronic disease|chronic disease
Disorder|Disease or Syndrome|Hospital Course|10745,10752|false|false|false|C0012634|Disease|disease
Event|Event|Hospital Course|10745,10752|false|false|false|||disease
Attribute|Clinical Attribute|Hospital Course|10759,10770|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|10759,10770|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|10759,10770|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|10759,10770|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|10759,10783|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|10774,10783|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|10774,10783|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|10785,10795|false|false|false|C0051696|amlodipine|amlodipine
Drug|Pharmacologic Substance|Hospital Course|10785,10795|false|false|false|C0051696|amlodipine|amlodipine
Drug|Biomedical or Dental Material|Hospital Course|10801,10807|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10813,10819|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|10823,10831|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10826,10831|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10826,10831|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|10832,10841|false|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|Hospital Course|10832,10841|false|false|false|C1170480|One Daily|one daily
Drug|Vitamin|Hospital Course|10832,10841|false|false|false|C1170480|One Daily|one daily
Drug|Organic Chemical|Hospital Course|10844,10856|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|10844,10856|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|10844,10856|false|false|false|||atorvastatin
Drug|Organic Chemical|Hospital Course|10858,10865|false|false|false|C0593906|Lipitor|Lipitor
Drug|Pharmacologic Substance|Hospital Course|10858,10865|false|false|false|C0593906|Lipitor|Lipitor
Drug|Biomedical or Dental Material|Hospital Course|10873,10879|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|10885,10891|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|10895,10903|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10898,10903|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10898,10903|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|10916,10926|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Pharmacologic Substance|Hospital Course|10916,10926|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Vitamin|Hospital Course|10916,10926|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Event|Event|Hospital Course|10916,10926|false|false|false|||calcitriol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10936,10943|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10936,10943|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10936,10943|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10947,10954|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|10947,10954|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|10947,10954|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|10958,10966|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|10961,10966|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|10961,10966|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|10967,10971|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|10967,10977|false|false|false|C3537736|Once A Day|once a day
Event|Event|Hospital Course|10974,10977|false|false|false|||day
Finding|Idea or Concept|Hospital Course|10974,10977|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|10974,10977|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|10978,10989|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|10978,10989|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|Hospital Course|10978,10989|false|false|false|||clopidogrel
Drug|Organic Chemical|Hospital Course|10991,10997|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Hospital Course|10991,10997|false|false|false|C0633084|Plavix|Plavix
Drug|Biomedical or Dental Material|Hospital Course|11005,11011|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11014,11020|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|11024,11032|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11027,11032|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11027,11032|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|11033,11037|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|Hospital Course|11041,11044|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11041,11044|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|11046,11056|false|false|false|C0016410|folic acid|folic acid
Drug|Pharmacologic Substance|Hospital Course|11046,11056|false|false|false|C0016410|folic acid|folic acid
Drug|Vitamin|Hospital Course|11046,11056|false|false|false|C0016410|folic acid|folic acid
Procedure|Laboratory Procedure|Hospital Course|11046,11056|false|false|false|C0523631|Folic acid measurement|folic acid
Event|Event|Hospital Course|11052,11056|false|false|false|||acid
Drug|Biomedical or Dental Material|Hospital Course|11063,11069|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11074,11080|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|11084,11092|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11087,11092|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11087,11092|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11093,11102|false|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|Hospital Course|11093,11102|false|false|false|C1170480|One Daily|one daily
Drug|Vitamin|Hospital Course|11093,11102|false|false|false|C1170480|One Daily|one daily
Drug|Organic Chemical|Hospital Course|11104,11114|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|11104,11114|false|false|false|C0016860|furosemide|furosemide
Event|Event|Hospital Course|11104,11114|false|false|false|||furosemide
Drug|Biomedical or Dental Material|Hospital Course|11121,11127|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11131,11137|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|11141,11149|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11144,11149|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11144,11149|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11156,11166|false|false|false|C0023992|loperamide|loperamide
Drug|Pharmacologic Substance|Hospital Course|11156,11166|false|false|false|C0023992|loperamide|loperamide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11172,11179|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|11172,11179|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|11172,11179|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11185,11192|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|11185,11192|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|11185,11192|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|11196,11204|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11199,11204|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11199,11204|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|11225,11231|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|11233,11242|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|11233,11242|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|11233,11242|false|false|false|||lorazepam
Drug|Biomedical or Dental Material|Hospital Course|11250,11256|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11261,11267|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11261,11267|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|11271,11279|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11274,11279|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11274,11279|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Hospital Course|11293,11299|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|11304,11310|false|false|false|C4255480||Nausea
Event|Event|Hospital Course|11304,11310|false|false|false|||Nausea
Finding|Sign or Symptom|Hospital Course|11304,11310|false|false|false|C0027497|Nausea|Nausea
Drug|Organic Chemical|Hospital Course|11312,11322|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|11312,11322|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|11312,11331|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|Hospital Course|11312,11331|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|Hospital Course|11323,11331|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|Hospital Course|11323,11331|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|Hospital Course|11323,11331|false|false|false|||tartrate
Drug|Organic Chemical|Hospital Course|11333,11342|false|false|false|C0700776|Lopressor|Lopressor
Drug|Pharmacologic Substance|Hospital Course|11333,11342|false|false|false|C0700776|Lopressor|Lopressor
Drug|Biomedical or Dental Material|Hospital Course|11350,11356|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11362,11368|false|false|false|C0039225|Tablet Dosage Form|Tablet
Anatomy|Body Location or Region|Hospital Course|11376,11381|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11376,11381|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11405,11413|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|11405,11413|false|false|false|C0040610|tramadol|tramadol
Event|Event|Hospital Course|11405,11413|false|false|false|||tramadol
Procedure|Laboratory Procedure|Hospital Course|11405,11413|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|11420,11426|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11443,11449|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11443,11449|false|false|false|||Tablet
Finding|Functional Concept|Hospital Course|11453,11461|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11456,11461|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11456,11461|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|11469,11474|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|11469,11474|false|false|false|||times
Finding|Idea or Concept|Hospital Course|11477,11480|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11477,11480|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|11484,11490|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|11495,11499|false|false|false|C2598155||Pain
Event|Event|Hospital Course|11495,11499|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|11495,11499|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|11495,11499|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|11502,11511|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|Hospital Course|11502,11511|false|false|false|C0040805|trazodone|trazodone
Event|Event|Hospital Course|11502,11511|false|false|false|||trazodone
Drug|Biomedical or Dental Material|Hospital Course|11518,11524|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11530,11536|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|11540,11548|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11543,11548|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11543,11548|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11549,11558|false|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|Hospital Course|11549,11558|false|false|false|C1170480|One Daily|one daily
Drug|Vitamin|Hospital Course|11549,11558|false|false|false|C1170480|One Daily|one daily
Event|Event|Hospital Course|11563,11569|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|11571,11578|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|11571,11578|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|11571,11578|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Hospital Course|11585,11591|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11585,11591|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|11585,11601|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Biomedical or Dental Material|Hospital Course|11605,11611|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|11615,11623|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|11618,11623|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11618,11623|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11624,11633|false|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|Hospital Course|11624,11633|false|false|false|C1170480|One Daily|one daily
Drug|Vitamin|Hospital Course|11624,11633|false|false|false|C1170480|One Daily|one daily
Drug|Organic Chemical|Hospital Course|11635,11645|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|11635,11645|false|false|false|C0034665|ranitidine|ranitidine
Drug|Organic Chemical|Hospital Course|11635,11649|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Drug|Pharmacologic Substance|Hospital Course|11635,11649|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Disorder|Neoplastic Process|Hospital Course|11646,11649|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|11646,11649|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|11646,11649|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|11646,11649|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|11646,11649|false|false|false|||HCl
Drug|Organic Chemical|Hospital Course|11651,11663|false|false|false|C4765118|Acid Control|Acid Control
Drug|Pharmacologic Substance|Hospital Course|11651,11663|false|false|false|C4765118|Acid Control|Acid Control
Drug|Organic Chemical|Hospital Course|11656,11663|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|Control
Drug|Pharmacologic Substance|Hospital Course|11656,11663|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|Control
Drug|Substance|Hospital Course|11656,11663|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|Control
Event|Event|Hospital Course|11656,11663|false|false|false|||Control
Finding|Conceptual Entity|Hospital Course|11656,11663|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|Control
Finding|Functional Concept|Hospital Course|11656,11663|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|Control
Finding|Idea or Concept|Hospital Course|11656,11663|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|Control
Drug|Biomedical or Dental Material|Hospital Course|11672,11678|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11684,11690|false|false|false|C0039225|Tablet Dosage Form|Tablet
Anatomy|Body Location or Region|Hospital Course|11698,11703|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|11698,11703|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Organic Chemical|Hospital Course|11704,11713|false|false|false|C1170480|One Daily|one daily
Drug|Pharmacologic Substance|Hospital Course|11704,11713|false|false|false|C1170480|One Daily|one daily
Drug|Vitamin|Hospital Course|11704,11713|false|false|false|C1170480|One Daily|one daily
Event|Event|Hospital Course|11717,11726|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|11717,11726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11717,11726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11717,11726|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11717,11726|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11717,11738|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|11727,11738|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11727,11738|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|11727,11738|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|11727,11738|false|false|false|C4284232|Medications|Medications
Drug|Biologically Active Substance|Hospital Course|11743,11749|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|11743,11749|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|11743,11749|false|false|false|C0030054|oxygen|oxygen
Event|Event|Hospital Course|11743,11749|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11743,11749|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Hospital Course|11754,11764|false|false|false|||continuous
Finding|Idea or Concept|Hospital Course|11754,11764|false|false|false|C0549178|Continuous|continuous
Attribute|Clinical Attribute|Hospital Course|11766,11771|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|Hospital Course|11766,11771|false|false|false|||pulse
Finding|Physiologic Function|Hospital Course|11766,11771|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|Hospital Course|11766,11771|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|Hospital Course|11766,11771|false|false|false|C0034107|Pulse taking|pulse
Event|Event|Hospital Course|11772,11776|false|false|false|||dose
Event|Event|Hospital Course|11781,11792|false|false|false|||portability
Anatomy|Body Location or Region|Hospital Course|11797,11801|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11797,11801|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|11797,11801|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|11797,11801|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|11797,11808|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Hospital Course|11802,11808|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Hospital Course|11802,11808|false|false|false|||cancer
Drug|Antibiotic|Hospital Course|11812,11824|false|false|false|C0282386|levofloxacin|levofloxacin
Drug|Organic Chemical|Hospital Course|11812,11824|false|false|false|C0282386|levofloxacin|levofloxacin
Event|Event|Hospital Course|11812,11824|false|false|false|||levofloxacin
Drug|Biomedical or Dental Material|Hospital Course|11832,11838|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11852,11858|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11852,11858|false|false|false|||Tablet
Event|Event|Hospital Course|11862,11866|false|false|false|||Q48H
Event|Event|Hospital Course|11868,11873|false|false|false|||every
Finding|Intellectual Product|Hospital Course|11868,11873|false|false|false|C1720374|Every - dosing instruction fragment|every
Finding|Idea or Concept|Hospital Course|11903,11906|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|11903,11906|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|11920,11926|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11920,11926|false|false|false|||Tablet
Finding|Idea or Concept|Hospital Course|11931,11938|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|11946,11958|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11946,11958|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|11946,11958|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|11965,11971|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|11985,11991|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|11992,11994|false|false|false|||PO
Drug|Organic Chemical|Hospital Course|12016,12026|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|12016,12026|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Hospital Course|12016,12026|false|false|false|||metoprolol
Drug|Organic Chemical|Hospital Course|12016,12035|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|Hospital Course|12016,12035|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|Hospital Course|12027,12035|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|Hospital Course|12027,12035|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|Hospital Course|12027,12035|false|false|false|||tartrate
Drug|Biomedical or Dental Material|Hospital Course|12042,12048|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|12062,12068|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|12081,12084|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12081,12084|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|12098,12102|false|false|false|||THIS
Event|Event|Hospital Course|12108,12114|false|false|false|||CHANGE
Finding|Functional Concept|Hospital Course|12108,12114|false|false|false|C0392747|Changing|CHANGE
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12108,12114|false|false|false|C4319952|Change - procedure|CHANGE
Event|Event|Hospital Course|12134,12141|false|false|false|||EVENING
Event|Event|Hospital Course|12143,12149|false|false|false|||DOSING
Drug|Organic Chemical|Hospital Course|12156,12164|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|12156,12164|false|false|false|C1692318|docusate|docusate
Event|Event|Hospital Course|12156,12164|false|false|false|||docusate
Drug|Organic Chemical|Hospital Course|12156,12171|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|12156,12171|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|12165,12171|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|12165,12171|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|12165,12171|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|12165,12171|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|12165,12171|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|12165,12171|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12179,12186|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|12179,12186|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|12179,12186|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12200,12207|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|12200,12207|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|12200,12207|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12211,12214|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12211,12214|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12211,12214|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|12211,12214|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|12211,12214|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|12219,12224|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|12227,12230|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12227,12230|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|12233,12237|false|false|false|C1948035|Hold (action)|hold
Event|Event|Hospital Course|12233,12237|false|false|false|||hold
Finding|Functional Concept|Hospital Course|12233,12237|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|Hospital Course|12233,12237|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Sign or Symptom|Hospital Course|12241,12253|false|false|false|C0011991;C2129214|Diarrhea;Loose stool|loose stools
Attribute|Clinical Attribute|Hospital Course|12247,12253|false|false|false|C0489144||stools
Event|Event|Hospital Course|12247,12253|false|false|false|||stools
Finding|Body Substance|Hospital Course|12247,12253|false|false|false|C0015733|Feces|stools
Drug|Organic Chemical|Hospital Course|12260,12269|false|false|false|C0040805|trazodone|trazodone
Drug|Pharmacologic Substance|Hospital Course|12260,12269|false|false|false|C0040805|trazodone|trazodone
Event|Event|Hospital Course|12260,12269|false|false|false|||trazodone
Drug|Biomedical or Dental Material|Hospital Course|12276,12282|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|12296,12302|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12296,12302|false|false|false|||Tablet
Event|Event|Hospital Course|12326,12332|false|false|false|||needed
Drug|Pharmacologic Substance|Hospital Course|12337,12345|false|false|false|C1950154|Insomnia homeopathic medication|insomnia
Event|Event|Hospital Course|12337,12345|false|false|false|||insomnia
Finding|Sign or Symptom|Hospital Course|12337,12345|false|false|false|C0917801|Sleeplessness|insomnia
Drug|Organic Chemical|Hospital Course|12352,12363|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|12352,12363|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Biomedical or Dental Material|Hospital Course|12370,12376|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|12390,12396|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12390,12396|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|12421,12431|false|false|false|C0034665|ranitidine|ranitidine
Drug|Pharmacologic Substance|Hospital Course|12421,12431|false|false|false|C0034665|ranitidine|ranitidine
Event|Event|Hospital Course|12421,12431|false|false|false|||ranitidine
Drug|Organic Chemical|Hospital Course|12421,12435|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Drug|Pharmacologic Substance|Hospital Course|12421,12435|false|false|false|C0700466|ranitidine hydrochloride|ranitidine HCl
Disorder|Neoplastic Process|Hospital Course|12432,12435|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|12432,12435|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|12432,12435|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|12432,12435|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Hospital Course|12432,12435|false|false|false|||HCl
Drug|Biomedical or Dental Material|Hospital Course|12443,12449|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|12463,12469|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12463,12469|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|12494,12504|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Pharmacologic Substance|Hospital Course|12494,12504|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Drug|Vitamin|Hospital Course|12494,12504|false|false|false|C0006674;C3714610|Calcitriol Drug Class;calcitriol|calcitriol
Event|Event|Hospital Course|12494,12504|false|false|false|||calcitriol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12514,12521|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|12514,12521|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|12514,12521|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12535,12542|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|12535,12542|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|12535,12542|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|Hospital Course|12568,12578|false|false|false|C0016410|folic acid|folic acid
Drug|Pharmacologic Substance|Hospital Course|12568,12578|false|false|false|C0016410|folic acid|folic acid
Drug|Vitamin|Hospital Course|12568,12578|false|false|false|C0016410|folic acid|folic acid
Procedure|Laboratory Procedure|Hospital Course|12568,12578|false|false|false|C0523631|Folic acid measurement|folic acid
Event|Event|Hospital Course|12574,12578|false|false|false|||acid
Drug|Biomedical or Dental Material|Hospital Course|12584,12590|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12591,12594|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|12604,12610|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12604,12610|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|12636,12643|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|12636,12643|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|12636,12643|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Hospital Course|12650,12656|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|12650,12666|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12667,12670|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12667,12670|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|12667,12670|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|12667,12670|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|12680,12686|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|12680,12686|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Hospital Course|12680,12696|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Event|Event|Hospital Course|12688,12696|false|false|false|||Chewable
Event|Event|Hospital Course|12721,12730|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12721,12730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12721,12730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12721,12730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12721,12730|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|12721,12742|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|12721,12742|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|12731,12742|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|12731,12742|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|12731,12742|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|12744,12748|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|12744,12748|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|12744,12748|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|12744,12748|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|12754,12761|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|12754,12761|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|12764,12772|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|12764,12772|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|12780,12789|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|12780,12789|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12780,12789|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12780,12789|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12780,12789|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12780,12799|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|12790,12799|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|12790,12799|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|12790,12799|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|12790,12799|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|12790,12799|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|12820,12829|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Hospital Course|12820,12829|false|false|false|||pneumonia
Disorder|Neoplastic Process|Hospital Course|12836,12858|false|false|false|C0149925|Small cell carcinoma of lung|small cell lung cancer
Disorder|Neoplastic Process|Hospital Course|12836,12864|false|false|false|C0280249|stage, small cell lung cancer|small cell lung cancer stage
Anatomy|Cell|Hospital Course|12842,12846|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|12842,12846|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Anatomy|Body Location or Region|Hospital Course|12847,12851|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12847,12851|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|12847,12851|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|12847,12851|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Hospital Course|12847,12858|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Hospital Course|12847,12867|false|false|false|C0855005|Stage IV Lung Cancer AJCC v7|lung cancer stage IV
Disorder|Neoplastic Process|Hospital Course|12852,12858|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Diagnostic Procedure|Hospital Course|12852,12864|false|false|false|C0027646|Diagnostic Neoplasm Staging|cancer stage
Attribute|Clinical Attribute|Hospital Course|12859,12864|false|false|false|C1300072|Tumor stage|stage
Event|Event|Hospital Course|12859,12864|false|false|false|||stage
Finding|Intellectual Product|Hospital Course|12859,12867|false|false|false|C0441772|Stage level 4|stage IV
Event|Event|Hospital Course|12869,12880|false|false|false|||progressing
Finding|Functional Concept|Hospital Course|12869,12880|false|false|false|C0205329|Progressive|progressing
Disorder|Neoplastic Process|Hospital Course|12883,12892|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Hospital Course|12883,12892|false|false|false|C1522484|metastatic qualifier|SECONDARY
Event|Event|Hospital Course|12893,12902|false|false|false|||DIAGNOSES
Procedure|Diagnostic Procedure|Hospital Course|12893,12902|false|false|false|C0011900|Diagnosis|DIAGNOSES
Disorder|Disease or Syndrome|Hospital Course|12906,12912|false|false|false|C0002871|Anemia|anemia
Event|Event|Hospital Course|12906,12912|false|false|false|||anemia
Finding|Intellectual Product|Hospital Course|12916,12921|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|Hospital Course|12916,12934|false|false|false|C0333361|Acute inflammation|acute inflammation
Event|Event|Hospital Course|12922,12934|false|false|false|||inflammation
Finding|Pathologic Function|Hospital Course|12922,12934|false|false|false|C0021368|Inflammation|inflammation
Disorder|Disease or Syndrome|Hospital Course|12937,12940|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12937,12940|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|12937,12940|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|12937,12940|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|12937,12940|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|12937,12940|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|12937,12940|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12937,12940|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|Hospital Course|12950,12957|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|12950,12957|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|12950,12957|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|12950,12970|false|false|false|C1135194|Chronic systolic heart failure|chronic systolic CHF
Finding|Organ or Tissue Function|Hospital Course|12958,12966|false|false|false|C0039155|Systole|systolic
Disorder|Disease or Syndrome|Hospital Course|12958,12970|false|false|false|C2039715|systolic congestive heart failure|systolic CHF
Anatomy|Body Space or Junction|Hospital Course|12967,12970|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|12967,12970|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|12967,12970|false|false|false|||CHF
Disorder|Disease or Syndrome|Hospital Course|12973,12976|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|12973,12976|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|12979,12982|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Hospital Course|12983,12988|false|false|false|C1300072|Tumor stage|stage
Finding|Mental Process|Discharge Condition|13017,13023|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|13017,13030|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|13017,13030|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|13024,13030|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|13024,13030|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|13032,13037|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|13032,13037|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|13042,13050|false|false|false|||coherent
Finding|Finding|Discharge Condition|13042,13050|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|13052,13057|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|13052,13074|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|13052,13074|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|13061,13074|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|13061,13074|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|13061,13074|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|13076,13081|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|13076,13081|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|13076,13081|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|13076,13081|false|false|false|||Alert
Finding|Finding|Discharge Condition|13076,13081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|13076,13081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|13076,13081|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|13086,13097|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|13086,13097|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|13099,13107|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|13099,13107|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|13099,13107|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|13108,13114|false|false|false|C5889824||Status
Event|Event|Discharge Condition|13108,13114|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|13108,13114|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|13116,13126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|13116,13126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|13116,13126|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|13116,13126|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|13129,13137|false|false|false|||requires
Event|Event|Discharge Condition|13138,13148|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|13138,13148|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|13152,13155|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|13152,13155|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|13152,13155|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|13152,13155|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|13152,13155|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|13157,13163|false|false|false|||walker
Event|Event|Discharge Instructions|13211,13219|false|false|false|||admitted
Drug|Organic Chemical|Discharge Instructions|13225,13230|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Discharge Instructions|13225,13230|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Discharge Instructions|13225,13230|false|false|false|||cough
Finding|Sign or Symptom|Discharge Instructions|13225,13230|false|false|false|C0010200|Coughing|cough
Event|Event|Discharge Instructions|13235,13240|false|false|false|||found
Finding|Finding|Discharge Instructions|13249,13252|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|13249,13252|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Biologically Active Substance|Discharge Instructions|13253,13259|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|13253,13259|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|13253,13259|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13253,13259|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Instructions|13260,13266|false|false|false|||levels
Event|Event|Discharge Instructions|13274,13282|false|false|false|||required
Procedure|Health Care Activity|Discharge Instructions|13287,13301|false|false|false|C0085559|intensive care|Intensive Care
Finding|Idea or Concept|Discharge Instructions|13287,13306|false|false|false|C1549475|Room type - Intensive care unit|Intensive Care Unit
Event|Activity|Discharge Instructions|13297,13301|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|13297,13301|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|13297,13301|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Discharge Instructions|13316,13321|false|false|false|||shows
Event|Event|Discharge Instructions|13323,13334|false|false|false|||progression
Finding|Functional Concept|Discharge Instructions|13323,13334|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Discharge Instructions|13323,13334|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Anatomy|Body Location or Region|Discharge Instructions|13343,13347|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13343,13347|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|13343,13347|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|13343,13347|false|false|false|C0740941|Lung Problem|lung
Disorder|Neoplastic Process|Discharge Instructions|13343,13354|false|false|false|C0242379;C0684249|Carcinoma of lung;Malignant neoplasm of lung|lung cancer
Disorder|Neoplastic Process|Discharge Instructions|13348,13354|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Discharge Instructions|13348,13354|false|false|false|||cancer
Finding|Finding|Discharge Instructions|13362,13370|false|false|false|C0332148|Probable diagnosis|probable
Event|Event|Discharge Instructions|13371,13383|false|false|false|||superimposed
Disorder|Disease or Syndrome|Discharge Instructions|13385,13394|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|Discharge Instructions|13385,13394|false|false|false|||pneumonia
Event|Event|Discharge Instructions|13405,13412|false|false|false|||treated
Drug|Antibiotic|Discharge Instructions|13418,13429|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|13418,13429|false|false|false|||antibiotics
Drug|Biologically Active Substance|Discharge Instructions|13434,13440|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|13434,13440|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|13434,13440|false|false|false|C0030054|oxygen|oxygen
Event|Event|Discharge Instructions|13434,13440|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13434,13440|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Instructions|13446,13454|false|false|false|||improved
Event|Event|Discharge Instructions|13469,13479|false|false|false|||tranferred
Finding|Functional Concept|Discharge Instructions|13487,13494|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|13487,13494|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|13487,13494|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|13487,13494|false|false|false|C0199168|Medical service|medical
Anatomy|Anatomical Structure|Discharge Instructions|13495,13500|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Discharge Instructions|13512,13521|false|false|false|||continued
Drug|Antibiotic|Discharge Instructions|13525,13536|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|13525,13536|false|false|false|||antibiotics
Drug|Biologically Active Substance|Discharge Instructions|13547,13553|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|13547,13553|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|13547,13553|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13547,13553|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Event|Event|Discharge Instructions|13554,13560|false|false|false|||levels
Event|Event|Discharge Instructions|13566,13575|false|false|false|||monitored
Event|Event|Discharge Instructions|13589,13601|false|false|false|||communicated
Event|Event|Discharge Instructions|13651,13656|false|false|false|||weigh
Event|Event|Discharge Instructions|13661,13666|false|false|false|||risks
Finding|Idea or Concept|Discharge Instructions|13661,13666|false|false|false|C0035647|Risk|risks
Event|Event|Discharge Instructions|13671,13679|false|false|false|||benefits
Finding|Functional Concept|Discharge Instructions|13684,13694|false|false|false|C1524062|Additional|additional
Event|Event|Discharge Instructions|13695,13707|false|false|false|||chemotherapy
Finding|Functional Concept|Discharge Instructions|13695,13707|false|false|false|C0013217|pharmacotherapeutic|chemotherapy
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13695,13707|false|false|false|C0013216;C0392920;C3665472|Chemotherapy;Chemotherapy Regimen;Pharmacotherapy|chemotherapy
Event|Event|Discharge Instructions|13723,13734|false|false|false|||complicated
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13744,13750|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Discharge Instructions|13744,13750|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|Discharge Instructions|13744,13750|false|false|false|||kidney
Finding|Sign or Symptom|Discharge Instructions|13744,13750|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Discharge Instructions|13744,13750|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13744,13750|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Finding|Pathologic Function|Discharge Instructions|13744,13762|false|false|false|C0151746|Abnormal renal function|kidney dysfunction
Disorder|Disease or Syndrome|Discharge Instructions|13751,13762|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|Discharge Instructions|13751,13762|false|false|false|||dysfunction
Finding|Conceptual Entity|Discharge Instructions|13751,13762|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Discharge Instructions|13751,13762|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|Discharge Instructions|13751,13762|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|Discharge Instructions|13773,13780|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|13773,13780|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|13773,13780|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|13773,13780|false|false|false|C0199168|Medical service|medical
Event|Event|Discharge Instructions|13781,13789|false|false|false|||problems
Finding|Idea or Concept|Discharge Instructions|13781,13789|false|false|false|C1546466|Problems - What subject filter|problems
Event|Event|Discharge Instructions|13794,13799|false|false|false|||plans
Procedure|Diagnostic Procedure|Discharge Instructions|13816,13823|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|Discharge Instructions|13819,13823|false|false|false|||scan
Procedure|Diagnostic Procedure|Discharge Instructions|13819,13823|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|Discharge Instructions|13833,13839|false|false|false|||finish
Drug|Antibiotic|Discharge Instructions|13845,13856|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|Discharge Instructions|13845,13856|false|false|false|||antibiotics
Event|Event|Discharge Instructions|13869,13877|false|false|false|||evaluate
Event|Activity|Discharge Instructions|13882,13886|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|13882,13886|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|13882,13886|false|false|false|C1549480|Amount type - Rate|rate
Disorder|Disease or Syndrome|Discharge Instructions|13895,13902|false|false|false|C0012634|Disease|disease
Event|Event|Discharge Instructions|13895,13902|false|false|false|||disease
Finding|Pathologic Function|Discharge Instructions|13895,13914|false|false|false|C0242656|Disease Progression|disease progression
Event|Event|Discharge Instructions|13903,13914|false|false|false|||progression
Finding|Functional Concept|Discharge Instructions|13903,13914|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Finding|Pathologic Function|Discharge Instructions|13903,13914|false|false|false|C0242656;C0449258|Disease Progression;Progression|progression
Disorder|Disease or Syndrome|Discharge Instructions|13922,13946|false|false|false|C0018802|Congestive heart failure|congestive heart failure
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13933,13938|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|13933,13938|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|13933,13938|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|13933,13946|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|heart failure
Event|Event|Discharge Instructions|13939,13946|false|false|false|||failure
Finding|Functional Concept|Discharge Instructions|13939,13946|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Discharge Instructions|13939,13946|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Discharge Instructions|13939,13946|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Event|Event|Discharge Instructions|13956,13962|false|false|false|||stable
Finding|Intellectual Product|Discharge Instructions|13956,13962|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Discharge Instructions|13971,13975|false|false|false|||note
Event|Event|Discharge Instructions|13980,13987|false|false|false|||stopped
Drug|Organic Chemical|Discharge Instructions|13993,13998|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Discharge Instructions|13993,13998|false|false|false|C0699992|Lasix|lasix
Event|Event|Discharge Instructions|13993,13998|false|false|false|||lasix
Drug|Organic Chemical|Discharge Instructions|14003,14013|false|false|false|C0051696|amlodipine|amlodipine
Drug|Pharmacologic Substance|Discharge Instructions|14003,14013|false|false|false|C0051696|amlodipine|amlodipine
Event|Event|Discharge Instructions|14003,14013|false|false|false|||amlodipine
Event|Event|Discharge Instructions|14036,14040|false|false|false|||need
Event|Event|Discharge Instructions|14048,14060|false|false|false|||re-evaluated
Disorder|Disease or Syndrome|Discharge Instructions|14069,14072|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|14069,14072|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|14069,14072|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|14069,14072|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|14069,14072|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|14069,14072|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|14069,14072|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|14069,14072|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Discharge Instructions|14069,14072|false|false|false|||PCP
Finding|Gene or Genome|Discharge Instructions|14069,14072|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|14069,14072|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Discharge Instructions|14076,14079|false|false|false|||see
Event|Event|Discharge Instructions|14096,14103|false|false|false|||restart
Event|Event|Discharge Instructions|14119,14128|false|false|false|||decreased
Event|Event|Discharge Instructions|14142,14146|false|false|false|||dose
Drug|Organic Chemical|Discharge Instructions|14150,14160|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Discharge Instructions|14150,14160|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|Discharge Instructions|14150,14160|false|false|false|||metoprolol
Event|Event|Discharge Instructions|14180,14185|false|false|false|||weigh
Finding|Functional Concept|Discharge Instructions|14214,14218|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Gene or Genome|Discharge Instructions|14214,14218|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Intellectual Product|Discharge Instructions|14214,14218|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Finding|Mental Process|Discharge Instructions|14214,14218|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|call
Attribute|Clinical Attribute|Discharge Instructions|14225,14231|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|14225,14231|false|false|false|||weight
Finding|Finding|Discharge Instructions|14225,14231|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|14225,14231|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|14225,14231|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|14232,14236|false|false|false|||goes
Procedure|Laboratory Procedure|Discharge Instructions|14253,14256|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Procedure|Health Care Activity|Discharge Instructions|14260,14268|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|14269,14281|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|14269,14281|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|14269,14281|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

