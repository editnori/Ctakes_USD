CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|penicillins|Drug|false|false||Penicillins
null|penicillins|Drug|false|false||Penicillinsnull|Poisoning by, adverse effect of and underdosing of penicillins|Disorder|false|false||Penicillins
null|Poisoning by penicillin|Disorder|false|false||Penicillinsnull|Adverse reaction to penicillins|Finding|false|false||Penicillinsnull|Dilantin|Drug|false|false||Dilantin
null|Dilantin|Drug|false|false||Dilantinnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|true|false||History of Present Illnessnull|null|Attribute|true|false||History of Present Illnessnull|Medical History|Finding|true|false||History ofnull|History of present illness (finding)|Finding|true|false||History
null|History of previous events|Finding|true|false||History
null|Historical aspects qualifier|Finding|true|false||History
null|Medical History|Finding|true|false||History
null|Concept History|Finding|true|false||Historynull|History|Subject|true|false||Historynull|Present illness|Finding|true|false||Present Illnessnull|Present|Finding|true|false||Present
null|Presentation|Finding|true|false||Presentnull|Illness (finding)|Finding|true|false||Illnessnull|Medical History|Finding|false|false||medical historynull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Medical History|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|History of present illness (finding)|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Irritable Bowel Syndrome|Disorder|false|false||irritable bowel syndromenull|Irritable Bowel Syndrome|Disorder|false|false||irritable bowelnull|Irritable Mood|Finding|false|false||irritable
null|Irritability - emotion|Finding|false|false||irritablenull|Intestines|Anatomy|false|false||bowelnull|Syndrome|Disorder|false|false||syndromenull|Presenile dementia|Disorder|false|false||dementia
null|Dementia|Disorder|false|false||dementianull|Problems - What subject filter|Finding|true|false||problemsnull|Intestines|Anatomy|true|false||bowelsnull|year|Time|true|false||yearsnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||acute onsetnull|Sudden onset (attribute)|Time|false|false||acute onset
null|acute|Time|false|false||acute onsetnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onset ofnull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Morning|Time|false|false||morningnull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Event|Event|false|false||eventnull|Recent|Time|true|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Illness (finding)|Finding|true|false||sicknull|Contacts|Procedure|true|false||contactsnull|Corned beef|Drug|false|false||corned beefnull|beef allergenic extract|Drug|false|false||beef
null|Beef preparation|Drug|false|false||beef
null|Beef preparation|Drug|false|false||beef
null|beef allergenic extract|Drug|false|false||beef
null|Beef (dietary)|Drug|false|false||beef
null|Beef Antigen|Drug|false|false||beefnull|Cattle for beef production|Entity|false|false||beefnull|cabbage allergenic extract|Drug|false|false||cabbage
null|cabbage preparation|Drug|false|false||cabbage
null|cabbage preparation|Drug|false|false||cabbage
null|null|Drug|false|false||cabbage
null|cabbage allergenic extract|Drug|false|false||cabbagenull|Brassica oleracea|Entity|false|false||cabbagenull|Local Remote Control State - Local|Finding|false|false||localnull|Local|Modifier|false|false||localnull|Last|Modifier|false|false||lastnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Loose|Modifier|false|false||loosenull|Watery diarrhoea|Finding|false|false||watery diarrheanull|Watery|Modifier|false|false||waterynull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Abdominal Cramps|Finding|true|false||abdominal crampingnull|Abdomen|Anatomy|true|false||abdominalnull|Abdominal (qualifier value)|Modifier|true|false||abdominalnull|Muscle Cramp|Finding|true|false||crampingnull|Cramping sensation quality|Modifier|true|false||crampingnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|rectal discharge diarrhea (physical finding)|Finding|true|false||diarrhea
null|Diarrhea|Finding|true|false||diarrheanull|Imodium|Drug|true|false||Imodium
null|Imodium|Drug|true|false||Imodiumnull|Unable|Finding|false|false||unablenull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Food|Drug|false|false||foodsnull|Presentation|Finding|false|false||presentednull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|White Blood Cell Count procedure|Procedure|false|false||WBC countnull|Leukocytes|Anatomy|false|false||WBCnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Blood urea increased|Finding|false|false||elevated BUNnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|liter|LabModifier|false|false||liternull|Saline Solution|Drug|false|false||saline
null|Saline Solution|Drug|false|false||salinenull|Saline method|Procedure|false|false||salinenull|Review of systems (procedure)|Procedure|false|false||Review of Systemsnull|null|Attribute|false|false||Review of Systems
null|null|Attribute|false|false||Review of Systemsnull|Review of|Finding|false|false||Review ofnull|Review (Publication Type)|Finding|false|false||Review
null|Act Class - review|Finding|false|false||Reviewnull|System|Finding|false|false||Systemsnull|Pain Measurement|Procedure|false|false||Pain assessmentnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Knowledge acquisition using a method of assessment|Finding|false|false||assessmentnull|assessment of cognitive functions|Procedure|false|false||assessment
null|Physical Examination|Procedure|false|false||assessment
null|Nutrition Assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Personal care assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Evaluation procedure|Procedure|false|false||assessment
null|Evaluation|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessmentnull|Assessed|Event|false|false||assessmentnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Recent|Time|true|false||recentnull|Illness (finding)|Finding|true|false||illnessesnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Night time|Time|true|false||nightnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Dyspnea|Finding|true|false||SOBnull|Cough (guaifenesin)|Drug|true|false||cough
null|Cough (guaifenesin)|Drug|true|false||coughnull|Coughing|Finding|true|false||coughnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Urinary symptoms|Finding|true|false||urinary symptomsnull|Urinary tract|Anatomy|true|false||urinarynull|urinary|Modifier|true|false||urinarynull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|System|Finding|false|false||systemsnull|detail - Response Level|Finding|false|false||detailnull|Details|Modifier|false|false||detailnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|Osteoporosis|Disorder|false|false||Osteoporosisnull|Encounter due to family history of osteoporosis|Finding|false|false||Osteoporosisnull|Irritable Bowel Syndrome|Disorder|false|false||Irritable bowel syndromenull|Irritable Bowel Syndrome|Disorder|false|false||Irritable bowelnull|Irritable Mood|Finding|false|false||Irritable
null|Irritability - emotion|Finding|false|false||Irritablenull|Intestines|Anatomy|false|false||bowelnull|Syndrome|Disorder|false|false||syndromenull|Macrocytosis (morphologic abnormality)|Disorder|false|false||Macrocytosis
null|Macrocytosis|Disorder|false|false||Macrocytosisnull|Macrocytosis (finding)|Lab|false|false||Macrocytosisnull|Science of Etiology|Finding|false|false||etiology
null|Etiology aspects|Finding|false|false||etiology
null|Etiology|Finding|false|false||etiologynull|left ear symptoms (symptom)|Finding|false|false||Left earnull|Left ear structure|Anatomy|false|false||Left earnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Ear and labyrinth disorders|Disorder|false|false||earnull|SpecimenType - Ear|Finding|false|false||ear
null|null|Finding|false|false||earnull|Ear structure|Anatomy|false|false||ear
null|null|Anatomy|false|false||earnull|hearing impairment|Disorder|false|false||hearing lossnull|hearing loss by exam|Finding|false|false||hearing loss
null|Partial Hearing Loss|Finding|false|false||hearing loss
null|Hearing Loss|Finding|false|false||hearing loss
null|Deafness|Finding|false|false||hearing lossnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Appendectomy; for ruptured appendix with abscess or generalized peritonitis|Procedure|false|false||appendectomy
null|Appendectomy|Procedure|false|false||appendectomynull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Removal of ovarian cyst|Procedure|false|false||ovarian cyst removalnull|Ovarian Cysts|Disorder|false|false||ovarian cystnull|Ovarian|Anatomy|false|false||ovariannull|Cyst removal|Procedure|false|false||cyst removalnull|Cyst|Disorder|false|false||cystnull|SpecimenType - Cyst|Finding|false|false||cyst
null|null|Finding|false|false||cystnull|Cyst form of protozoa|Entity|false|false||cystnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|reported history of cataract surgery|Finding|false|false||Cataract surgery
null|Consent Type - Cataract Surgery|Finding|false|false||Cataract surgerynull|Cataract surgery|Procedure|false|false||Cataract surgery
null|Cataract Extraction|Procedure|false|false||Cataract surgerynull|Cataract surgery specialty (qualifier value)|Title|false|false||Cataract surgerynull|Cataract|Disorder|false|false||Cataractnull|cataract on exam (physical finding)|Finding|false|false||Cataractnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Glaucoma|Disorder|false|false||Glaucomanull|Glaucoma <Glaucomidae>|Entity|false|false||Glaucomanull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Relevance|Modifier|true|false||relevantnull|Electrical Current|Phenomenon|true|false||currentnull|Current (present time)|Time|true|false||currentnull|Admission activity|Procedure|true|false||admission
null|Hospital admission|Procedure|true|false||admissionnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Taking vital signs|Procedure|false|false||Vital Signsnull|null|Attribute|false|false||Vital Signs
null|Vital signs|Attribute|false|false||Vital Signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||Signs
null|Physical findings|Finding|false|false||Signsnull|Manufactured sign|Device|false|false||Signsnull|physical examination (physical finding)|Finding|false|false||Physical examinationnull|Physical Examination|Procedure|false|false||Physical examinationnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Physical Examination|Procedure|false|false||examination
null|Medical Examination|Procedure|false|false||examinationnull|Examination|Event|false|false||examinationnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Elderly (population group)|Subject|false|false||Elderlynull|Old age|Time|false|false||Elderlynull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|hearing impairment|Disorder|false|false||Hard of hearingnull|Partial Hearing Loss|Finding|false|false||Hard of hearingnull|Hardness|Modifier|false|false||Hardnull|outcomes otolaryngology hearing|Finding|false|false||hearing
null|Hearing finding|Finding|false|false||hearing
null|Hearing|Finding|false|false||hearingnull|right ear symptoms (symptom)|Finding|false|false||Right earnull|Right ear structure|Anatomy|false|false||Right earnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Ear and labyrinth disorders|Disorder|false|false||earnull|SpecimenType - Ear|Finding|false|false||ear
null|null|Finding|false|false||earnull|Ear structure|Anatomy|false|false||ear
null|null|Anatomy|false|false||earnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Respiration|Finding|false|false||respirationsnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Auscultation|Procedure|false|false||auscultationnull|Regular|Modifier|false|false||Regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Jugular venous pressure|Finding|false|false||JVPnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Ankle edema (finding)|Finding|true|false||ankle edemanull|Lower extremity>Ankle|Anatomy|true|false||ankle
null|Ankle|Anatomy|true|false||ankle
null|Ankle joint structure|Anatomy|true|false||anklenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Daughter|Subject|false|false||daughternull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|Timing, LOINC Axis 3|Finding|true|false||timingnull|Timing|Time|true|false||timingnull|recent events relating to health|Finding|false|false||recent eventsnull|Recent|Time|false|false||recentnull|Event|Event|false|false||eventsnull|Poor short-term memory|Disorder|false|false||short-term memory impairmentnull|Memory, Short-Term|Finding|false|false||short-term memorynull|short-term|Time|false|false||short-termnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Term (lexical)|Finding|false|false||term
null|Term Birth|Finding|false|false||termnull|Term (temporal)|Time|false|false||termnull|Memory impairment|Disorder|false|false||memory impairmentnull|Forgetful|Finding|false|false||memory impairmentnull|Memory observations|Finding|false|false||memory
null|Memory G-code|Finding|false|false||memory
null|Memory|Finding|false|false||memorynull|Memory Device|Device|false|false||memorynull|Impaired health|Finding|false|false||impairment
null|Impaired|Finding|false|false||impairmentnull|Speech|Finding|false|false||Speechnull|Speech assessment|Procedure|false|false||Speechnull|Programming Languages|Finding|false|false||languagenull|null|Attribute|false|false||languagenull|Languages|Entity|false|false||languagenull|Psychiatric problem|Disorder|false|false||Psych
null|Mental disorders|Disorder|false|false||Psychnull|patient appearance regarding mental status exam|Procedure|false|false||Appearancenull|null|Attribute|false|false||Appearancenull|Personal appearance|Subject|false|false||Appearancenull|Appearance|Modifier|false|false||Appearancenull|Kind of quantity - Appearance|LabModifier|false|false||Appearancenull|Behavior|Finding|false|false||behaviornull|null|Attribute|false|false||behaviornull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Laboratory test finding|Lab|false|false||Labsnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Bands|Device|false|false||Bandsnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipase
null|lipase|Drug|false|false||Lipasenull|Lipase measurement|Procedure|false|false||Lipasenull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Yellow color|Modifier|false|false||Yellownull|Cloudy|Modifier|false|false||Hazynull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Leukocytes|Anatomy|false|false||WBCnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|true|false||MODnull|Yeast, Dried|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeast
null|Candida albicans allergenic extract|Drug|true|false||Yeastnull|Saccharomyces cerevisiae|Entity|true|false||Yeast
null|Yeasts|Entity|true|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|epinephrine|Drug|true|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|true|false||Epinull|Exocrine pancreatic insufficiency|Disorder|true|false||Epinull|Eysenck personality inventory|Finding|true|false||Epi
null|TFPI wt Allele|Finding|true|false||Epi
null|TFPI gene|Finding|true|false||Epinull|Electronic Portal Imaging|Procedure|true|false||Epi
null|Echo-Planar Imaging|Procedure|true|false||Epinull|Microbiology Diagnostic Service Section ID|Finding|false|false||Microbiology
null|Microbiological|Finding|false|false||Microbiology
null|Microbiology - Laboratory Class|Finding|false|false||Microbiologynull|Microbiology procedure|Procedure|false|false||Microbiologynull|Science of Microbiology|Title|false|false||Microbiologynull|Feces|Finding|false|false||Stoolnull|Stool seat|Device|false|false||Stoolnull|Culture (Anthropological)|Finding|false|false||Culturesnull|Consistency of stool|Finding|false|false||STOOL     CONSISTENCYnull|Feces|Finding|false|false||STOOLnull|Stool seat|Device|false|false||STOOLnull|Consistency|Modifier|false|false||CONSISTENCYnull|Kind of quantity - Consistency|LabModifier|false|false||CONSISTENCYnull|Watery|Modifier|false|false||WATERYnull|Source (property) (qualifier value)|Finding|false|false||Source
null|Term Source|Finding|false|false||Source
null|Source|Finding|false|false||Sourcenull|Feces|Finding|false|false||Stoolnull|Stool seat|Device|false|false||Stoolnull|Stool culture|Procedure|false|false||FECAL CULTUREnull|Feces|Finding|false|false||FECALnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Pending - Allergy Clinical Status|Finding|false|false||Pending
null|Pending - referral status|Finding|false|false||Pendingnull|Pending - status|Time|false|false||Pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||Pending
null|pending - RoleStatus|Modifier|false|false||Pending
null|Pending - Day type|Modifier|false|false||Pendingnull|Campylobacter culture|Procedure|false|false||CAMPYLOBACTER CULTUREnull|Campylobacter|Entity|false|false||CAMPYLOBACTERnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Pending - Allergy Clinical Status|Finding|false|false||Pending
null|Pending - referral status|Finding|false|false||Pendingnull|Pending - status|Time|false|false||Pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||Pending
null|pending - RoleStatus|Modifier|false|false||Pending
null|Pending - Day type|Modifier|false|false||Pendingnull|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN A
null|tcdA protein, Clostridium difficile|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN Anull|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXIN
null|Clostridium difficile toxin|Drug|false|false||CLOSTRIDIUM DIFFICILE TOXINnull|Clostridioides difficile|Entity|false|false||CLOSTRIDIUM DIFFICILEnull|Genus Clostridium (organism)|Entity|false|false||CLOSTRIDIUMnull|Toxin|Drug|false|false||TOXIN
null|Toxin|Drug|false|false||TOXINnull|Toxin (disposition)|Modifier|false|false||TOXINnull|Tests (qualifier value)|Finding|false|false||TEST
null|Testing|Finding|false|false||TESTnull|Laboratory Procedures|Procedure|false|false||TESTnull|Test - temporal region|Anatomy|false|false||TESTnull|Test Result|Lab|false|false||TESTnull|Test Dosing Unit|LabModifier|false|false||TESTnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Feces|Finding|true|false||Fecesnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Toxin|Drug|false|false||toxin
null|Toxin|Drug|false|false||toxinnull|Toxin (disposition)|Modifier|false|false||toxinnull|Endocrine Therapy-Induced Alopecia|Disorder|false|false||EIA
null|Equine Infectious Anemia|Disorder|false|false||EIAnull|Enzyme Immunoassay|Procedure|false|false||EIAnull|Reference range (qualifier value)|Modifier|false|false||Reference Rangenull|null|LabModifier|false|false||Reference Rangenull|Reference - MdfHmdMetSourceType|Finding|false|false||Reference
null|Reference Object|Finding|false|false||Reference
null|Reference source|Finding|false|false||Reference
null|Bibliographic Reference|Finding|false|false||Reference
null|Reference - HL7UpdateMode|Finding|false|false||Referencenull|Concept model range (foundation metadata concept)|Finding|false|false||Rangenull|Sample Range|LabModifier|false|false||Range
null|Range|LabModifier|false|false||Rangenull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Culture (Anthropological)|Finding|false|false||Culturesnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Ichthyosis Bullosa of Siemens|Disorder|false|false||IBS
null|Irritable Bowel Syndrome|Disorder|false|false||IBSnull|Presenile dementia|Disorder|false|false||Dementia
null|Dementia|Disorder|false|false||Dementianull|day|Time|false|false||daysnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Dehydration|Disorder|false|false||dehydratednull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Kidney Failure, Acute|Disorder|false|false||acute renal failurenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Kidney Failure|Disorder|false|false||renal failurenull|Urologic Diseases|Disorder|false|false||renalnull|Kidney|Anatomy|false|false||renalnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Symptomatic|Finding|false|false||symptomaticnull|Orthostasis|Finding|false|false||orthostasis
null|Orthostatic intolerance|Finding|false|false||orthostasisnull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false||IVFnull|SCN5A wt Allele|Finding|false|false||IVF
null|SCN5A gene|Finding|false|false||IVFnull|Assisted Reproductive Technologies|Procedure|false|false||IVF
null|Fertilization in Vitro|Procedure|false|false||IVFnull|Structure of interventricular foramen|Anatomy|false|false||IVFnull|Intestines|Anatomy|false|false||bowelnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Presentation|Finding|false|false||presentationnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Slow|Modifier|false|false||slowlynull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Renal function|Finding|false|false||Renal functionnull|Kidney Function Tests|Procedure|false|false||Renal functionnull|Urologic Diseases|Disorder|false|false||Renalnull|Kidney|Anatomy|false|false||Renalnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Ventricular Fibrillation, Paroxysmal Familial, 1|Disorder|false|false||IVFnull|SCN5A wt Allele|Finding|false|false||IVF
null|SCN5A gene|Finding|false|false||IVFnull|Assisted Reproductive Technologies|Procedure|false|false||IVF
null|Fertilization in Vitro|Procedure|false|false||IVFnull|Structure of interventricular foramen|Anatomy|false|false||IVFnull|Bland diet|Finding|true|false||bland dietnull|Diet (animal life circumstance)|Drug|true|false||diet
null|Diet|Drug|true|false||dietnull|diet - supply|Finding|true|false||dietnull|Diet therapy|Procedure|true|false||dietnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Orthostasis|Finding|true|false||orthostasis
null|Orthostatic intolerance|Finding|true|false||orthostasisnull|Transaction counts and value totals - day|Finding|true|false||day
null|Precision - day|Finding|true|false||daynull|Land Dayak Languages|Entity|true|false||daynull|day|Time|true|false||day
null|Daily|Time|true|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|SAFE-Biopharma Standard|Finding|true|false||safenull|Discharge to home|Procedure|true|false||discharge homenull|Body Substance Discharge|Finding|true|false||discharge
null|Discharge Body Fluid|Finding|true|false||discharge
null|Body Fluid Discharge|Finding|true|false||discharge
null|null|Finding|true|false||dischargenull|Patient Discharge|Procedure|true|false||dischargenull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|Clinical Service|Procedure|true|false||servicesnull|Services|Event|true|false||servicesnull|Conjunctivitis|Disorder|false|false||Conjunctivitisnull|examination of left eye|Procedure|false|false||left eyenull|Left eye structure|Anatomy|false|false||left eyenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Drops - Drug Form|Drug|false|false||dropsnull|Drop Dosing Unit|LabModifier|false|false||dropsnull|examination of left eye|Procedure|false|false||left eyenull|Left eye structure|Anatomy|false|false||left eyenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Conjunctivitis|Disorder|false|false||conjunctivitisnull|Continuous|Finding|false|false||ongoingnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|Ointments|Drug|false|false||ointmentnull|Improvement|Finding|false|false||improvementnull|Conjunctival hyperemia|Finding|false|false||conjunctival injectionnull|Conjunctival Route of Administration|Finding|false|false||conjunctivalnull|conjunctiva|Anatomy|false|false||conjunctivalnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Eye symptom|Finding|true|false||eye symptomsnull|Carcinoma in situ of eye|Disorder|true|false||eye
null|Disorder of eye|Disorder|true|false||eyenull|Eye - Specimen Source Code|Finding|true|false||eye
null|Eye problem|Finding|true|false||eye
null|Eye Specimen|Finding|true|false||eyenull|Head>Eye|Anatomy|true|false||eye
null|Eye|Anatomy|true|false||eye
null|Orbital region|Anatomy|true|false||eyenull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Chronic - Admission Level of Care Code|Finding|true|false||chronicnull|Provision of recurring care for chronic illness|Procedure|true|false||chronicnull|chronic|Time|true|false||chronicnull|Pharmaceutical Preparations|Drug|true|false||medicationnull|medication - HL7 publishing domain|Finding|true|false||medication
null|Medications|Finding|true|false||medicationnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|CODE STATUS|Procedure|false|false||Code Statusnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|daunorubicin|Drug|false|false||DNR
null|daunorubicin|Drug|false|false||DNRnull|Do-Not-Resuscitate Orders|Finding|false|false||DNR
null|Do not resuscitate status|Finding|false|false||DNRnull|null|Attribute|false|false||DNRnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Primary caregiver|Subject|false|false||primary caregivernull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Caregiver|Subject|false|false||caregivernull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Daily|Time|false|false||dailynull|Namenda|Drug|false|false||Namenda
null|Namenda|Drug|false|false||Namendanull|Daily|Time|false|false||dailynull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||dailynull|raloxifene|Drug|false|false||Raloxifene
null|raloxifene|Drug|false|false||Raloxifenenull|Evista|Drug|false|false||Evista
null|Evista|Drug|false|false||Evistanull|Daily|Time|false|false||dailynull|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitamin
null|Multivitamin preparation|Drug|false|false||Multivitaminnull|Daily|Time|false|false||dailynull|glucosamine|Drug|false|false||Glucosamine
null|glucosamine|Drug|false|false||Glucosaminenull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium supplement
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium supplementnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Dietary Supplements|Drug|false|false||supplementnull|Supplement - Diet Code Specification Type|Finding|false|false||supplement
null|Supplement|Finding|false|false||supplement
null|Supplement (document)|Finding|false|false||supplementnull|cholecalciferol|Drug|false|false||Cholecalciferol (Vitamin D3)
null|cholecalciferol|Drug|false|false||Cholecalciferol (Vitamin D3)
null|cholecalciferol|Drug|false|false||Cholecalciferol (Vitamin D3)null|cholecalciferol|Drug|false|false||Cholecalciferol
null|cholecalciferol|Drug|false|false||Cholecalciferol
null|cholecalciferol|Drug|false|false||Cholecalciferolnull|vitamin D3|Drug|false|false||Vitamin D3
null|vitamin D3|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3
null|cholecalciferol|Drug|false|false||Vitamin D3null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Daily|Time|false|false||dailynull|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acid
null|ascorbic acid|Drug|false|false||Ascorbic Acidnull|Ascorbic acid measurement|Procedure|false|false||Ascorbic Acidnull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|donepezil|Drug|false|false||donepezil
null|donepezil|Drug|false|false||donepezilnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Namenda|Drug|false|false||Namenda
null|Namenda|Drug|false|false||Namendanull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||qhsnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Delayed Release Dosage Form|Drug|false|false||Delayed Releasenull|Views delayed|Attribute|false|false||Delayednull|Deferred|Time|false|false||Delayednull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|raloxifene|Drug|false|false||raloxifene
null|raloxifene|Drug|false|false||raloxifenenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a week|Time|false|false||once a weeknull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitamin
null|Multivitamin preparation|Drug|false|false||multivitaminnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|glucosamine|Drug|false|false||Glucosamine
null|glucosamine|Drug|false|false||Glucosaminenull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|ascorbic acid|Drug|false|false||ascorbic acid
null|ascorbic acid|Drug|false|false||ascorbic acid
null|ascorbic acid|Drug|false|false||ascorbic acidnull|Ascorbic acid measurement|Procedure|false|false||ascorbic acidnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Oral Dosage Form|Drug|false|false||Oralnull|Oral Route of Administration|Finding|false|false||Oral
null|Oral (intended site)|Finding|false|false||Oralnull|Oral cavity|Anatomy|false|false||Oralnull|Oral|Modifier|false|false||Oralnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|gram|LabModifier|false|false||gramnull|Ointments|Drug|false|false||Ointmentnull|Inch Unit of Length|LabModifier|false|false||inchnull|Ophthalmic Dosage Form|Drug|false|false||Ophthalmicnull|Ophthalmic Route of Administration|Finding|false|false||Ophthalmicnull|Eye|Anatomy|false|false||Ophthalmicnull|Four times daily|Time|false|false||four times a daynull|Four Times|LabModifier|false|false||four timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|examination of left eye|Procedure|false|false||left eyenull|Left eye structure|Anatomy|false|false||left eyenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|refill|Finding|false|false||Refillsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Gastrointestinal attachment|Finding|false|false||Gastrointestinalnull|gastrointestinal|Modifier|false|false||Gastrointestinalnull|Virus Diseases|Disorder|false|false||Virus
null|AS virus|Disorder|false|false||Virus
null|Virus|Disorder|false|false||Virusnull|dehydration (Na, H2O)|Disorder|false|false||Dehydration
null|Dehydration|Disorder|false|false||Dehydrationnull|Dehydration procedure|Procedure|false|false||Dehydrationnull|Symptomatic|Finding|false|false||Symptomaticnull|Orthostasis|Finding|false|false||orthostasis
null|Orthostatic intolerance|Finding|false|false||orthostasisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Illness (finding)|Finding|false|false||illnessnull|dehydration (Na, H2O)|Disorder|false|false||dehydration
null|Dehydration|Disorder|false|false||dehydrationnull|Dehydration procedure|Procedure|false|false||dehydrationnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Virus Diseases|Disorder|false|false||virus
null|AS virus|Disorder|false|false||virus
null|Virus|Disorder|false|false||virusnull|Very|Modifier|false|false||verynull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Supportive assistance|Finding|false|false||supportivenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Improvement|Finding|false|false||improvementnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|SAFE-Biopharma Standard|Finding|false|false||safenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Much|Finding|false|false||muchnull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Hydration status|Finding|false|false||hydration
null|Hydration|Finding|false|false||hydrationnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Appointments|Event|false|false||appointmentnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|examination of left eye|Procedure|false|false||left eyenull|Left eye structure|Anatomy|false|false||left eyenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Conjunctivitis|Disorder|false|false||conjunctivitisnull|null|Drug|false|false||erythromycin ointmentnull|erythromycin|Drug|false|false||erythromycin
null|erythromycin|Drug|false|false||erythromycinnull|Ointments|Drug|false|false||ointmentnull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|true|false||facenull|FANCE wt Allele|Finding|true|false||face
null|FANCE gene|Finding|true|false||face
null|ELOVL6 gene|Finding|true|false||facenull|Head>Face|Anatomy|true|false||face
null|Face|Anatomy|true|false||facenull|Face (spatial concept)|Modifier|true|false||facenull|Fever|Finding|true|false||feversnull|Visual changes|Finding|false|false||visual changesnull|Visual|Finding|false|false||visualnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Eye symptom|Finding|false|false||eye symptomsnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Return to (contextual qualifier) (qualifier value)|Modifier|false|false||returnnull|Certification patient type - Urgent|Finding|false|false||urgent
null|Admission Type - Urgent|Finding|false|false||urgent
null|Triage Code - Urgent|Finding|false|false||urgent
null|Visit Priority Code - Urgent|Finding|false|false||urgentnull|Act Priority - urgent|Time|false|false||urgentnull|Urgent|Modifier|false|false||urgentnull|urgent - premium|LabModifier|false|false||urgentnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|true|false||changesnull|Pharmaceutical Preparations|Drug|true|false||medicationsnull|Medications|Finding|true|false||medicationsnull|null|Attribute|true|false||medications
null|null|Attribute|true|false||medicationsnull|follow-up|Procedure|true|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions