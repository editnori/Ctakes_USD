 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|44,53|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|44,53|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|44,58|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|78,87|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|78,87|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|78,92|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|134,137|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|145,152|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|145,152|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|154,162|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|165,174|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|165,174|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|165,174|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|186,195|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|186,195|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|186,195|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|198,220|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|206,210|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|206,210|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|206,220|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|211,220|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|223,232|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|223,232|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|246,255|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|257,266|false|false|false|||Epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|257,266|false|false|false|C0014591|Epistaxis|Epistaxis
Finding|Classification|SIMPLE_SEGMENT|269,274|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|287,305|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|296,305|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|296,305|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|296,305|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|296,305|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|296,305|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|315,322|true|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|315,322|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|315,322|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|315,322|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|315,325|true|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|315,341|true|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|315,341|true|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|326,333|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|326,333|true|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|326,341|true|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|334,341|true|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|366,373|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|366,376|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|377,380|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|377,380|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|SIMPLE_SEGMENT|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|SIMPLE_SEGMENT|377,380|false|false|false|||AAA
Finding|Gene or Genome|SIMPLE_SEGMENT|377,380|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|SIMPLE_SEGMENT|385,391|false|false|false|||repair
Finding|Functional Concept|SIMPLE_SEGMENT|385,391|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|385,391|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|385,391|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|385,391|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|SIMPLE_SEGMENT|393,404|false|false|false|||complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|412,424|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|412,424|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|430,444|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|430,444|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|430,444|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|449,457|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|464,472|false|false|false|||transfer
Finding|Functional Concept|SIMPLE_SEGMENT|464,472|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|464,472|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|464,472|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|SIMPLE_SEGMENT|486,494|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|486,494|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|500,505|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|500,505|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|500,505|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|506,515|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|506,515|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|506,515|false|false|false|C4554413|Fractured|fractures
Event|Event|SIMPLE_SEGMENT|521,530|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|521,530|false|false|false|C0014591|Epistaxis|epistaxis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|531,540|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|531,540|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|531,540|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|544,548|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|544,548|false|false|false|C0085639|Falls|fall
Finding|Body Substance|SIMPLE_SEGMENT|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|562,569|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|624,632|false|false|false|||coughing
Event|Event|SIMPLE_SEGMENT|637,644|false|false|false|||tripped
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|653,657|false|false|false|C0263940|Curb|curb
Event|Event|SIMPLE_SEGMENT|653,657|false|false|false|||curb
Event|Event|SIMPLE_SEGMENT|662,670|false|false|false|||suffered
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|671,677|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|671,677|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|671,677|false|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|685,689|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|685,689|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|685,689|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|685,689|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|701,705|true|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|701,705|true|false|false|C5890125|Loss (adaptation)|loss
Event|Event|SIMPLE_SEGMENT|710,723|true|false|false|||consciousness
Finding|Finding|SIMPLE_SEGMENT|710,723|true|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|SIMPLE_SEGMENT|710,723|true|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Event|Event|SIMPLE_SEGMENT|754,763|false|false|false|||nosebleed
Event|Event|SIMPLE_SEGMENT|769,777|false|false|false|||appeared
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|791,797|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|791,797|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|791,797|false|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|805,809|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|805,809|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|805,809|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|805,809|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|820,831|false|false|false|||transferred
Event|Activity|SIMPLE_SEGMENT|852,856|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|852,856|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|852,856|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|852,856|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|867,874|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|870,874|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|870,874|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Location or Region|SIMPLE_SEGMENT|883,887|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|883,887|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|883,887|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|883,887|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|883,887|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|889,893|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|889,893|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|889,893|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|899,903|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|899,903|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|SIMPLE_SEGMENT|899,903|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|909,919|false|false|false|||remarkable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|926,931|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|926,931|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|926,931|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|926,936|false|false|false|C0027422|Nasal bone structure|nasal bone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|932,936|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|932,936|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|932,936|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|949,957|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|949,957|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|976,985|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|976,985|false|false|false|C0014591|Epistaxis|epistaxis
Event|Event|SIMPLE_SEGMENT|998,1010|false|false|false|||RhinoRockets
Event|Event|SIMPLE_SEGMENT|1016,1022|false|false|false|||placed
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1039,1047|false|false|false|C0043242;C0518443;C1302752|Abrasion;Superficial abrasion;skin abrasion|abrasion
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1039,1047|false|false|false|C1627366|Abrasion Pharmacologic Substance|abrasion
Event|Event|SIMPLE_SEGMENT|1039,1047|false|false|false|||abrasion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1039,1047|false|false|false|C0580209|Surgical abrasion|abrasion
Event|Event|SIMPLE_SEGMENT|1055,1061|false|false|false|||bridge
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1055,1061|false|false|false|C0399080|Fixation of dental bridge|bridge
Event|Event|SIMPLE_SEGMENT|1089,1095|true|false|false|||closed
Event|Event|SIMPLE_SEGMENT|1097,1105|false|false|false|||Bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|1097,1105|false|false|false|C0019080|Hemorrhage|Bleeding
Finding|Finding|SIMPLE_SEGMENT|1110,1114|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|1115,1125|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|1159,1166|false|false|false|||episode
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1170,1176|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1170,1176|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1170,1176|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|1181,1188|false|false|false|||coughed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1198,1203|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|1198,1203|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|1198,1203|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|1222,1227|false|false|false|||began
Event|Event|SIMPLE_SEGMENT|1231,1235|false|false|false|||feel
Event|Event|SIMPLE_SEGMENT|1236,1247|false|false|false|||lightheaded
Finding|Sign or Symptom|SIMPLE_SEGMENT|1236,1247|false|false|false|C0220870|Lightheadedness|lightheaded
Event|Event|SIMPLE_SEGMENT|1257,1262|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|1269,1280|false|false|false|||hypotensive
Finding|Pathologic Function|SIMPLE_SEGMENT|1269,1280|false|false|false|C0857353|Hypotensive|hypotensive
Event|Event|SIMPLE_SEGMENT|1285,1296|false|false|false|||bradycardic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1302,1308|false|false|false|C4255046||report
Event|Event|SIMPLE_SEGMENT|1302,1308|false|false|false|||report
Finding|Intellectual Product|SIMPLE_SEGMENT|1302,1308|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|1302,1308|false|false|false|C0700287|Reporting|report
Finding|Intellectual Product|SIMPLE_SEGMENT|1320,1325|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1320,1347|false|false|false|C0234431|Brief loss of consciousness|brief loss of consciousness
Event|Event|SIMPLE_SEGMENT|1326,1330|false|false|false|||loss
Finding|Finding|SIMPLE_SEGMENT|1326,1330|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|SIMPLE_SEGMENT|1326,1347|false|false|false|C0041657|Unconscious State|loss of consciousness
Event|Event|SIMPLE_SEGMENT|1334,1347|false|false|false|||consciousness
Finding|Finding|SIMPLE_SEGMENT|1334,1347|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|SIMPLE_SEGMENT|1334,1347|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Event|Event|SIMPLE_SEGMENT|1364,1372|false|false|false|||returned
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1381,1389|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1381,1389|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1381,1389|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|SIMPLE_SEGMENT|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|SIMPLE_SEGMENT|1402,1407|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1417,1421|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1417,1421|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|1422,1428|false|false|false|||rolled
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1444,1448|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1444,1448|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1444,1448|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|1444,1448|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1444,1448|false|false|false|C0876917|Procedure on head|head
Finding|Body Substance|SIMPLE_SEGMENT|1454,1461|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1454,1461|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1454,1461|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1462,1469|true|false|false|||recalls
Event|Event|SIMPLE_SEGMENT|1474,1479|true|false|false|C0441471|Event|event
Event|Event|SIMPLE_SEGMENT|1484,1490|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1491,1501|true|false|false|||post-event
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1503,1512|true|false|false|C0009676|Confusion|confusion
Event|Event|SIMPLE_SEGMENT|1503,1512|true|false|false|||confusion
Finding|Finding|SIMPLE_SEGMENT|1503,1512|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|SIMPLE_SEGMENT|1532,1540|true|false|false|||episodes
Event|Event|SIMPLE_SEGMENT|1544,1551|true|false|false|||syncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|1544,1551|true|false|false|C0039070|Syncope|syncope
Event|Event|SIMPLE_SEGMENT|1555,1566|true|false|false|||hemodynamic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1555,1566|true|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1555,1566|true|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Event|Event|SIMPLE_SEGMENT|1568,1575|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1568,1575|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|1597,1602|false|false|false|C0441471|Event|event
Event|Event|SIMPLE_SEGMENT|1607,1616|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|1607,1616|false|false|false|C0014591|Epistaxis|epistaxis
Finding|Body Substance|SIMPLE_SEGMENT|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1635,1646|false|false|false|||transferred
Event|Activity|SIMPLE_SEGMENT|1659,1663|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|1659,1663|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|1659,1663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|1659,1663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|SIMPLE_SEGMENT|1677,1684|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|SIMPLE_SEGMENT|1685,1690|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1685,1696|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|1685,1696|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|SIMPLE_SEGMENT|1691,1696|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|1691,1696|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1691,1696|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1724,1728|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|SIMPLE_SEGMENT|1735,1742|false|false|false|||notable
Anatomy|Cell|SIMPLE_SEGMENT|1747,1750|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|1779,1782|false|false|false|||plt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1779,1782|false|false|false|C0201617|Primed lymphocyte test|plt
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1788,1791|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1788,1791|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|SIMPLE_SEGMENT|1788,1791|false|false|false|||BUN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1788,1791|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Event|Event|SIMPLE_SEGMENT|1804,1808|false|false|false|||HCTs
Event|Event|SIMPLE_SEGMENT|1814,1822|false|false|false|||repeated
Event|Event|SIMPLE_SEGMENT|1834,1840|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|1834,1840|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|1844,1854|false|false|false|||urinalysis
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1844,1854|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|urinalysis
Event|Event|SIMPLE_SEGMENT|1860,1868|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|1860,1868|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|1860,1868|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1860,1868|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|1872,1875|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1872,1875|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|1876,1888|false|false|false|||demonstrated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1897,1910|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|1897,1910|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|1918,1922|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1924,1928|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1924,1928|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1924,1928|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1924,1928|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1924,1933|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1929,1933|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Event|Event|SIMPLE_SEGMENT|1929,1933|false|false|false|||base
Finding|Gene or Genome|SIMPLE_SEGMENT|1929,1933|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|1929,1933|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Finding|SIMPLE_SEGMENT|1935,1943|false|false|false|C0332149|Possible|possibly
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1957,1967|false|false|false|C1720922|Respiratory Aspiration|aspiration
Event|Event|SIMPLE_SEGMENT|1957,1967|false|false|false|||aspiration
Finding|Finding|SIMPLE_SEGMENT|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1957,1967|false|false|false|C0349707||aspiration
Event|Event|SIMPLE_SEGMENT|1971,1981|false|false|false|||developing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1983,1992|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|SIMPLE_SEGMENT|1983,1992|false|false|false|||pneumonia
Finding|Body Substance|SIMPLE_SEGMENT|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Immunologic Factor|SIMPLE_SEGMENT|2016,2020|false|false|false|C3526553;C3644171|diphtheria, tetanus toxoids and acellular pertussis vaccine;tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Tdap
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2016,2020|false|false|false|C3526553;C3644171|diphtheria, tetanus toxoids and acellular pertussis vaccine;tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Tdap
Drug|Antibiotic|SIMPLE_SEGMENT|2022,2033|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|2022,2033|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|SIMPLE_SEGMENT|2022,2033|false|false|false|||amoxicillin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2022,2045|false|false|false|C0054066|amoxicillin / clavulanate|amoxicillin-clavulanate
Drug|Antibiotic|SIMPLE_SEGMENT|2034,2045|false|false|false|C0110038|clavulanate|clavulanate
Drug|Organic Chemical|SIMPLE_SEGMENT|2034,2045|false|false|false|C0110038|clavulanate|clavulanate
Event|Event|SIMPLE_SEGMENT|2034,2045|false|false|false|||clavulanate
Drug|Antibiotic|SIMPLE_SEGMENT|2051,2061|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2051,2073|false|false|false|C0282638|Antibiotic Prophylaxis|antibiotic prophylaxis
Event|Event|SIMPLE_SEGMENT|2062,2073|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2062,2073|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Organic Chemical|SIMPLE_SEGMENT|2075,2086|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2075,2086|false|false|false|C0061851|ondansetron|ondansetron
Event|Event|SIMPLE_SEGMENT|2075,2086|false|false|false|||ondansetron
Drug|Organic Chemical|SIMPLE_SEGMENT|2103,2113|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2103,2113|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|2103,2113|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|2103,2122|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2103,2122|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|2114,2122|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2114,2122|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|2123,2127|false|false|false|||50mg
Drug|Organic Chemical|SIMPLE_SEGMENT|2129,2140|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2129,2140|false|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|SIMPLE_SEGMENT|2129,2140|false|false|false|||Clopidogrel
Event|Event|SIMPLE_SEGMENT|2145,2149|false|false|false|||held
Finding|Finding|SIMPLE_SEGMENT|2153,2173|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2158,2165|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2158,2165|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2158,2165|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2158,2165|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2158,2165|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2158,2173|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2166,2173|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2166,2173|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2166,2173|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2184,2187|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2184,2187|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|SIMPLE_SEGMENT|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|SIMPLE_SEGMENT|2184,2187|false|false|false|||AAA
Finding|Gene or Genome|SIMPLE_SEGMENT|2184,2187|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|SIMPLE_SEGMENT|2188,2194|false|false|false|||repair
Finding|Functional Concept|SIMPLE_SEGMENT|2188,2194|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|2188,2194|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|2188,2194|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2188,2194|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2215,2218|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|2215,2218|false|false|false|||HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2219,2239|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|SIMPLE_SEGMENT|2219,2239|false|false|false|||Hypercholesterolemia
Finding|Finding|SIMPLE_SEGMENT|2219,2239|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Finding|Functional Concept|SIMPLE_SEGMENT|2242,2248|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2242,2256|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2249,2256|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2249,2256|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2249,2256|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2249,2256|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2262,2268|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2262,2268|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2262,2268|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2262,2268|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2262,2276|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2269,2276|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2269,2276|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2269,2276|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2269,2276|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Body Substance|SIMPLE_SEGMENT|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|2289,2296|false|false|false|||unaware
Procedure|Research Activity|SIMPLE_SEGMENT|2289,2296|false|false|false|C0150114|unaware|unaware
Finding|Classification|SIMPLE_SEGMENT|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|2302,2316|false|false|false|C0241889|Family Medical History|family history
Finding|Finding|SIMPLE_SEGMENT|2302,2319|false|false|false|C0241889|Family Medical History|family history of
Event|Event|SIMPLE_SEGMENT|2309,2316|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2309,2319|false|false|false|C0262926|Medical History|history of
Finding|Pathologic Function|SIMPLE_SEGMENT|2320,2328|false|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2320,2338|false|false|false|C0005779|Blood Coagulation Disorders|bleeding diathesis
Finding|Pathologic Function|SIMPLE_SEGMENT|2320,2338|false|false|false|C1458140|Bleeding tendency|bleeding diathesis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2329,2338|false|false|false|C0012655|Disease susceptibility|diathesis
Event|Event|SIMPLE_SEGMENT|2329,2338|false|false|false|||diathesis
Event|Event|SIMPLE_SEGMENT|2343,2351|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2343,2351|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2343,2351|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2343,2351|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2343,2356|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2343,2356|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2352,2356|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2352,2356|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2352,2356|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2358,2367|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2396,2403|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2396,2403|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2396,2403|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2405,2410|true|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2405,2410|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2405,2410|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2405,2410|true|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2405,2410|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2405,2410|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2405,2410|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|2412,2420|true|false|false|||oriented
Finding|Intellectual Product|SIMPLE_SEGMENT|2425,2430|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|2431,2439|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2431,2439|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2431,2439|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2442,2447|true|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2457,2466|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2457,2466|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2468,2471|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2468,2471|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2473,2483|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|2484,2489|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2484,2489|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2491,2499|false|false|false|C0009938|Contusions|bruising
Event|Event|SIMPLE_SEGMENT|2491,2499|false|false|false|||bruising
Finding|Finding|SIMPLE_SEGMENT|2491,2499|false|false|false|C2136686|reported bruising (history)|bruising
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2507,2516|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2512,2516|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2512,2516|false|false|false|C5848506||eyes
Finding|Finding|SIMPLE_SEGMENT|2518,2525|false|false|false|C0038999|Swelling|swollen
Finding|Finding|SIMPLE_SEGMENT|2518,2530|false|false|false|C0240577|Swollen nose|swollen nose
Event|Event|SIMPLE_SEGMENT|2526,2530|false|false|false|||nose
Finding|Intellectual Product|SIMPLE_SEGMENT|2536,2540|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|2541,2551|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2541,2551|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2541,2551|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Activity|SIMPLE_SEGMENT|2570,2575|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|2570,2575|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|2570,2575|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|2570,2575|false|false|false|C1533810||place
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2578,2582|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2578,2582|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2578,2582|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|2584,2590|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|2584,2590|true|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2600,2603|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2600,2603|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|2600,2603|true|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2600,2603|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2606,2610|true|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2606,2610|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Event|Event|SIMPLE_SEGMENT|2606,2610|true|false|false|||RESP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2622,2625|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|2622,2625|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2622,2625|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2622,2625|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|SIMPLE_SEGMENT|2644,2647|false|false|false|||RRR
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2669,2672|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2669,2672|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|2669,2672|true|false|false|||ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2674,2678|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|2674,2678|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|2710,2718|false|false|false|||Deferred
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2720,2723|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|SIMPLE_SEGMENT|2720,2723|false|false|false|||EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|2720,2723|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|SIMPLE_SEGMENT|2725,2729|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|2725,2729|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2725,2729|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|2731,2735|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2736,2744|true|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|2749,2755|true|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2749,2755|true|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2749,2755|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2749,2755|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2760,2768|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|2760,2768|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|2770,2778|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|2770,2778|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2783,2788|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2783,2788|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2783,2788|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|2816,2822|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2816,2822|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|SIMPLE_SEGMENT|2824,2829|false|false|false|C1513492|motor movement|motor
Finding|Finding|SIMPLE_SEGMENT|2824,2838|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2824,2838|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|SIMPLE_SEGMENT|2830,2838|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|2847,2853|false|false|false|||normal
Anatomy|Body System|SIMPLE_SEGMENT|2854,2858|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2854,2858|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2854,2858|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|2854,2858|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|2854,2858|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|2854,2858|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2863,2875|true|false|false|C0015256|Excoriation|excoriations
Event|Event|SIMPLE_SEGMENT|2863,2875|true|false|false|||excoriations
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2879,2883|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|2879,2883|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|2879,2883|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|2879,2883|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|2886,2895|false|false|false|||DISCHARGE
Finding|Body Substance|SIMPLE_SEGMENT|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2886,2895|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2924,2931|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2924,2931|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2924,2931|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2933,2938|true|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2933,2938|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2933,2938|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2933,2938|true|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2933,2938|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2933,2938|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2933,2938|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|2940,2948|true|false|false|||oriented
Finding|Intellectual Product|SIMPLE_SEGMENT|2953,2958|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|2959,2967|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2959,2967|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2959,2967|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2970,2975|true|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2985,2994|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2985,2994|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2996,2999|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2996,2999|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3001,3011|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|3012,3017|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3012,3017|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3019,3027|false|false|false|C0009938|Contusions|bruising
Event|Event|SIMPLE_SEGMENT|3019,3027|false|false|false|||bruising
Finding|Finding|SIMPLE_SEGMENT|3019,3027|false|false|false|C2136686|reported bruising (history)|bruising
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3035,3044|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3040,3044|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3040,3044|false|false|false|C5848506||eyes
Finding|Finding|SIMPLE_SEGMENT|3046,3053|false|false|false|C0038999|Swelling|swollen
Finding|Finding|SIMPLE_SEGMENT|3046,3058|false|false|false|C0240577|Swollen nose|swollen nose
Event|Event|SIMPLE_SEGMENT|3054,3058|false|false|false|||nose
Finding|Intellectual Product|SIMPLE_SEGMENT|3064,3068|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|3069,3079|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3069,3079|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3069,3079|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Activity|SIMPLE_SEGMENT|3098,3103|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3098,3103|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3098,3103|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3098,3103|false|false|false|C1533810||place
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3106,3110|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3106,3110|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3106,3110|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|SIMPLE_SEGMENT|3112,3118|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|3112,3118|true|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3128,3131|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3128,3131|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|3128,3131|true|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3128,3131|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3134,3138|true|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3134,3138|true|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Event|Event|SIMPLE_SEGMENT|3134,3138|true|false|false|||RESP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3150,3153|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|SIMPLE_SEGMENT|3150,3153|false|false|false|||CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|3150,3153|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3150,3153|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|SIMPLE_SEGMENT|3172,3175|false|false|false|||RRR
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3197,3200|true|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|3197,3200|true|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|3197,3200|true|false|false|||ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3202,3206|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|SIMPLE_SEGMENT|3202,3206|false|false|false|||Soft
Event|Event|SIMPLE_SEGMENT|3238,3246|false|false|false|||Deferred
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3248,3251|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|SIMPLE_SEGMENT|3248,3251|false|false|false|||EXT
Finding|Gene or Genome|SIMPLE_SEGMENT|3248,3251|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|SIMPLE_SEGMENT|3253,3257|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|3253,3257|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3253,3257|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3259,3263|true|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3264,3272|true|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3277,3283|true|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3277,3283|true|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3277,3283|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3277,3283|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|3288,3296|true|false|false|C0149651|Clubbing|clubbing
Event|Event|SIMPLE_SEGMENT|3288,3296|true|false|false|||clubbing
Event|Event|SIMPLE_SEGMENT|3298,3306|true|false|false|||cyanosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3298,3306|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3311,3316|true|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|3311,3316|true|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|3311,3316|true|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3344,3350|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3344,3350|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|SIMPLE_SEGMENT|3352,3357|false|false|false|C1513492|motor movement|motor
Finding|Finding|SIMPLE_SEGMENT|3352,3366|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3352,3366|false|false|false|C0234130|Motor function (observable entity)|motor function
Event|Event|SIMPLE_SEGMENT|3358,3366|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|3375,3381|false|false|false|||normal
Anatomy|Body System|SIMPLE_SEGMENT|3382,3386|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3382,3386|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3382,3386|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3382,3386|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3382,3386|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3382,3386|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3391,3403|true|false|false|C0015256|Excoriation|excoriations
Event|Event|SIMPLE_SEGMENT|3391,3403|true|false|false|||excoriations
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3407,3411|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|3407,3411|true|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|3407,3411|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|3407,3411|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Procedure|Health Care Activity|SIMPLE_SEGMENT|3434,3443|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3457,3462|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3457,3462|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3457,3462|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3463,3466|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3473,3476|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3473,3476|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3473,3476|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3483,3486|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3483,3486|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3483,3486|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3483,3486|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3492,3495|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3492,3495|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3502,3505|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3502,3505|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3502,3505|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3502,3505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3502,3505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3509,3512|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3509,3512|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3509,3512|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3509,3512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3509,3512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3509,3512|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3519,3523|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3539,3542|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3559,3564|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3559,3564|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3559,3564|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3577,3583|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3599,3602|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3599,3602|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3599,3602|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3629,3634|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3629,3634|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3629,3634|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3639,3642|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3639,3642|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3639,3642|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3664,3669|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3664,3669|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3664,3669|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3664,3677|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3664,3677|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3664,3677|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3670,3677|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3670,3677|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3670,3677|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|3670,3677|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3670,3677|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3670,3677|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3725,3729|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3725,3729|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3725,3729|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3755,3760|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3755,3760|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3755,3760|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3764,3767|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|3764,3767|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|3764,3767|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|3764,3767|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3764,3767|false|false|false|C0201973|Creatine kinase measurement|CPK
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3775,3782|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3775,3782|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3775,3789|false|false|false|C1271630|Cardiac markers|CARDIAC MARKER
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3790,3795|false|false|false|C4554533||TREND
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3809,3814|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3809,3814|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3809,3814|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3841,3846|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3841,3846|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3841,3846|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3847,3852|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3847,3852|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3847,3852|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3847,3852|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3896,3901|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3896,3901|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3896,3901|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3902,3907|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3902,3907|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3902,3907|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3902,3907|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3950,3955|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3950,3955|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3950,3955|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3956,3961|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3956,3961|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3956,3961|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3956,3961|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3990,3995|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3990,3995|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3990,3995|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3996,4001|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|3996,4001|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|3996,4001|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3996,4001|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|3999,4003|false|false|false|C0602256|MB 5|MB-5
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4030,4035|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4030,4035|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4030,4035|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4036,4041|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4036,4041|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4036,4041|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4036,4041|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4070,4075|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4070,4075|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4070,4075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4076,4081|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|4076,4081|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|4076,4081|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4076,4081|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|SIMPLE_SEGMENT|4079,4083|false|false|false|C0602249|MB 2|MB-2
Finding|Body Substance|SIMPLE_SEGMENT|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|4099,4108|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|4109,4113|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4109,4113|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4127,4132|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4127,4132|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4127,4132|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4133,4136|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4141,4144|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4151,4154|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4151,4154|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4151,4154|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4151,4154|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4161,4164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4161,4164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4172,4175|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4172,4175|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4172,4175|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4172,4175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4172,4175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4179,4182|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4179,4182|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4179,4182|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4179,4182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4179,4182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4179,4182|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4189,4193|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4208,4211|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4228,4233|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4228,4233|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4228,4233|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4228,4241|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4228,4241|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4228,4241|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4234,4241|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4234,4241|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4234,4241|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4234,4241|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4234,4241|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4234,4241|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4289,4293|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4289,4293|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4289,4293|false|false|false|C0202059|Bicarbonate measurement|HCO3
Event|Event|SIMPLE_SEGMENT|4307,4314|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4307,4314|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4307,4314|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|4320,4323|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4320,4323|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|4339,4344|false|false|false|||views
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4352,4357|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|4352,4357|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|4358,4366|false|false|false|||provided
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4372,4377|false|false|false|C0024109|Lung|lungs
Event|Event|SIMPLE_SEGMENT|4395,4402|false|false|false|||aerated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4421,4434|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|4421,4434|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|4442,4446|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4442,4451|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4442,4456|false|false|false|C0225732|Structure of base of left lung|left lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4447,4451|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4447,4451|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4447,4451|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|4447,4451|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4447,4456|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4452,4456|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|SIMPLE_SEGMENT|4452,4456|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|SIMPLE_SEGMENT|4452,4456|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Event|Event|SIMPLE_SEGMENT|4458,4466|false|false|false|||adjacent
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4482,4495|false|false|false|C1269845|Structure of hemidiaphragm|hemidiaphragm
Finding|Intellectual Product|SIMPLE_SEGMENT|4506,4510|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4511,4519|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4521,4532|false|false|false|C0020452|Hyperemia|engorgement
Event|Event|SIMPLE_SEGMENT|4521,4532|false|false|false|||engorgement
Finding|Finding|SIMPLE_SEGMENT|4521,4532|false|false|false|C1706102|Tick Engorgement|engorgement
Finding|Finding|SIMPLE_SEGMENT|4553,4578|false|false|false|C5139173|Apical pulmonary opacity|apical pleural thickening
Anatomy|Tissue|SIMPLE_SEGMENT|4560,4567|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4560,4567|false|false|false|C0032226|Pleural Diseases|pleural
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4560,4578|false|false|false|C0264545|Thickening of pleura|pleural thickening
Event|Event|SIMPLE_SEGMENT|4568,4578|false|false|false|||thickening
Finding|Finding|SIMPLE_SEGMENT|4568,4578|false|false|false|C0205400|Thickened|thickening
Event|Event|SIMPLE_SEGMENT|4603,4613|false|false|false|||silhouette
Event|Event|SIMPLE_SEGMENT|4617,4627|false|false|false|||remarkable
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4632,4638|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4632,4643|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4632,4643|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|SIMPLE_SEGMENT|4639,4643|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|SIMPLE_SEGMENT|4639,4643|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Event|Event|SIMPLE_SEGMENT|4645,4659|false|false|false|||calcifications
Finding|Finding|SIMPLE_SEGMENT|4645,4659|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4645,4659|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4665,4670|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4665,4670|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|4665,4670|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|4665,4670|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|4678,4684|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|4700,4704|false|false|false|||ECHO
Procedure|Health Care Activity|SIMPLE_SEGMENT|4700,4704|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4700,4704|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|SIMPLE_SEGMENT|4709,4713|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4709,4720|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4714,4720|false|false|false|C0018792|Heart Atrium|atrium
Event|Event|SIMPLE_SEGMENT|4731,4738|false|false|false|||dilated
Finding|Functional Concept|SIMPLE_SEGMENT|4740,4744|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4740,4761|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4745,4756|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4745,4761|false|false|false|C0507618|Wall of ventricle|ventricular wall
Event|Event|SIMPLE_SEGMENT|4763,4774|false|false|false|||thicknesses
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4779,4785|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4779,4785|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4779,4785|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|4786,4790|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|4795,4801|false|false|false|||normal
Finding|Intellectual Product|SIMPLE_SEGMENT|4812,4816|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|4827,4831|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4827,4864|false|false|false|C1277187|Left ventricular systolic dysfunction|left ventricular systolic dysfunction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4832,4843|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4844,4852|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|SIMPLE_SEGMENT|4844,4864|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4853,4864|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|4853,4864|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Event|Event|SIMPLE_SEGMENT|4884,4895|false|false|false|||hypokinesis
Finding|Finding|SIMPLE_SEGMENT|4884,4895|false|false|false|C0086439|Hypokinesia|hypokinesis
Event|Event|SIMPLE_SEGMENT|4911,4919|false|false|false|||segments
Event|Event|SIMPLE_SEGMENT|4920,4928|false|false|false|||contract
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4939,4943|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Event|Event|SIMPLE_SEGMENT|4939,4943|false|false|false|||LVEF
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4939,4943|false|false|false|C3837267|LVEF (procedure)|LVEF
Event|Event|SIMPLE_SEGMENT|4957,4963|true|false|false|||masses
Event|Event|SIMPLE_SEGMENT|4967,4974|true|false|false|||thrombi
Finding|Pathologic Function|SIMPLE_SEGMENT|4967,4974|true|false|false|C0087086|Thrombus|thrombi
Event|Event|SIMPLE_SEGMENT|4979,4983|true|false|false|||seen
Finding|Functional Concept|SIMPLE_SEGMENT|4991,4995|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4991,5005|false|false|false|C0225897;C4266612|Chest>Heart.ventricle.left;Left ventricular structure|left ventricle
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4996,5005|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4996,5005|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Finding|Functional Concept|SIMPLE_SEGMENT|5007,5012|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5014,5025|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5026,5033|false|false|false|C0935616|chamber [body part]|chamber
Event|Event|SIMPLE_SEGMENT|5034,5038|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|5043,5047|false|false|false|||free
Finding|Functional Concept|SIMPLE_SEGMENT|5043,5047|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5048,5059|false|false|false|C1980023|Wall motion|wall motion
Event|Event|SIMPLE_SEGMENT|5053,5059|false|false|false|||motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5053,5059|false|false|false|C0026597|Motion|motion
Event|Event|SIMPLE_SEGMENT|5064,5070|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5089,5095|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5089,5101|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5096,5101|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5102,5110|false|false|false|||leaflets
Finding|Intellectual Product|SIMPLE_SEGMENT|5121,5125|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5126,5132|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5126,5138|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5133,5138|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5140,5148|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5140,5148|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5150,5155|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|SIMPLE_SEGMENT|5150,5160|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|SIMPLE_SEGMENT|5156,5160|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5164,5167|false|false|false|C0555206|Chiari malformation type II|cm2
Finding|Intellectual Product|SIMPLE_SEGMENT|5170,5174|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5180,5186|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5180,5200|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Event|Event|SIMPLE_SEGMENT|5187,5200|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5187,5200|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5187,5200|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5187,5200|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|5205,5209|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5215,5227|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5222,5227|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5228,5236|false|false|false|||leaflets
Event|Event|SIMPLE_SEGMENT|5248,5257|false|false|false|||thickened
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5268,5288|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Event|Event|SIMPLE_SEGMENT|5275,5288|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5275,5288|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5275,5288|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5275,5288|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Event|Event|SIMPLE_SEGMENT|5292,5296|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5302,5311|true|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5302,5311|true|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|5302,5311|true|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5302,5318|true|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5312,5318|true|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|5312,5318|true|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|5319,5327|true|false|false|||systolic
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5319,5327|true|false|false|C0039155|Systole|systolic
Event|Event|SIMPLE_SEGMENT|5329,5337|true|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|5329,5337|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|5329,5337|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5329,5337|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5329,5337|true|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|5351,5361|true|false|false|||determined
Finding|Functional Concept|SIMPLE_SEGMENT|5382,5393|false|false|false|C0205463|Physiological|physiologic
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5395,5406|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5395,5406|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5395,5415|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|SIMPLE_SEGMENT|5395,5415|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|SIMPLE_SEGMENT|5407,5415|false|false|false|||effusion
Finding|Body Substance|SIMPLE_SEGMENT|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|SIMPLE_SEGMENT|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|SIMPLE_SEGMENT|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Event|Event|SIMPLE_SEGMENT|5419,5429|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5419,5429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5419,5429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Functional Concept|SIMPLE_SEGMENT|5438,5442|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5438,5461|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5438,5466|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5443,5454|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5443,5461|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5455,5461|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5455,5461|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5455,5461|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Event|Event|SIMPLE_SEGMENT|5462,5466|false|false|false|||size
Event|Event|SIMPLE_SEGMENT|5472,5476|false|false|false|||mild
Finding|Intellectual Product|SIMPLE_SEGMENT|5472,5476|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5487,5495|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|SIMPLE_SEGMENT|5487,5507|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5496,5507|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Event|Event|SIMPLE_SEGMENT|5496,5507|false|false|false|||dysfunction
Finding|Conceptual Entity|SIMPLE_SEGMENT|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|SIMPLE_SEGMENT|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|SIMPLE_SEGMENT|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5517,5520|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5517,5520|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|5517,5520|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|5517,5520|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5517,5520|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5522,5528|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5529,5532|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5529,5532|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|SIMPLE_SEGMENT|5529,5532|false|false|false|||LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5529,5532|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|SIMPLE_SEGMENT|5534,5546|false|false|false|||distribution
Finding|Cell Function|SIMPLE_SEGMENT|5534,5546|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|SIMPLE_SEGMENT|5534,5546|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Intellectual Product|SIMPLE_SEGMENT|5549,5553|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5549,5575|false|false|false|C3276923|Mild aortic valve stenosis|Mild aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5554,5560|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5554,5566|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5554,5575|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5554,5575|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5554,5575|false|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5561,5566|false|false|false|C1186983|Anatomical valve|valve
Event|Event|SIMPLE_SEGMENT|5567,5575|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5567,5575|false|false|false|C1261287|Stenosis|stenosis
Finding|Intellectual Product|SIMPLE_SEGMENT|5577,5581|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5582,5588|false|false|false|C0003483|Aorta|aortic
Event|Event|SIMPLE_SEGMENT|5590,5603|false|false|false|||regurgitation
Finding|Finding|SIMPLE_SEGMENT|5590,5603|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5590,5603|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5590,5603|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Intellectual Product|SIMPLE_SEGMENT|5608,5613|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5614,5622|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5614,5629|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5614,5629|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|5654,5661|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5654,5664|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5665,5668|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5665,5668|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|SIMPLE_SEGMENT|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|SIMPLE_SEGMENT|5665,5668|false|false|false|||AAA
Finding|Gene or Genome|SIMPLE_SEGMENT|5665,5668|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|SIMPLE_SEGMENT|5673,5679|false|false|false|||repair
Finding|Functional Concept|SIMPLE_SEGMENT|5673,5679|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|5673,5679|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|5673,5679|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5673,5679|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|SIMPLE_SEGMENT|5681,5692|false|false|false|||complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5700,5712|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|5700,5712|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5718,5732|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|5718,5732|false|false|false|||hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|5718,5732|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|SIMPLE_SEGMENT|5738,5747|false|false|false|||presented
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5753,5758|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|5753,5758|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|5753,5758|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5759,5768|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|5759,5768|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|5759,5768|false|false|false|C4554413|Fractured|fractures
Event|Event|SIMPLE_SEGMENT|5773,5782|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|5773,5782|false|false|false|C0014591|Epistaxis|epistaxis
Event|Event|SIMPLE_SEGMENT|5789,5799|false|false|false|||mechanical
Finding|Functional Concept|SIMPLE_SEGMENT|5789,5799|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5789,5799|false|false|false|C0699886|Mechanical Treatments|mechanical
Event|Event|SIMPLE_SEGMENT|5801,5805|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|5801,5805|false|false|false|C0085639|Falls|fall
Finding|Idea or Concept|SIMPLE_SEGMENT|5811,5819|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5811,5826|false|false|false|C0488549||hospital course
Finding|Finding|SIMPLE_SEGMENT|5811,5826|false|false|false|C0489547|Hospital course|hospital course
Event|Event|SIMPLE_SEGMENT|5820,5826|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|5827,5838|false|false|false|||complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5842,5848|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|5842,5848|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|5842,5848|false|false|false|C3537184||NSTEMI
Event|Event|SIMPLE_SEGMENT|5852,5861|false|false|false|||Epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|5852,5861|false|false|false|C0014591|Epistaxis|Epistaxis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5863,5868|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|5863,5868|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|5863,5868|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5869,5878|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|5869,5878|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|5869,5878|false|false|false|C4554413|Fractured|fractures
Finding|Body Substance|SIMPLE_SEGMENT|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|5887,5897|false|false|false|||presenting
Event|Event|SIMPLE_SEGMENT|5904,5914|false|false|false|||mechanical
Finding|Functional Concept|SIMPLE_SEGMENT|5904,5914|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5904,5914|false|false|false|C0699886|Mechanical Treatments|mechanical
Event|Event|SIMPLE_SEGMENT|5915,5919|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|5915,5919|false|false|false|C0085639|Falls|fall
Event|Event|SIMPLE_SEGMENT|5925,5937|false|false|false|||Rhinorockets
Event|Event|SIMPLE_SEGMENT|5939,5945|false|false|false|||placed
Finding|Idea or Concept|SIMPLE_SEGMENT|5957,5965|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|5970,5977|false|false|false|C0549178|Continuous|ongoing
Event|Event|SIMPLE_SEGMENT|5978,5987|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|5978,5987|false|false|false|C0014591|Epistaxis|epistaxis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5989,5996|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Event|Event|SIMPLE_SEGMENT|5992,5996|false|false|false|||scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5992,5996|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Event|SIMPLE_SEGMENT|6008,6016|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|6008,6016|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|6017,6029|false|false|false|||demonstrated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6030,6035|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|6030,6035|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|6030,6035|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6030,6040|false|false|false|C0027422|Nasal bone structure|nasal bone
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6036,6040|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|6036,6040|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|6036,6040|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|6052,6061|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|6052,6061|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|6052,6061|false|false|false|C4554413|Fractured|fractures
Event|Event|SIMPLE_SEGMENT|6086,6096|false|false|false|||maintained
Event|Event|SIMPLE_SEGMENT|6103,6112|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|6103,6112|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|6103,6112|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|6117,6129|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|6140,6149|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6140,6149|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|6158,6168|false|false|false|||encouraged
Event|Event|SIMPLE_SEGMENT|6172,6175|false|false|false|||use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6190,6195|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|6190,6195|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|6190,6195|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6197,6202|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|SIMPLE_SEGMENT|6197,6202|false|false|false|C2003858|Spray (action)|spray
Event|Event|SIMPLE_SEGMENT|6197,6202|false|false|false|||spray
Finding|Functional Concept|SIMPLE_SEGMENT|6197,6202|false|false|false|C4521772|Spray (administration method)|spray
Event|Activity|SIMPLE_SEGMENT|6207,6211|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|SIMPLE_SEGMENT|6207,6211|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|SIMPLE_SEGMENT|6207,6211|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Event|Event|SIMPLE_SEGMENT|6212,6220|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6212,6220|false|false|false|C0033095||pressure
Event|Event|SIMPLE_SEGMENT|6228,6236|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|6228,6236|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|6237,6244|false|false|false|||reoccur
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6249,6255|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|6249,6255|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|6249,6255|false|false|false|C3537184||NSTEMI
Finding|Body Substance|SIMPLE_SEGMENT|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6264,6269|false|false|false|||found
Finding|Intellectual Product|SIMPLE_SEGMENT|6278,6282|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|6283,6292|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6283,6292|false|false|false|C0439775|Elevation procedure|elevation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6296,6304|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6296,6304|false|false|false|C0041199|Troponin|troponin
Event|Event|SIMPLE_SEGMENT|6296,6304|false|false|false|||troponin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6296,6304|false|false|false|C0523952|Troponin measurement|troponin
Event|Event|SIMPLE_SEGMENT|6326,6333|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|6349,6353|false|false|false|||rose
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6372,6381|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6372,6381|false|false|false|C1179435|Protein Component|component
Event|Event|SIMPLE_SEGMENT|6372,6381|false|false|false|||component
Finding|Conceptual Entity|SIMPLE_SEGMENT|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|SIMPLE_SEGMENT|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|SIMPLE_SEGMENT|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|SIMPLE_SEGMENT|6383,6394|false|false|false|||downtrended
Event|Event|SIMPLE_SEGMENT|6402,6408|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|6412,6421|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6412,6421|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|SIMPLE_SEGMENT|6427,6434|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6427,6434|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6427,6434|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6448,6453|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|6448,6453|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6448,6458|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6448,6458|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6454,6458|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6454,6458|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6454,6458|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6454,6458|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6468,6475|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|6468,6475|true|false|false|C1314974|Cardiac attachment|cardiac
Finding|Sign or Symptom|SIMPLE_SEGMENT|6468,6484|true|false|false|C0741933|cardiac symptom|cardiac symptoms
Event|Event|SIMPLE_SEGMENT|6476,6484|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|6476,6484|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|6476,6484|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body System|SIMPLE_SEGMENT|6486,6496|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Event|SIMPLE_SEGMENT|6501,6510|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|6516,6523|false|false|false|||thought
Finding|Idea or Concept|SIMPLE_SEGMENT|6538,6549|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|6543,6549|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6543,6549|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6550,6559|false|true|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|6550,6559|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6550,6559|false|true|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|6563,6569|false|false|false|||demand
Finding|Idea or Concept|SIMPLE_SEGMENT|6563,6569|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6563,6569|false|false|false|C0441516|Demand (clinical)|demand
Event|Event|SIMPLE_SEGMENT|6571,6579|false|false|false|||ischemia
Finding|Pathologic Function|SIMPLE_SEGMENT|6571,6579|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6571,6579|false|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Gene or Genome|SIMPLE_SEGMENT|6581,6585|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|6581,6585|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6593,6602|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|SIMPLE_SEGMENT|6593,6602|false|false|false|||secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6593,6602|false|false|false|C1522484|metastatic qualifier|secondary
Event|Event|SIMPLE_SEGMENT|6610,6614|false|false|false|||fall
Finding|Finding|SIMPLE_SEGMENT|6610,6614|false|false|false|C0085639|Falls|fall
Event|Event|SIMPLE_SEGMENT|6619,6633|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6619,6633|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|6635,6647|false|false|false|||demonstrated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6648,6654|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|SIMPLE_SEGMENT|6648,6663|false|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Event|Event|SIMPLE_SEGMENT|6655,6663|false|false|false|||stenosis
Finding|Pathologic Function|SIMPLE_SEGMENT|6655,6663|false|false|false|C1261287|Stenosis|stenosis
Finding|Finding|SIMPLE_SEGMENT|6668,6674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6668,6674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6675,6681|false|true|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6682,6685|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6682,6685|false|true|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|6682,6685|false|true|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6686,6693|false|true|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|6686,6693|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6704,6715|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6709,6715|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|6716,6729|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|6716,6729|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|6716,6729|false|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|SIMPLE_SEGMENT|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|6745,6755|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6745,6755|false|false|false|C0025859|metoprolol|metoprolol
Event|Event|SIMPLE_SEGMENT|6745,6755|false|false|false|||metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|6777,6788|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6777,6788|false|false|false|C0085542|pravastatin|pravastatin
Event|Event|SIMPLE_SEGMENT|6777,6788|false|false|false|||pravastatin
Event|Event|SIMPLE_SEGMENT|6793,6802|false|false|false|||converted
Drug|Organic Chemical|SIMPLE_SEGMENT|6806,6818|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6806,6818|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|6806,6818|false|false|false|||atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|6825,6836|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6825,6836|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|SIMPLE_SEGMENT|6825,6836|false|false|false|||clopidogrel
Event|Event|SIMPLE_SEGMENT|6841,6851|false|false|false|||maintained
Event|Event|SIMPLE_SEGMENT|6864,6871|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|6875,6882|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6875,6882|false|false|false|C0004057|aspirin|aspirin
Event|Event|SIMPLE_SEGMENT|6875,6882|false|false|false|||aspirin
Event|Event|SIMPLE_SEGMENT|6886,6895|false|false|false|||Hypoxemia
Finding|Finding|SIMPLE_SEGMENT|6886,6895|false|false|false|C0700292;C5548348|Blood oxygen concentration below reference range (finding);Hypoxemia|Hypoxemia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6906,6919|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|6906,6919|false|false|false|||consolidation
Finding|Body Substance|SIMPLE_SEGMENT|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|6928,6936|false|false|false|||reported
Event|Event|SIMPLE_SEGMENT|6950,6957|false|false|false|||hypoxic
Finding|Pathologic Function|SIMPLE_SEGMENT|6950,6957|false|false|false|C0242184|Hypoxia|hypoxic
Event|Event|SIMPLE_SEGMENT|6980,6990|false|false|false|||maintained
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6998,7004|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6998,7004|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6998,7004|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6998,7004|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6998,7016|false|false|false|C0483415|Oxygen Saturation|oxygen saturations
Event|Event|SIMPLE_SEGMENT|7005,7016|false|false|false|||saturations
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7005,7016|false|false|false|C0522534|Saturated|saturations
Finding|Finding|SIMPLE_SEGMENT|7017,7028|false|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7020,7028|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Event|Event|SIMPLE_SEGMENT|7025,7028|false|false|false|||air
Finding|Finding|SIMPLE_SEGMENT|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|SIMPLE_SEGMENT|7033,7039|false|false|false|||denied
Event|Event|SIMPLE_SEGMENT|7041,7050|true|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7041,7060|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|7041,7060|true|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|SIMPLE_SEGMENT|7054,7060|true|false|false|||breath
Finding|Body Substance|SIMPLE_SEGMENT|7054,7060|true|false|false|C0225386|Breath|breath
Drug|Organic Chemical|SIMPLE_SEGMENT|7064,7069|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7064,7069|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|7064,7069|true|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|7064,7069|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|7071,7077|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|7071,7077|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7088,7098|true|false|false|C0009450|Communicable Diseases|infectious
Event|Event|SIMPLE_SEGMENT|7088,7098|true|false|false|||infectious
Event|Event|SIMPLE_SEGMENT|7100,7108|true|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|7100,7108|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|7100,7108|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7120,7132|true|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|7120,7132|true|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|7120,7132|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|7136,7139|false|false|false|||CXR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7136,7139|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|SIMPLE_SEGMENT|7140,7148|false|false|false|||revealed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7149,7162|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|SIMPLE_SEGMENT|7149,7162|false|false|false|||consolidation
Finding|Functional Concept|SIMPLE_SEGMENT|7167,7171|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7167,7176|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7172,7176|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7172,7176|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7172,7176|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|7172,7176|false|false|false|C0740941|Lung Problem|lung
Event|Event|SIMPLE_SEGMENT|7178,7185|false|false|false|||thought
Finding|Idea or Concept|SIMPLE_SEGMENT|7178,7185|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|SIMPLE_SEGMENT|7178,7185|false|false|false|C0039869;C4319827|Thought|thought
Finding|Finding|SIMPLE_SEGMENT|7192,7200|false|false|false|C0332149|Possible|possibly
Drug|Organic Chemical|SIMPLE_SEGMENT|7201,7208|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|7201,7208|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|7201,7208|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|7201,7208|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7212,7221|false|false|false|C1720922|Respiratory Aspiration|aspirated
Event|Event|SIMPLE_SEGMENT|7212,7221|false|false|false|||aspirated
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7212,7221|false|false|false|C0700198|Pulmonary aspiration|aspirated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7222,7227|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|7222,7227|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|7222,7227|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7231,7238|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|SIMPLE_SEGMENT|7231,7238|false|false|false|C0728873|Monitor brand of insecticide|monitor
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7239,7252|false|false|false|C0523807|Oxygen saturation measurement|O2 saturation
Event|Event|SIMPLE_SEGMENT|7242,7252|false|false|false|||saturation
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7242,7252|false|false|false|C0522534|Saturated|saturation
Event|Event|SIMPLE_SEGMENT|7254,7265|false|false|false|||temperature
Procedure|Health Care Activity|SIMPLE_SEGMENT|7254,7265|false|false|false|C0886414|Body temperature measurement|temperature
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7267,7272|false|false|false|C4554533||trend
Anatomy|Cell|SIMPLE_SEGMENT|7273,7276|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|7273,7276|false|false|false|||WBC
Event|Event|SIMPLE_SEGMENT|7285,7293|false|false|false|||convered
Drug|Antibiotic|SIMPLE_SEGMENT|7300,7311|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|7300,7311|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|7318,7327|false|false|false|||inpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7318,7327|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|7318,7327|false|false|false|C1555324|inpatient encounter|inpatient
Event|Event|SIMPLE_SEGMENT|7343,7354|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7343,7354|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|SIMPLE_SEGMENT|7391,7403|false|false|false|||discontinued
Event|Event|SIMPLE_SEGMENT|7409,7418|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7409,7418|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7422,7427|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7422,7441|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7422,7441|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7428,7434|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7428,7434|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|SIMPLE_SEGMENT|7428,7434|false|false|false|||kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|7428,7434|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7428,7434|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7428,7434|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7428,7441|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7435,7441|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|7435,7441|false|false|false|||injury
Finding|Body Substance|SIMPLE_SEGMENT|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7450,7459|false|false|false|||presented
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7465,7475|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7465,7475|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7465,7475|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7465,7475|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7465,7475|false|false|false|C0201975|Creatinine measurement|creatinine
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7493,7503|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7493,7503|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7493,7503|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7493,7503|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7493,7503|false|false|false|C0201975|Creatinine measurement|creatinine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|7508,7511|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|7508,7511|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|7508,7511|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|SIMPLE_SEGMENT|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7529,7536|false|false|false|||unaware
Procedure|Research Activity|SIMPLE_SEGMENT|7529,7536|false|false|false|C0150114|unaware|unaware
Event|Event|SIMPLE_SEGMENT|7542,7549|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7542,7552|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|7542,7567|false|false|false|C0455686||history of kidney disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7553,7559|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7553,7559|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|7553,7559|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7553,7559|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7553,7559|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7553,7567|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7560,7567|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7560,7567|false|false|false|||disease
Finding|Body Substance|SIMPLE_SEGMENT|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|7586,7596|false|false|false|||discharged
Finding|Intellectual Product|SIMPLE_SEGMENT|7604,7610|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7611,7621|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|7611,7621|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|7611,7621|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|7611,7621|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7611,7621|false|false|false|C0201975|Creatinine measurement|creatinine
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7625,7652|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7636,7644|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7636,7652|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7645,7652|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7645,7652|false|false|false|||disease
Finding|Body Substance|SIMPLE_SEGMENT|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7667,7674|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7667,7677|true|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|7678,7681|true|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7678,7681|true|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7678,7681|true|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7678,7681|true|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|SIMPLE_SEGMENT|7678,7681|true|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7678,7681|true|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Event|Event|SIMPLE_SEGMENT|7678,7681|true|false|false|||AAA
Finding|Gene or Genome|SIMPLE_SEGMENT|7678,7681|true|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Event|Event|SIMPLE_SEGMENT|7682,7688|true|false|false|||repair
Finding|Functional Concept|SIMPLE_SEGMENT|7682,7688|true|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|SIMPLE_SEGMENT|7682,7688|true|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|SIMPLE_SEGMENT|7682,7688|true|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7682,7688|true|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|SIMPLE_SEGMENT|7704,7711|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7704,7714|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7723,7726|true|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7723,7726|true|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7723,7726|true|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7723,7726|true|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|7723,7726|true|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7723,7726|true|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|7723,7726|true|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7723,7726|true|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|7723,7726|true|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|7723,7726|true|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|7723,7726|true|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|SIMPLE_SEGMENT|7728,7735|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7728,7735|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7728,7735|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7736,7742|false|false|false|||denied
Event|Event|SIMPLE_SEGMENT|7743,7750|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|7743,7753|true|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|7754,7758|true|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7754,7758|true|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7762,7769|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|7762,7769|true|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|7782,7788|false|false|false|||stents
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7792,7799|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|7792,7799|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|SIMPLE_SEGMENT|7800,7807|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|7800,7807|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7800,7807|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|7812,7821|false|false|false|||continued
Finding|Idea or Concept|SIMPLE_SEGMENT|7826,7831|false|false|false|C1552828|Table Frame - above|above
Finding|Idea or Concept|SIMPLE_SEGMENT|7834,7846|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Classification|SIMPLE_SEGMENT|7855,7865|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7855,7865|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7866,7872|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|7866,7872|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7866,7872|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Event|Event|SIMPLE_SEGMENT|7866,7872|false|false|false|||stress
Finding|Finding|SIMPLE_SEGMENT|7866,7872|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7866,7877|false|false|false|C0920208|Echocardiography, Stress|stress echo
Event|Event|SIMPLE_SEGMENT|7873,7877|false|false|false|||echo
Procedure|Health Care Activity|SIMPLE_SEGMENT|7873,7877|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7873,7877|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Event|Event|SIMPLE_SEGMENT|7889,7899|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|7889,7899|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|7889,7899|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7900,7906|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7907,7910|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7907,7910|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7907,7910|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7911,7918|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7911,7918|false|false|false|||disease
Finding|Finding|SIMPLE_SEGMENT|7921,7929|false|false|false|C0332149|Possible|possibly
Finding|Gene or Genome|SIMPLE_SEGMENT|7932,7937|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Tissue|SIMPLE_SEGMENT|7938,7948|false|false|false|C0027061|Myocardium|myocardial
Event|Event|SIMPLE_SEGMENT|7949,7958|false|false|false|||territory
Event|Event|SIMPLE_SEGMENT|7962,7966|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|7962,7966|false|false|false|C0035647|Risk|risk
Finding|Functional Concept|SIMPLE_SEGMENT|7971,7977|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|SIMPLE_SEGMENT|7978,7992|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7978,7992|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|SIMPLE_SEGMENT|8009,8016|false|false|false|||monitor
Finding|Intellectual Product|SIMPLE_SEGMENT|8017,8021|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|8033,8042|false|false|false|||epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|8033,8042|false|false|false|C0014591|Epistaxis|epistaxis
Event|Event|SIMPLE_SEGMENT|8043,8050|false|false|false|||returns
Event|Event|SIMPLE_SEGMENT|8056,8059|false|false|false|||use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8074,8079|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|8074,8079|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|8074,8079|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8074,8085|false|false|false|C2608294|Nasal Spray brand of phenylephrine|nasal spray
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8080,8085|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|SIMPLE_SEGMENT|8080,8085|false|false|false|C2003858|Spray (action)|spray
Event|Event|SIMPLE_SEGMENT|8080,8085|false|false|false|||spray
Finding|Functional Concept|SIMPLE_SEGMENT|8080,8085|false|false|false|C4521772|Spray (administration method)|spray
Finding|Functional Concept|SIMPLE_SEGMENT|8088,8094|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8095,8100|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|8095,8100|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8095,8106|false|false|false|C0039985|Plain chest X-ray|chest x-ray
Event|Event|SIMPLE_SEGMENT|8101,8106|false|false|false|||x-ray
Finding|Functional Concept|SIMPLE_SEGMENT|8101,8106|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|SIMPLE_SEGMENT|8101,8106|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|8101,8106|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8101,8106|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Event|Event|SIMPLE_SEGMENT|8123,8129|false|false|false|||ensure
Event|Event|SIMPLE_SEGMENT|8130,8140|false|false|false|||resolution
Finding|Conceptual Entity|SIMPLE_SEGMENT|8130,8140|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|SIMPLE_SEGMENT|8130,8140|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8148,8151|false|false|false|C1261077|Structure of left lower lobe of lung|LLL
Event|Event|SIMPLE_SEGMENT|8153,8165|false|false|false|||infiltrative
Finding|Finding|SIMPLE_SEGMENT|8153,8165|false|false|false|C4527217|Infiltrative Tumor Margin|infiltrative
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8166,8173|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8166,8173|false|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|SIMPLE_SEGMENT|8166,8173|false|false|false|||process
Finding|Functional Concept|SIMPLE_SEGMENT|8166,8173|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8166,8173|false|false|false|C1522240|Process|process
Finding|Idea or Concept|SIMPLE_SEGMENT|8176,8184|false|false|false|C0750591|consider|Consider
Event|Event|SIMPLE_SEGMENT|8185,8191|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|8185,8191|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8185,8191|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8185,8194|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8185,8194|false|false|false|C1522577|follow-up|follow-up
Event|Event|SIMPLE_SEGMENT|8192,8194|false|false|false|||up
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8200,8203|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8200,8203|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|SIMPLE_SEGMENT|8200,8203|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|SIMPLE_SEGMENT|8200,8203|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Drug|Substance|SIMPLE_SEGMENT|8207,8214|false|false|false|C0032167|Plastics|Plastic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8207,8222|false|false|false|C0677616|Plastic Surgical Procedures|Plastic Surgery
Event|Event|SIMPLE_SEGMENT|8215,8222|false|false|false|||Surgery
Finding|Finding|SIMPLE_SEGMENT|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|SIMPLE_SEGMENT|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|SIMPLE_SEGMENT|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8215,8222|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Event|Event|SIMPLE_SEGMENT|8234,8244|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|8234,8244|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|8234,8244|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8248,8253|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|SIMPLE_SEGMENT|8248,8253|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|SIMPLE_SEGMENT|8248,8253|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8254,8263|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|8254,8263|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|8254,8263|false|false|false|C4554413|Fractured|fractures
Finding|Functional Concept|SIMPLE_SEGMENT|8266,8272|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Anatomy|Cell Component|SIMPLE_SEGMENT|8273,8276|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|SIMPLE_SEGMENT|8273,8276|false|false|false|||CBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8273,8276|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Intellectual Product|SIMPLE_SEGMENT|8284,8288|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|8292,8298|false|false|false|||ensure
Event|Event|SIMPLE_SEGMENT|8299,8308|false|false|false|||stability
Event|Event|SIMPLE_SEGMENT|8312,8315|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8312,8315|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8312,8315|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Anatomy|Cell|SIMPLE_SEGMENT|8321,8330|false|false|false|C0005821|Blood Platelets|platelets
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8321,8330|false|false|false|C0443116|Platelets Product|platelets
Event|Event|SIMPLE_SEGMENT|8321,8330|false|false|false|||platelets
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8321,8330|false|false|false|C0032181|Platelet count (procedure)|platelets
Finding|Idea or Concept|SIMPLE_SEGMENT|8333,8341|false|false|false|C0750591|consider|Consider
Event|Event|SIMPLE_SEGMENT|8342,8352|false|false|false|||conversion
Finding|Functional Concept|SIMPLE_SEGMENT|8342,8352|false|false|false|C0439836|Conversions (qualifier value)|conversion
Drug|Organic Chemical|SIMPLE_SEGMENT|8356,8366|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8356,8366|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8356,8375|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8356,8375|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8367,8375|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8367,8375|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|8367,8375|false|false|false|||tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8379,8388|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Finding|Mental Process|SIMPLE_SEGMENT|8394,8398|false|false|false|C1331418|Comfort|ease
Event|Event|SIMPLE_SEGMENT|8402,8416|false|false|false|||administration
Event|Occupational Activity|SIMPLE_SEGMENT|8402,8416|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8402,8416|false|false|false|C1533734|Administration (procedure)|administration
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8420,8431|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8420,8431|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8420,8431|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8420,8431|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|8420,8444|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|8435,8444|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8435,8444|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8463,8473|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8463,8473|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|8463,8478|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|8474,8478|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|8474,8478|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|8482,8490|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|8495,8503|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|8495,8503|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|8495,8503|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|8508,8519|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8508,8519|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|SIMPLE_SEGMENT|8550,8558|false|false|false|||Tartrate
Event|Event|SIMPLE_SEGMENT|8568,8571|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|8576,8587|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8576,8587|false|false|false|C0085542|pravastatin|Pravastatin
Event|Event|SIMPLE_SEGMENT|8597,8600|false|false|false|||QPM
Event|Event|SIMPLE_SEGMENT|8605,8614|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8605,8614|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|8605,8626|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8615,8626|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8615,8626|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|8615,8626|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8615,8626|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8631,8642|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8631,8642|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|8662,8675|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8662,8675|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|8662,8675|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8662,8675|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|8690,8693|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8694,8698|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|8694,8698|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|8694,8698|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|8694,8698|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|8707,8712|false|false|false|||avoid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8713,8718|false|false|false|C0003211;C3536840|Anti-Inflammatory Agents, Non-Steroidal|NSAID
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8719,8730|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8719,8730|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|8719,8730|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|8719,8730|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|SIMPLE_SEGMENT|8736,8745|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8736,8745|false|false|false|C0020740|ibuprofen|ibuprofen
Event|Event|SIMPLE_SEGMENT|8736,8745|false|false|false|||ibuprofen
Event|Event|SIMPLE_SEGMENT|8758,8766|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|8758,8766|false|false|false|C0019080|Hemorrhage|bleeding
Drug|Organic Chemical|SIMPLE_SEGMENT|8772,8779|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8772,8779|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8795,8803|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Drug|Organic Chemical|SIMPLE_SEGMENT|8817,8827|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8817,8827|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8817,8836|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8817,8836|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8828,8836|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8828,8836|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Event|Event|SIMPLE_SEGMENT|8828,8836|false|false|false|||Tartrate
Event|Event|SIMPLE_SEGMENT|8846,8849|false|false|false|||TID
Drug|Organic Chemical|SIMPLE_SEGMENT|8855,8865|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8855,8865|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|8855,8874|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8855,8874|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|8866,8874|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8866,8874|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Event|Event|SIMPLE_SEGMENT|8866,8874|false|false|false|||tartrate
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8883,8889|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|8893,8901|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8896,8901|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8896,8901|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8908,8913|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8932,8938|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|8939,8946|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|8939,8946|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|8953,8965|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8953,8965|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|8975,8978|false|false|false|||QPM
Event|Event|SIMPLE_SEGMENT|8980,8982|false|false|false|||RX
Drug|Organic Chemical|SIMPLE_SEGMENT|8984,8996|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8984,8996|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|8984,8996|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9005,9011|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|9015,9023|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9018,9023|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|9018,9023|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|9038,9042|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|9038,9042|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9049,9055|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|9056,9063|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9056,9063|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|9070,9083|false|false|false|C0030071|oxymetazoline|Oxymetazoline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9070,9083|false|false|false|C0030071|oxymetazoline|Oxymetazoline
Event|Event|SIMPLE_SEGMENT|9086,9090|false|false|false|||SPRY
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9094,9097|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9094,9097|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9094,9097|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9094,9097|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9094,9097|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|9098,9101|false|false|false|||PRN
Finding|Gene or Genome|SIMPLE_SEGMENT|9098,9101|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|9102,9111|false|false|false|||nosebleed
Event|Event|SIMPLE_SEGMENT|9125,9134|false|false|false|||purchased
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9144,9151|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|SIMPLE_SEGMENT|9144,9151|false|false|false|C0702263|Counter brand of Terbufos|counter
Event|Event|SIMPLE_SEGMENT|9144,9151|false|false|false|||counter
Finding|Intellectual Product|SIMPLE_SEGMENT|9157,9167|false|false|false|C0592503|Proprietary Name|brand name
Finding|Intellectual Product|SIMPLE_SEGMENT|9163,9167|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Event|Event|SIMPLE_SEGMENT|9181,9190|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9181,9190|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9181,9202|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|9181,9202|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9191,9202|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|9191,9202|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|9191,9202|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|9204,9208|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9204,9208|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9204,9208|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9204,9208|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|SIMPLE_SEGMENT|9214,9221|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|9214,9221|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|9224,9232|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9224,9232|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|9240,9249|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9240,9249|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9240,9259|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9250,9259|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9250,9259|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9250,9259|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9250,9259|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9250,9259|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9261,9266|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|9261,9266|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|9261,9266|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9261,9275|false|false|false|C0339848|Fractured nasal bones|Nasal fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|9267,9275|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|9267,9275|false|false|false|||fracture
Event|Event|SIMPLE_SEGMENT|9276,9285|false|false|false|||Epistaxis
Finding|Pathologic Function|SIMPLE_SEGMENT|9276,9285|false|false|false|C0014591|Epistaxis|Epistaxis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9286,9292|false|false|false|C4255010||NSTEMI
Event|Event|SIMPLE_SEGMENT|9286,9292|false|false|false|||NSTEMI
Finding|Finding|SIMPLE_SEGMENT|9286,9292|false|false|false|C3537184||NSTEMI
Event|Event|SIMPLE_SEGMENT|9296,9305|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9296,9305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9296,9305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9296,9305|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9296,9305|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9306,9315|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9306,9315|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9306,9315|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9306,9315|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9317,9323|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9317,9330|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9317,9330|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9324,9330|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9324,9330|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9332,9337|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9332,9337|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|9342,9350|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|9342,9350|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|9352,9357|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9352,9374|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9352,9374|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9361,9374|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9361,9374|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9361,9374|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9376,9381|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|9376,9381|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9376,9381|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|9376,9381|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|9386,9397|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|9386,9397|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|9399,9407|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9399,9407|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9399,9407|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9408,9414|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9408,9414|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9408,9414|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9416,9426|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9416,9426|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9429,9440|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|9429,9440|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|9429,9440|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|9445,9454|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9445,9454|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9445,9454|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9445,9454|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9445,9454|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9445,9467|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9445,9467|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9445,9467|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9455,9467|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9455,9467|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9455,9467|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|9487,9495|false|false|false|||admitted
Event|Event|SIMPLE_SEGMENT|9506,9510|false|false|false|||fell
Event|Event|SIMPLE_SEGMENT|9515,9520|false|false|false|||broke
Event|Event|SIMPLE_SEGMENT|9526,9530|false|false|false|||nose
Event|Event|SIMPLE_SEGMENT|9546,9552|false|false|false|||bleeds
Finding|Pathologic Function|SIMPLE_SEGMENT|9546,9552|false|false|false|C0019080|Hemorrhage|bleeds
Event|Event|SIMPLE_SEGMENT|9563,9572|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|9563,9572|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|9576,9583|false|false|false|||control
Event|Event|SIMPLE_SEGMENT|9602,9608|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|9625,9629|false|false|false|||stop
Event|Event|SIMPLE_SEGMENT|9634,9642|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|9634,9642|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|9656,9664|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|9656,9664|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|9683,9688|false|false|false|||found
Finding|Finding|SIMPLE_SEGMENT|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9702,9711|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9702,9711|false|false|false|C0041199|Troponin|troponins
Event|Event|SIMPLE_SEGMENT|9702,9711|false|false|false|||troponins
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9715,9720|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9715,9720|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9715,9720|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9715,9725|false|false|false|C0018941|Hematologic Tests|blood test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9721,9725|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|9721,9725|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|9721,9725|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|9721,9725|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9721,9725|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9721,9725|false|false|false|C0022885|Laboratory Procedures|test
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9735,9740|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9735,9740|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|9735,9740|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9735,9740|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|9744,9754|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|9744,9754|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|9744,9754|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9744,9754|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9763,9768|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9763,9768|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Event|Event|SIMPLE_SEGMENT|9763,9768|false|false|false|||heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|9763,9768|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|SIMPLE_SEGMENT|9796,9802|false|false|false|||follow
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|SIMPLE_SEGMENT|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|SIMPLE_SEGMENT|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|SIMPLE_SEGMENT|9816,9819|false|false|false|||PCP
Finding|Gene or Genome|SIMPLE_SEGMENT|9816,9819|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|SIMPLE_SEGMENT|9816,9819|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|SIMPLE_SEGMENT|9823,9830|false|false|false|||discuss
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9831,9837|false|false|true|C1718621|W stress|stress
Drug|Organic Chemical|SIMPLE_SEGMENT|9831,9837|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9831,9837|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|SIMPLE_SEGMENT|9831,9837|false|false|true|C0038435|Stress|stress
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9831,9842|false|false|true|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9838,9842|false|false|false|C4318744|Test - temporal region|test
Event|Event|SIMPLE_SEGMENT|9838,9842|false|false|false|||test
Finding|Functional Concept|SIMPLE_SEGMENT|9838,9842|false|false|true|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|SIMPLE_SEGMENT|9838,9842|false|false|true|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9838,9842|false|false|true|C0456984|Test Result|test
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9838,9842|false|false|true|C0022885|Laboratory Procedures|test
Event|Event|SIMPLE_SEGMENT|9854,9862|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|9854,9862|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|9854,9862|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|SIMPLE_SEGMENT|9863,9876|false|false|false|||participating
Event|Activity|SIMPLE_SEGMENT|9885,9889|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|9885,9889|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|9885,9889|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Activity|SIMPLE_SEGMENT|9906,9914|false|false|false|C1707391|Choose (action)|choosing
Procedure|Health Care Activity|SIMPLE_SEGMENT|9922,9930|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9931,9943|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9931,9943|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9931,9943|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

