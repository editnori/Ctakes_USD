 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
<EOL>|232,233
<EOL>|234,235
Shortness|252,261
of|262,264
breath|265,271
<EOL>|271,272
<EOL>|273,274
Major|274,279
Surgical|280,288
or|289,291
Invasive|292,300
Procedure|301,310
:|310,311
<EOL>|311,312
None|312,316
<EOL>|316,317
<EOL>|318,319
_|347,348
_|348,349
_|349,350
yo|351,353
woman|354,359
with|360,364
h|365,366
/|366,367
o|367,368
hypertension|369,381
,|381,382
hyperlipidemia|383,397
,|397,398
diabetes|399,407
<EOL>|408,409
mellitus|409,417
on|418,420
insulin|421,428
therapy|429,436
,|436,437
h|438,439
/|439,440
o|440,441
cerebellar|442,452
-|452,453
medullary|453,462
stroke|463,469
in|470,472
<EOL>|473,474
_|474,475
_|475,476
_|476,477
,|477,478
CKD|479,482
stage|483,488
III|489,492
-|492,493
IV|493,495
presenting|496,506
with|507,511
fatigue|512,519
and|520,523
dyspnea|524,531
on|532,534
<EOL>|535,536
exertion|536,544
(|545,546
DOE|546,549
)|549,550
for|551,554
a|555,556
few|557,560
weeks|561,566
,|566,567
markedly|568,576
worse|577,582
this|583,587
morning|588,595
.|595,596
<EOL>|597,598
Over|598,602
the|603,606
past|607,611
few|612,615
weeks|616,621
,|621,622
the|623,626
patient|627,634
noted|635,640
DOE|641,644
and|645,648
shortness|649,658
of|659,661
<EOL>|662,663
breath|663,669
(|670,671
SOB|671,674
)|674,675
even|676,680
at|681,683
rest|684,688
.|688,689
She|690,693
has|694,697
also|698,702
felt|703,707
more|708,712
tired|713,718
than|719,723
<EOL>|724,725
usual|725,730
.|730,731
She|732,735
notes|736,741
no|742,744
respiratory|745,756
issues|757,763
like|764,768
this|769,773
before|774,780
.|780,781
She|782,785
<EOL>|786,787
can|787,790
not|790,793
walk|794,798
up|799,801
stair|802,807
due|808,811
to|812,814
DOE|815,818
,|818,819
and|820,823
feels|824,829
SOB|830,833
after|834,839
only|840,844
a|845,846
<EOL>|847,848
short|848,853
distance|854,862
.|862,863
She|864,867
is|868,870
unsure|871,877
how|878,881
long|882,886
the|887,890
episodes|891,899
last|900,904
,|904,905
but|906,909
<EOL>|910,911
states|911,917
that|918,922
her|923,926
breathing|927,936
improves|937,945
with|946,950
albuterol|951,960
which|961,966
she|967,970
gets|971,975
<EOL>|976,977
from|977,981
her|982,985
husband|986,993
.|993,994
She|995,998
had|999,1002
a|1003,1004
bad|1005,1008
cough|1009,1014
around|1015,1021
a|1022,1023
month|1024,1029
ago|1030,1033
,|1033,1034
but|1035,1038
<EOL>|1039,1040
denies|1040,1046
any|1047,1050
recent|1051,1057
fevers|1058,1064
,|1064,1065
chills|1066,1072
,|1072,1073
or|1074,1076
night|1077,1082
sweats|1083,1089
.|1089,1090
No|1091,1093
chest|1094,1099
<EOL>|1100,1101
pain|1101,1105
,|1105,1106
nausea|1107,1113
,|1113,1114
or|1115,1117
dizziness|1118,1127
.|1127,1128
<EOL>|1128,1129
<EOL>|1130,1131
1.|1153,1155
CAD|1156,1159
RISK|1160,1164
FACTORS|1165,1172
:|1172,1173
+|1174,1175
Diabetes|1175,1183
,|1183,1184
+|1185,1186
Dyslipidemia|1186,1198
,|1198,1199
+|1200,1201
Hypertension|1201,1213
<EOL>|1213,1214
2.|1214,1216
CARDIAC|1217,1224
MI|1235,1237
in|1238,1240
_|1241,1242
_|1242,1243
_|1243,1244
<EOL>|1244,1245
3.|1245,1247
OTHER|1248,1253
PAST|1254,1258
MEDICAL|1259,1266
Hypertension|1278,1290
<EOL>|1290,1291
Hyperlipidemia|1291,1305
<EOL>|1305,1306
Diabetes|1306,1314
mellitus|1315,1323
on|1324,1326
insulin|1327,1334
therapy|1335,1342
<EOL>|1342,1343
h|1343,1344
/|1344,1345
o|1345,1346
cerebellar|1347,1357
-|1357,1358
medullary|1358,1367
stroke|1368,1374
in|1375,1377
_|1378,1379
_|1379,1380
_|1380,1381
<EOL>|1381,1382
CKD|1382,1385
stage|1386,1391
III|1392,1395
-|1395,1396
IV|1396,1398
<EOL>|1398,1399
PVD|1399,1402
<EOL>|1402,1403
<EOL>|1404,1405
:|1419,1420
<EOL>|1420,1421
_|1421,1422
_|1422,1423
_|1423,1424
<EOL>|1424,1425
:|1439,1440
<EOL>|1440,1441
Denies|1441,1447
cardiac|1448,1455
family|1456,1462
history|1463,1470
.|1470,1471
Family|1472,1478
hx|1479,1481
of|1482,1484
DM|1485,1487
and|1488,1491
HTN|1492,1495
;|1495,1496
<EOL>|1497,1498
otherwise|1498,1507
non-contributory|1508,1524
.|1524,1525
<EOL>|1525,1526
<EOL>|1527,1528
Admission|1543,1552
exam|1553,1557
:|1557,1558
<EOL>|1558,1559
GENERAL|1559,1566
-|1566,1567
Oriented|1568,1576
x3|1577,1579
.|1579,1580
Mood|1581,1585
,|1585,1586
affect|1587,1593
appropriate|1594,1605
.|1605,1606
<EOL>|1606,1607
VS|1607,1609
-|1609,1610
T|1611,1612
=|1612,1613
98.1|1614,1618
BP|1619,1621
=|1621,1622
200|1623,1626
/|1626,1627
103|1627,1630
HR|1631,1633
=|1633,1634
65|1635,1637
RR|1638,1640
=|1640,1641
26|1642,1644
O2|1645,1647
sat|1648,1651
=|1651,1652
100|1653,1656
%|1656,1657
on|1658,1660
RA|1661,1663
<EOL>|1663,1664
HEENT|1664,1669
-|1669,1670
NCAT|1671,1675
.|1675,1676
Sclera|1677,1683
anicteric|1684,1693
.|1693,1694
PERRL|1695,1700
,|1700,1701
EOMI|1702,1706
.|1706,1707
Conjunctiva|1708,1719
were|1720,1724
<EOL>|1725,1726
pink|1726,1730
,|1730,1731
no|1732,1734
pallor|1735,1741
or|1742,1744
cyanosis|1745,1753
of|1754,1756
the|1757,1760
oral|1761,1765
mucosa|1766,1772
.|1772,1773
No|1774,1776
xanthalesma|1777,1788
.|1788,1789
<EOL>|1789,1790
NECK|1790,1794
-|1794,1795
JVD|1796,1799
to|1800,1802
angle|1803,1808
of|1809,1811
mandible|1812,1820
<EOL>|1820,1821
CARDIAC|1821,1828
-|1828,1829
RR|1830,1832
,|1832,1833
normal|1834,1840
S1|1841,1843
,|1843,1844
S2|1845,1847
.|1847,1848
No|1849,1851
murmurs|1852,1859
,|1859,1860
rubs|1861,1865
or|1866,1868
gallops|1869,1876
.|1876,1877
No|1878,1880
<EOL>|1881,1882
thrills|1882,1889
,|1889,1890
lifts|1891,1896
.|1896,1897
<EOL>|1897,1898
LUNGS|1898,1903
-|1903,1904
Kyphosis|1905,1913
.|1913,1914
Resp|1915,1919
were|1920,1924
labored|1925,1932
,|1932,1933
mild|1934,1938
exp|1939,1942
wheezes|1943,1950
<EOL>|1951,1952
bilaterally|1952,1963
.|1963,1964
<EOL>|1964,1965
ABDOMEN|1965,1972
-|1972,1973
Soft|1974,1978
,|1978,1979
non-tender|1980,1990
,|1990,1991
not|1992,1995
distended|1996,2005
.|2005,2006
Abd|2007,2010
aorta|2011,2016
not|2017,2020
enlarged|2021,2029
<EOL>|2030,2031
by|2031,2033
palpation|2034,2043
.|2043,2044
No|2045,2047
abdominal|2048,2057
bruits|2058,2064
.|2064,2065
<EOL>|2065,2066
EXTREMITIES|2066,2077
-|2077,2078
No|2079,2081
clubbing|2082,2090
,|2090,2091
cyanosis|2092,2100
or|2101,2103
edema|2104,2109
.|2109,2110
No|2111,2113
femoral|2114,2121
bruits|2122,2128
.|2128,2129
<EOL>|2129,2130
SKIN|2130,2134
-|2134,2135
No|2136,2138
stasis|2139,2145
dermatitis|2146,2156
,|2156,2157
ulcers|2158,2164
,|2164,2165
scars|2166,2171
,|2171,2172
or|2173,2175
xanthomas|2176,2185
.|2185,2186
<EOL>|2186,2187
NEURO|2187,2192
-|2192,2193
CNII|2194,2198
-|2198,2199
XII|2199,2202
grossly|2203,2210
intact|2211,2217
.|2217,2218
Strength|2219,2227
_|2228,2229
_|2229,2230
_|2230,2231
in|2232,2234
LEs|2235,2238
and|2239,2242
UEs|2243,2246
.|2246,2247
<EOL>|2248,2249
Diminished|2249,2259
sensation|2260,2269
along|2270,2275
lateral|2276,2283
aspect|2284,2290
of|2291,2293
left|2294,2298
leg|2299,2302
to|2303,2305
light|2306,2311
<EOL>|2312,2313
touch|2313,2318
<EOL>|2318,2319
<EOL>|2319,2320
Discharge|2320,2329
exam|2330,2334
:|2334,2335
<EOL>|2335,2336
Lungs|2336,2341
:|2341,2342
CTAB|2343,2347
<EOL>|2347,2348
Otherwise|2348,2357
unchanged|2358,2367
<EOL>|2367,2368
<EOL>|2369,2370
Pertinent|2370,2379
Results|2380,2387
:|2387,2388
<EOL>|2388,2389
Admission|2389,2398
Labs|2399,2403
<EOL>|2403,2404
_|2404,2405
_|2405,2406
_|2406,2407
01|2408,2410
:|2410,2411
18PM|2411,2415
BLOOD|2416,2421
WBC|2422,2425
-|2425,2426
6|2426,2427
.|2427,2428
4|2428,2429
#|2429,2430
RBC|2431,2434
-|2434,2435
3|2435,2436
.|2436,2437
15|2437,2439
*|2439,2440
Hgb|2441,2444
-|2444,2445
9|2445,2446
.|2446,2447
5|2447,2448
*|2448,2449
Hct|2450,2453
-|2453,2454
30|2454,2456
.|2456,2457
1|2457,2458
*|2458,2459
<EOL>|2460,2461
MCV|2461,2464
-|2464,2465
96|2465,2467
MCH|2468,2471
-|2471,2472
30.1|2472,2476
MCHC|2477,2481
-|2481,2482
31.5|2482,2486
RDW|2487,2490
-|2490,2491
14.1|2491,2495
Plt|2496,2499
_|2500,2501
_|2501,2502
_|2502,2503
<EOL>|2503,2504
_|2504,2505
_|2505,2506
_|2506,2507
01|2508,2510
:|2510,2511
18PM|2511,2515
BLOOD|2516,2521
Glucose|2522,2529
-|2529,2530
150|2530,2533
*|2533,2534
UreaN|2535,2540
-|2540,2541
33|2541,2543
*|2543,2544
Creat|2545,2550
-|2550,2551
1|2551,2552
.|2552,2553
6|2553,2554
*|2554,2555
Na|2556,2558
-|2558,2559
144|2559,2562
<EOL>|2563,2564
K|2564,2565
-|2565,2566
4.8|2566,2569
Cl|2570,2572
-|2572,2573
111|2573,2576
*|2576,2577
HCO3|2578,2582
-|2582,2583
18|2583,2585
*|2585,2586
AnGap|2587,2592
-|2592,2593
20|2593,2595
<EOL>|2595,2596
_|2596,2597
_|2597,2598
_|2598,2599
01|2600,2602
:|2602,2603
18PM|2603,2607
BLOOD|2608,2613
CK|2614,2616
(|2616,2617
CPK|2617,2620
)|2620,2621
-|2621,2622
245|2622,2625
*|2625,2626
<EOL>|2626,2627
_|2627,2628
_|2628,2629
_|2629,2630
01|2631,2633
:|2633,2634
18PM|2634,2638
BLOOD|2639,2644
cTropnT|2645,2652
-|2652,2653
0|2653,2654
.|2654,2655
05|2655,2657
*|2657,2658
<EOL>|2658,2659
_|2659,2660
_|2660,2661
_|2661,2662
01|2663,2665
:|2665,2666
18PM|2666,2670
BLOOD|2671,2676
CK|2677,2679
-|2679,2680
MB|2680,2682
-|2682,2683
6|2683,2684
proBNP|2685,2691
-|2691,2692
4571|2692,2696
*|2696,2697
<EOL>|2697,2698
_|2698,2699
_|2699,2700
_|2700,2701
03|2702,2704
:|2704,2705
56AM|2705,2709
BLOOD|2710,2715
Calcium|2716,2723
-|2723,2724
9.4|2724,2727
Phos|2728,2732
-|2732,2733
4|2733,2734
.|2734,2735
9|2735,2736
*|2736,2737
Mg|2738,2740
-|2740,2741
2.0|2741,2744
Cholest|2745,2752
-|2752,2753
230|2753,2756
*|2756,2757
<EOL>|2757,2758
<EOL>|2758,2759
Pertinent|2759,2768
Labs|2769,2773
<EOL>|2773,2774
_|2774,2775
_|2775,2776
_|2776,2777
06|2778,2780
:|2780,2781
09AM|2781,2785
BLOOD|2786,2791
WBC|2792,2795
-|2795,2796
4.3|2796,2799
RBC|2800,2803
-|2803,2804
3|2804,2805
.|2805,2806
27|2806,2808
*|2808,2809
Hgb|2810,2813
-|2813,2814
9|2814,2815
.|2815,2816
9|2816,2817
*|2817,2818
Hct|2819,2822
-|2822,2823
31|2823,2825
.|2825,2826
4|2826,2827
*|2827,2828
<EOL>|2829,2830
MCV|2830,2833
-|2833,2834
96|2834,2836
MCH|2837,2840
-|2840,2841
30.4|2841,2845
MCHC|2846,2850
-|2850,2851
31.6|2851,2855
RDW|2856,2859
-|2859,2860
14.5|2860,2864
Plt|2865,2868
_|2869,2870
_|2870,2871
_|2871,2872
<EOL>|2872,2873
_|2873,2874
_|2874,2875
_|2875,2876
06|2877,2879
:|2879,2880
09AM|2880,2884
BLOOD|2885,2890
Glucose|2891,2898
-|2898,2899
138|2899,2902
*|2902,2903
UreaN|2904,2909
-|2909,2910
31|2910,2912
*|2912,2913
Creat|2914,2919
-|2919,2920
1|2920,2921
.|2921,2922
4|2922,2923
*|2923,2924
Na|2925,2927
-|2927,2928
144|2928,2931
<EOL>|2932,2933
K|2933,2934
-|2934,2935
4.3|2935,2938
Cl|2939,2941
-|2941,2942
107|2942,2945
HCO3|2946,2950
-|2950,2951
26|2951,2953
AnGap|2954,2959
-|2959,2960
15|2960,2962
<EOL>|2962,2963
<EOL>|2963,2964
_|2964,2965
_|2965,2966
_|2966,2967
06|2968,2970
:|2970,2971
09AM|2971,2975
BLOOD|2976,2981
ALT|2982,2985
-|2985,2986
20|2986,2988
AST|2989,2992
-|2992,2993
17|2993,2995
<EOL>|2995,2996
_|2996,2997
_|2997,2998
_|2998,2999
03|3000,3002
:|3002,3003
56AM|3003,3007
BLOOD|3008,3013
Triglyc|3014,3021
-|3021,3022
97|3022,3024
HDL|3025,3028
-|3028,3029
65|3029,3031
CHOL|3032,3036
/|3036,3037
HD|3037,3039
-|3039,3040
3.5|3040,3043
<EOL>|3044,3045
LDLcalc|3045,3052
-|3052,3053
146|3053,3056
*|3056,3057
<EOL>|3057,3058
_|3058,3059
_|3059,3060
_|3060,3061
03|3062,3064
:|3064,3065
56AM|3065,3069
BLOOD|3070,3075
%|3076,3077
HbA1c|3077,3082
-|3082,3083
8|3083,3084
.|3084,3085
1|3085,3086
*|3086,3087
eAG|3088,3091
-|3091,3092
186|3092,3095
*|3095,3096
<EOL>|3096,3097
<EOL>|3097,3098
_|3098,3099
_|3099,3100
_|3100,3101
01|3102,3104
:|3104,3105
18PM|3105,3109
BLOOD|3110,3115
CK|3116,3118
(|3118,3119
CPK|3119,3122
)|3122,3123
-|3123,3124
245|3124,3127
*|3127,3128
CK|3129,3131
-|3131,3132
MB|3132,3134
-|3134,3135
6|3135,3136
cTropnT|3137,3144
-|3144,3145
0|3145,3146
.|3146,3147
05|3147,3149
*|3149,3150
<EOL>|3150,3151
_|3151,3152
_|3152,3153
_|3153,3154
08|3155,3157
:|3157,3158
43PM|3158,3162
BLOOD|3163,3168
CK|3169,3171
(|3171,3172
CPK|3172,3175
)|3175,3176
-|3176,3177
198|3177,3180
CK|3182,3184
-|3184,3185
MB|3185,3187
-|3187,3188
5|3188,3189
cTropnT|3190,3197
-|3197,3198
0|3198,3199
.|3199,3200
03|3200,3202
*|3202,3203
<EOL>|3203,3204
_|3204,3205
_|3205,3206
_|3206,3207
03|3208,3210
:|3210,3211
56AM|3211,3215
BLOOD|3216,3221
CK|3222,3224
(|3224,3225
CPK|3225,3228
)|3228,3229
-|3229,3230
173|3230,3233
CK|3235,3237
-|3237,3238
MB|3238,3240
-|3240,3241
5|3241,3242
cTropnT|3243,3250
-|3250,3251
0|3251,3252
.|3252,3253
04|3253,3255
*|3255,3256
<EOL>|3256,3257
_|3257,3258
_|3258,3259
_|3259,3260
06|3261,3263
:|3263,3264
09AM|3264,3268
BLOOD|3269,3274
cTropnT|3296,3303
-|3303,3304
0|3304,3305
.|3305,3306
01|3306,3308
<EOL>|3308,3309
<EOL>|3309,3310
_|3310,3311
_|3311,3312
_|3312,3313
01|3314,3316
:|3316,3317
18PM|3317,3321
proBNP|3322,3328
-|3328,3329
4571|3329,3333
*|3333,3334
<EOL>|3334,3335
<EOL>|3335,3336
ECG|3336,3339
_|3340,3341
_|3341,3342
_|3342,3343
7|3345,3346
:|3346,3347
56|3347,3349
:|3349,3350
06|3350,3352
_|3353,3354
_|3354,3355
_|3355,3356
<EOL>|3358,3359
Baseline|3359,3367
artifact|3368,3376
.|3376,3377
Sinus|3378,3383
rhythm|3384,3390
.|3390,3391
The|3392,3395
Q|3396,3397
-|3397,3398
T|3398,3399
interval|3400,3408
is|3409,3411
400|3412,3415
<EOL>|3416,3417
milliseconds|3417,3429
.|3429,3430
Q|3431,3432
waves|3433,3438
in|3439,3441
leads|3442,3447
V1|3448,3450
-|3450,3451
V2|3451,3453
with|3454,3458
ST|3459,3461
-|3461,3462
T|3462,3463
wave|3464,3468
<EOL>|3469,3470
abnormalities|3470,3483
extending|3484,3493
to|3494,3496
lead|3497,3501
V6|3502,3504
.|3504,3505
Consider|3506,3514
prior|3515,3520
anterior|3521,3529
<EOL>|3530,3531
myocardial|3531,3541
infarction|3542,3552
.|3552,3553
Since|3554,3559
the|3560,3563
previous|3564,3572
tracing|3573,3580
of|3581,3583
_|3584,3585
_|3585,3586
_|3586,3587
<EOL>|3588,3589
atrial|3589,3595
premature|3596,3605
beats|3606,3611
are|3612,3615
not|3616,3619
seen|3620,3624
.|3624,3625
The|3626,3629
Q|3630,3631
-|3631,3632
T|3632,3633
interval|3634,3642
is|3643,3645
<EOL>|3646,3647
shorter|3647,3654
.|3654,3655
ST|3656,3658
-|3658,3659
T|3659,3660
wave|3661,3665
abnormalities|3666,3679
are|3680,3683
less|3684,3688
prominent|3689,3698
.|3698,3699
<EOL>|3701,3702
<EOL>|3703,3704
CXR|3704,3707
_|3708,3709
_|3709,3710
_|3710,3711
:|3711,3712
<EOL>|3712,3713
PA|3713,3715
and|3716,3719
lateral|3720,3727
views|3728,3733
of|3734,3736
the|3737,3740
chest|3741,3746
demonstrate|3747,3758
low|3759,3762
lung|3763,3767
volumes|3768,3775
.|3775,3776
<EOL>|3777,3778
Tiny|3778,3782
bilateral|3783,3792
pleural|3793,3800
effusions|3801,3810
are|3811,3814
new|3815,3818
since|3819,3824
_|3825,3826
_|3826,3827
_|3827,3828
.|3828,3829
No|3830,3832
<EOL>|3833,3834
signs|3834,3839
of|3840,3842
pneumonia|3843,3852
or|3853,3855
pulmonary|3856,3865
vascular|3866,3874
congestion|3875,3885
.|3885,3886
Heart|3887,3892
is|3893,3895
<EOL>|3896,3897
top|3897,3900
normal|3901,3907
in|3908,3910
size|3911,3915
though|3916,3922
this|3923,3927
is|3928,3930
stable|3931,3937
.|3937,3938
Aorta|3939,3944
is|3945,3947
markedly|3948,3956
<EOL>|3957,3958
tortuous|3958,3966
,|3966,3967
unchanged|3968,3977
.|3977,3978
Aortic|3979,3985
arch|3986,3990
calcifications|3991,4005
are|4006,4009
seen|4010,4014
.|4014,4015
There|4016,4021
<EOL>|4022,4023
is|4023,4025
no|4026,4028
pneumothorax|4029,4041
.|4041,4042
No|4043,4045
focal|4046,4051
consolidation|4052,4065
.|4065,4066
Partially|4067,4076
imaged|4077,4083
<EOL>|4084,4085
upper|4085,4090
abdomen|4091,4098
is|4099,4101
unremarkable|4102,4114
.|4114,4115
<EOL>|4115,4116
IMPRESSION|4116,4126
:|4126,4127
Tiny|4128,4132
pleural|4133,4140
effusions|4141,4150
,|4150,4151
new|4152,4155
.|4155,4156
Otherwise|4157,4166
unremarkable|4167,4179
.|4179,4180
<EOL>|4180,4181
<EOL>|4181,4182
ECHO|4182,4186
_|4187,4188
_|4188,4189
_|4189,4190
:|4190,4191
<EOL>|4191,4192
The|4192,4195
left|4196,4200
atrium|4201,4207
is|4208,4210
mildly|4211,4217
dilated|4218,4225
.|4225,4226
The|4227,4230
estimated|4231,4240
right|4241,4246
atrial|4247,4253
<EOL>|4254,4255
pressure|4255,4263
is|4264,4266
_|4267,4268
_|4268,4269
_|4269,4270
mmHg|4271,4275
.|4275,4276
Left|4277,4281
ventricular|4282,4293
wall|4294,4298
thickness|4299,4308
,|4308,4309
cavity|4310,4316
<EOL>|4317,4318
size|4318,4322
and|4323,4326
regional|4327,4335
/|4335,4336
global|4336,4342
systolic|4343,4351
function|4352,4360
are|4361,4364
normal|4365,4371
(|4372,4373
LVEF|4373,4377
<EOL>|4378,4379
>|4379,4380
55|4380,4382
%|4382,4383
)|4383,4384
.|4384,4385
Right|4386,4391
ventricular|4392,4403
chamber|4404,4411
size|4412,4416
and|4417,4420
free|4421,4425
wall|4426,4430
motion|4431,4437
are|4438,4441
<EOL>|4442,4443
normal|4443,4449
.|4449,4450
The|4451,4454
diameters|4455,4464
of|4465,4467
aorta|4468,4473
at|4474,4476
the|4477,4480
sinus|4481,4486
,|4486,4487
ascending|4488,4497
and|4498,4501
arch|4502,4506
<EOL>|4507,4508
levels|4508,4514
are|4515,4518
normal|4519,4525
.|4525,4526
The|4527,4530
aortic|4531,4537
valve|4538,4543
leaflets|4544,4552
(|4553,4554
3|4554,4555
)|4555,4556
are|4557,4560
mildly|4561,4567
<EOL>|4568,4569
thickened|4569,4578
but|4579,4582
aortic|4583,4589
stenosis|4590,4598
is|4599,4601
not|4602,4605
present|4606,4613
.|4613,4614
No|4615,4617
masses|4618,4624
or|4625,4627
<EOL>|4628,4629
vegetations|4629,4640
are|4641,4644
seen|4645,4649
on|4650,4652
the|4653,4656
aortic|4657,4663
valve|4664,4669
,|4669,4670
but|4671,4674
can|4675,4678
not|4678,4681
be|4682,4684
fully|4685,4690
<EOL>|4691,4692
excluded|4692,4700
due|4701,4704
to|4705,4707
suboptimal|4708,4718
image|4719,4724
quality|4725,4732
.|4732,4733
Trace|4734,4739
aortic|4740,4746
<EOL>|4747,4748
regurgitation|4748,4761
is|4762,4764
seen|4765,4769
.|4769,4770
The|4771,4774
mitral|4775,4781
valve|4782,4787
leaflets|4788,4796
are|4797,4800
<EOL>|4801,4802
structurally|4802,4814
normal|4815,4821
.|4821,4822
An|4823,4825
eccentric|4826,4835
,|4835,4836
anteriorly|4837,4847
directed|4848,4856
jet|4857,4860
of|4861,4863
<EOL>|4864,4865
mild|4865,4869
to|4870,4872
moderate|4873,4881
(|4882,4883
_|4883,4884
_|4884,4885
_|4885,4886
)|4886,4887
mitral|4888,4894
regurgitation|4895,4908
is|4909,4911
seen|4912,4916
.|4916,4917
Moderate|4918,4926
<EOL>|4927,4928
[|4928,4929
2|4929,4930
+|4930,4931
]|4931,4932
tricuspid|4933,4942
regurgitation|4943,4956
is|4957,4959
seen|4960,4964
.|4964,4965
There|4966,4971
is|4972,4974
moderate|4975,4983
<EOL>|4984,4985
pulmonary|4985,4994
artery|4995,5001
systolic|5002,5010
hypertension|5011,5023
.|5023,5024
The|5025,5028
end|5029,5032
-|5032,5033
diastolic|5033,5042
<EOL>|5043,5044
pulmonic|5044,5052
regurgitation|5053,5066
velocity|5067,5075
is|5076,5078
increased|5079,5088
suggesting|5089,5099
<EOL>|5100,5101
pulmonary|5101,5110
artery|5111,5117
diastolic|5118,5127
hypertension|5128,5140
.|5140,5141
There|5142,5147
is|5148,5150
an|5151,5153
anterior|5154,5162
<EOL>|5163,5164
space|5164,5169
which|5170,5175
most|5176,5180
likely|5181,5187
represents|5188,5198
a|5199,5200
prominent|5201,5210
fat|5211,5214
pad|5215,5218
.|5218,5219
<EOL>|5219,5220
IMPRESSION|5220,5230
:|5230,5231
Suboptimal|5232,5242
image|5243,5248
quality|5249,5256
.|5256,5257
Normal|5258,5264
biventricular|5265,5278
<EOL>|5279,5280
cavity|5280,5286
sizes|5287,5292
with|5293,5297
preserved|5298,5307
global|5308,5314
and|5315,5318
regional|5319,5327
biventricular|5328,5341
<EOL>|5342,5343
systolic|5343,5351
function|5352,5360
.|5360,5361
Pulmonary|5362,5371
artery|5372,5378
hypertension|5379,5391
.|5391,5392
Mild|5393,5397
-|5397,5398
moderate|5398,5406
<EOL>|5407,5408
mitral|5408,5414
regurgitation|5415,5428
.|5428,5429
Moderate|5430,5438
tricuspid|5439,5448
regurgitation|5449,5462
.|5462,5463
<EOL>|5464,5465
Compared|5465,5473
with|5474,5478
the|5479,5482
prior|5483,5488
study|5489,5494
(|5495,5496
images|5496,5502
reviewed|5503,5511
)|5511,5512
of|5513,5515
_|5516,5517
_|5517,5518
_|5518,5519
,|5519,5520
the|5521,5524
<EOL>|5525,5526
severity|5526,5534
of|5535,5537
mitral|5538,5544
and|5545,5548
tricuspid|5549,5558
regurgitation|5559,5572
are|5573,5576
increased|5577,5586
and|5587,5590
<EOL>|5591,5592
moderate|5592,5600
PA|5601,5603
hypertension|5604,5616
is|5617,5619
now|5620,5623
identified|5624,5634
.|5634,5635
<EOL>|5635,5636
<EOL>|5637,5638
_|5661,5662
_|5662,5663
_|5663,5664
woman|5665,5670
with|5671,5675
h|5676,5677
/|5677,5678
o|5678,5679
hypertension|5680,5692
,|5692,5693
hypelipidemia|5694,5707
,|5707,5708
diabetes|5709,5717
<EOL>|5718,5719
mellitus|5719,5727
on|5728,5730
insulin|5731,5738
,|5738,5739
cerebellar|5740,5750
-|5750,5751
medullary|5751,5760
stroke|5761,5767
in|5768,5770
_|5771,5772
_|5772,5773
_|5773,5774
,|5774,5775
<EOL>|5776,5777
stage|5777,5782
_|5783,5784
_|5784,5785
_|5785,5786
CKD|5787,5790
followed|5791,5799
by|5800,5802
Dr|5803,5805
_|5806,5807
_|5807,5808
_|5808,5809
presenting|5810,5820
with|5821,5825
fatigue|5826,5833
and|5834,5837
<EOL>|5838,5839
DOE|5839,5842
for|5843,5846
a|5847,5848
few|5849,5852
weeks|5853,5858
,|5858,5859
markedly|5860,5868
worse|5869,5874
the|5875,5878
morning|5879,5886
of|5887,5889
admission|5890,5899
.|5899,5900
<EOL>|5901,5902
The|5902,5905
patient|5906,5913
has|5914,5917
known|5918,5923
diastolic|5924,5933
dysfunction|5934,5945
.|5945,5946
Of|5947,5949
note|5950,5954
,|5954,5955
she|5956,5959
has|5960,5963
<EOL>|5964,5965
been|5965,5969
noncompliant|5970,5982
with|5983,5987
her|5988,5991
medications|5992,6003
at|6004,6006
home|6007,6011
.|6011,6012
On|6013,6015
arrival|6016,6023
to|6024,6026
<EOL>|6027,6028
the|6028,6031
floor|6032,6037
,|6037,6038
she|6039,6042
required|6043,6051
hydralazine|6052,6063
20|6064,6066
mg|6067,6069
to|6070,6072
bring|6073,6078
down|6079,6083
her|6084,6087
BP|6088,6090
.|6090,6091
<EOL>|6092,6093
She|6093,6096
has|6097,6100
likely|6101,6107
had|6108,6111
elevated|6112,6120
BPs|6121,6124
at|6125,6127
home|6128,6132
for|6133,6136
a|6137,6138
while|6139,6144
,|6144,6145
which|6146,6151
is|6152,6154
<EOL>|6155,6156
contributing|6156,6168
to|6169,6171
her|6172,6175
SOB|6176,6179
,|6179,6180
CHF|6181,6184
exacerbation|6185,6197
,|6197,6198
and|6199,6202
secondary|6203,6212
demand|6213,6219
<EOL>|6220,6221
myonecrosis|6221,6232
(|6233,6234
hypertensive|6234,6246
urgency|6247,6254
)|6254,6255
with|6256,6260
mildly|6261,6267
elevated|6268,6276
<EOL>|6277,6278
troponin|6278,6286
.|6286,6287
<EOL>|6287,6288
<EOL>|6288,6289
#|6289,6290
CAD|6291,6294
:|6294,6295
Although|6296,6304
she|6305,6308
did|6309,6312
not|6313,6316
have|6317,6321
a|6322,6323
classic|6324,6331
anginal|6332,6339
presentation|6340,6352
,|6352,6353
<EOL>|6354,6355
patient|6355,6362
has|6363,6366
several|6367,6374
risk|6375,6379
factors|6380,6387
for|6388,6391
acute|6392,6397
coronary|6398,6406
syndrome|6407,6415
.|6415,6416
<EOL>|6417,6418
Her|6418,6421
only|6422,6426
symptom|6427,6434
was|6435,6438
SOB|6439,6442
in|6443,6445
the|6446,6449
setting|6450,6457
of|6458,6460
elevated|6461,6469
BPs|6470,6473
<EOL>|6474,6475
attributed|6475,6485
to|6486,6488
medication|6489,6499
noncompliance|6500,6513
at|6514,6516
home|6517,6521
.|6521,6522
Her|6523,6526
troponin|6527,6535
<EOL>|6536,6537
fell|6537,6541
from|6542,6546
0.05|6547,6551
at|6552,6554
admission|6555,6564
to|6565,6567
0.01|6568,6572
at|6573,6575
discharge|6576,6585
in|6586,6588
the|6589,6592
setting|6593,6600
<EOL>|6601,6602
of|6602,6604
renal|6605,6610
dysfunction|6611,6622
,|6622,6623
but|6624,6627
there|6628,6633
was|6634,6637
not|6638,6641
a|6642,6643
clear|6644,6649
rise|6650,6654
and|6655,6658
fall|6659,6663
to|6664,6666
<EOL>|6667,6668
suggest|6668,6675
an|6676,6678
acute|6679,6684
infarction|6685,6695
from|6696,6700
plaque|6701,6707
rupture|6708,6715
and|6716,6719
thrombosis|6720,6730
.|6730,6731
<EOL>|6732,6733
She|6733,6736
was|6737,6740
scheduled|6741,6750
for|6751,6754
an|6755,6757
outpatient|6758,6768
stress|6769,6775
test|6776,6780
to|6781,6783
evaluate|6784,6792
for|6793,6796
<EOL>|6797,6798
evidence|6798,6806
of|6807,6809
ischemia|6810,6818
from|6819,6823
flow|6824,6828
-|6828,6829
limiting|6829,6837
CAD|6838,6841
.|6841,6842
We|6843,6845
decreased|6846,6855
ASA|6856,6859
to|6860,6862
<EOL>|6863,6864
81|6864,6866
mg|6867,6869
from|6870,6874
325|6875,6878
mg|6879,6881
daily|6882,6887
to|6888,6890
decrease|6891,6899
the|6900,6903
risk|6904,6908
of|6909,6911
bleeding|6912,6920
.|6920,6921
Her|6922,6925
<EOL>|6926,6927
LDL|6927,6930
was|6931,6934
found|6935,6940
to|6941,6943
be|6944,6946
146|6947,6950
.|6950,6951
We|6952,6954
wanted|6955,6961
to|6962,6964
change|6965,6971
her|6972,6975
from|6976,6980
<EOL>|6981,6982
simvastatin|6982,6993
to|6994,6996
the|6997,7000
more|7001,7005
potent|7006,7012
atorvastatin|7013,7025
(|7026,7027
and|7027,7030
avoid|7031,7036
issues|7037,7043
<EOL>|7044,7045
with|7045,7049
drug|7050,7054
-|7054,7055
drug|7055,7059
interactions|7060,7072
)|7072,7073
,|7073,7074
but|7075,7078
her|7079,7082
insurance|7083,7092
would|7093,7098
not|7099,7102
cover|7103,7108
<EOL>|7109,7110
atorvastatin|7110,7122
.|7122,7123
She|7124,7127
was|7128,7131
therefore|7132,7141
switched|7142,7150
to|7151,7153
pravastatin|7154,7165
80|7166,7168
mg|7169,7171
at|7172,7174
<EOL>|7175,7176
discharge|7176,7185
.|7185,7186
From|7187,7191
a|7192,7193
cardiac|7194,7201
standpoint|7202,7212
,|7212,7213
we|7214,7216
did|7217,7220
not|7221,7224
feel|7225,7229
that|7230,7234
<EOL>|7235,7236
Plavix|7236,7242
was|7243,7246
necessary|7247,7256
for|7257,7260
CAD|7261,7264
,|7264,7265
but|7266,7269
her|7270,7273
neurologist|7274,7285
was|7286,7289
contacted|7290,7299
<EOL>|7300,7301
and|7301,7304
wanted|7305,7311
Plavix|7312,7318
continued|7319,7328
.|7328,7329
We|7330,7332
had|7333,7336
to|7337,7339
stop|7340,7344
metoprolol|7345,7355
due|7356,7359
to|7360,7362
HR|7363,7365
<EOL>|7366,7367
in|7367,7369
the|7370,7373
_|7374,7375
_|7375,7376
_|7376,7377
during|7378,7384
admission|7385,7394
even|7395,7399
off|7400,7403
metoprolol|7404,7414
.|7414,7415
<EOL>|7415,7416
<EOL>|7418,7419
#|7419,7420
Pump|7421,7425
:|7425,7426
Last|7427,7431
echo|7432,7436
in|7437,7439
_|7440,7441
_|7441,7442
_|7442,7443
showed|7444,7450
low|7451,7454
normal|7455,7461
LVEF|7462,7466
.|7466,7467
Her|7468,7471
current|7472,7479
<EOL>|7480,7481
presentation|7481,7493
was|7494,7497
consistent|7498,7508
with|7509,7513
CHF|7514,7517
exacerbation|7518,7530
with|7531,7535
bilateral|7536,7545
<EOL>|7546,7547
pleural|7547,7554
effusions|7555,7564
,|7564,7565
dyspnea|7566,7573
,|7573,7574
and|7575,7578
elevated|7579,7587
NT|7588,7590
-|7590,7591
Pro-BNP|7591,7598
.|7598,7599
Her|7600,7603
TTE|7604,7607
<EOL>|7608,7609
showed|7609,7615
mild|7616,7620
-|7620,7621
moderate|7621,7629
mitral|7630,7636
and|7637,7640
moderate|7641,7649
tricuspid|7650,7659
<EOL>|7660,7661
regurgitation|7661,7674
,|7674,7675
LVEF|7676,7680
50|7681,7683
-|7683,7684
55|7684,7686
%|7686,7687
,|7687,7688
and|7689,7692
pulmonary|7693,7702
hypertension|7703,7715
.|7715,7716
We|7717,7719
<EOL>|7720,7721
changed|7721,7728
her|7729,7732
HCTZ|7733,7737
to|7738,7740
Lasix|7741,7746
40|7747,7749
mg|7750,7752
PO|7753,7755
at|7756,7758
discharge|7759,7768
.|7768,7769
This|7770,7774
medication|7775,7785
<EOL>|7786,7787
can|7787,7790
be|7791,7793
uptitrated|7794,7804
as|7805,7807
needed|7808,7814
.|7814,7815
<EOL>|7815,7816
<EOL>|7816,7817
#|7817,7818
Hypertension|7819,7831
:|7831,7832
The|7833,7836
patient|7837,7844
's|7844,7846
nephrologist|7847,7859
,|7859,7860
Dr.|7861,7864
_|7865,7866
_|7866,7867
_|7867,7868
,|7868,7869
agreed|7870,7876
<EOL>|7877,7878
with|7878,7882
our|7883,7886
proposed|7887,7895
medication|7896,7906
adjustments|7907,7918
,|7918,7919
but|7920,7923
recommended|7924,7935
<EOL>|7936,7937
staying|7937,7944
away|7945,7949
from|7950,7954
clonidine|7955,7964
.|7964,7965
There|7966,7971
has|7972,7975
been|7976,7980
a|7981,7982
H|7983,7984
/|7984,7985
O|7985,7986
medication|7987,7997
<EOL>|7998,7999
non-adherence|7999,8012
.|8012,8013
Social|8014,8020
work|8021,8025
was|8026,8029
involved|8030,8038
in|8039,8041
discharge|8042,8051
planning|8052,8060
,|8060,8061
<EOL>|8062,8063
and|8063,8066
_|8067,8068
_|8068,8069
_|8069,8070
will|8071,8075
be|8076,8078
assisting|8079,8088
the|8089,8092
patient|8093,8100
at|8101,8103
home|8104,8108
.|8108,8109
We|8110,8112
added|8113,8118
<EOL>|8119,8120
lisinopril|8120,8130
20|8131,8133
mg|8134,8136
daily|8137,8142
,|8142,8143
Lasix|8144,8149
40|8150,8152
mg|8153,8155
daily|8156,8161
and|8162,8165
continued|8166,8175
<EOL>|8176,8177
nifedipine|8177,8187
120|8188,8191
mg|8192,8194
daily|8195,8200
.|8200,8201
Her|8202,8205
atenolol|8206,8214
was|8215,8218
stopped|8219,8226
due|8227,8230
to|8231,8233
her|8234,8237
<EOL>|8238,8239
renal|8239,8244
dysfunction|8245,8256
,|8256,8257
but|8258,8261
her|8262,8265
metoprolol|8266,8276
had|8277,8280
to|8281,8283
be|8284,8286
stopped|8287,8294
due|8295,8298
to|8299,8301
<EOL>|8302,8303
bradycardia|8303,8314
.|8314,8315
She|8316,8319
should|8320,8326
continue|8327,8335
on|8336,8338
once|8339,8343
a|8344,8345
day|8346,8349
medication|8350,8360
dosing|8361,8367
<EOL>|8368,8369
to|8369,8371
help|8372,8376
with|8377,8381
compliance|8382,8392
.|8392,8393
<EOL>|8393,8394
<EOL>|8394,8395
#|8395,8396
?|8397,8398
COPD|8399,8403
:|8403,8404
The|8405,8408
patient|8409,8416
may|8417,8420
have|8421,8425
a|8426,8427
component|8428,8437
of|8438,8440
COPD|8441,8445
as|8446,8448
she|8449,8452
was|8453,8456
<EOL>|8457,8458
wheezing|8458,8466
on|8467,8469
admission|8470,8479
and|8480,8483
responded|8484,8493
to|8494,8496
albuterol|8497,8506
.|8506,8507
She|8508,8511
was|8512,8515
given|8516,8521
<EOL>|8522,8523
a|8523,8524
prescription|8525,8537
for|8538,8541
albuterol|8542,8551
prn|8552,8555
.|8555,8556
<EOL>|8556,8557
<EOL>|8557,8558
Transitional|8558,8570
Issues|8571,8577
:|8577,8578
<EOL>|8578,8579
-|8579,8580
She|8581,8584
will|8585,8589
be|8590,8592
scheduled|8593,8602
for|8603,8606
outpt|8607,8612
stress|8613,8619
stress|8620,8626
test|8627,8631
<EOL>|8631,8632
-|8632,8633
She|8634,8637
has|8638,8641
follow|8642,8648
-|8648,8649
up|8649,8651
appointments|8652,8664
with|8665,8669
Dr.|8670,8673
_|8674,8675
_|8675,8676
_|8676,8677
and|8678,8681
Dr|8682,8684
.|8684,8685
<EOL>|8686,8687
_|8687,8688
_|8688,8689
_|8689,8690
and|8691,8694
both|8695,8699
can|8700,8703
work|8704,8708
on|8709,8711
uptitrating|8712,8723
her|8724,8727
BP|8728,8730
<EOL>|8731,8732
meds|8732,8736
as|8737,8739
needed|8740,8746
.|8746,8747
<EOL>|8747,8748
-|8748,8749
_|8750,8751
_|8751,8752
_|8752,8753
will|8754,8758
need|8759,8763
to|8764,8766
work|8767,8771
with|8772,8776
patient|8777,8784
on|8785,8787
medication|8788,8798
compliance|8799,8809
.|8809,8810
<EOL>|8810,8811
<EOL>|8812,8813
Medications|8813,8824
on|8825,8827
Admission|8828,8837
:|8837,8838
<EOL>|8838,8839
ATENOLOL|8839,8847
-|8848,8849
100|8850,8853
mg|8854,8856
Tablet|8857,8863
-|8864,8865
1.5|8866,8869
Tablet|8870,8876
(|8876,8877
s|8877,8878
)|8878,8879
by|8880,8882
mouth|8883,8888
once|8889,8893
a|8894,8895
day|8896,8899
<EOL>|8900,8901
CLONIDINE|8901,8910
-|8911,8912
0.1|8913,8916
mg|8917,8919
/|8919,8920
24|8920,8922
hour|8923,8927
Patch|8928,8933
Weekly|8934,8940
-|8941,8942
place|8943,8948
on|8949,8951
shoulder|8952,8960
once|8961,8965
<EOL>|8966,8967
a|8967,8968
week|8969,8973
<EOL>|8973,8974
CLOPIDOGREL|8974,8985
[|8986,8987
PLAVIX|8987,8993
]|8993,8994
-|8995,8996
75|8997,8999
mg|9000,9002
Tablet|9003,9009
-|9010,9011
1|9012,9013
Tablet|9014,9020
(|9020,9021
s|9021,9022
)|9022,9023
by|9024,9026
mouth|9027,9032
once|9033,9037
<EOL>|9038,9039
a|9039,9040
day|9041,9044
generic|9045,9052
is|9053,9055
available|9056,9065
preferable|9066,9076
,|9076,9077
please|9078,9084
call|9085,9089
Dr|9090,9092
_|9093,9094
_|9094,9095
_|9095,9096
<EOL>|9097,9098
an|9098,9100
appointment|9101,9112
<EOL>|9114,9115
FENOFIBRATE|9115,9126
MICRONIZED|9127,9137
-|9138,9139
134|9140,9143
mg|9144,9146
Capsule|9147,9154
-|9155,9156
1|9157,9158
Capsule|9159,9166
(|9166,9167
s|9167,9168
)|9168,9169
by|9170,9172
mouth|9173,9178
<EOL>|9179,9180
once|9180,9184
a|9185,9186
day|9187,9190
<EOL>|9190,9191
HYDROCHLOROTHIAZIDE|9191,9210
-|9211,9212
25|9213,9215
mg|9216,9218
Tablet|9219,9225
-|9226,9227
1|9228,9229
(|9230,9231
One|9231,9234
)|9234,9235
Tablet|9236,9242
(|9242,9243
s|9243,9244
)|9244,9245
by|9246,9248
mouth|9249,9254
<EOL>|9255,9256
once|9256,9260
a|9261,9262
day|9263,9266
<EOL>|9266,9267
NIFEDIPINE|9267,9277
[|9278,9279
NIFEDIAC|9279,9287
CC|9288,9290
]|9290,9291
-|9292,9293
60|9294,9296
mg|9297,9299
Tablet|9300,9306
Extended|9307,9315
Release|9316,9323
-|9324,9325
2|9326,9327
<EOL>|9328,9329
Tablet|9329,9335
(|9335,9336
s|9336,9337
)|9337,9338
by|9339,9341
mouth|9342,9347
once|9348,9352
a|9353,9354
day|9355,9358
<EOL>|9358,9359
NITROGLYCERIN|9359,9372
[|9373,9374
NITROSTAT|9374,9383
]|9383,9384
-|9385,9386
0.3|9387,9390
mg|9391,9393
Tablet|9394,9400
,|9400,9401
Sublingual|9402,9412
-|9413,9414
1|9415,9416
<EOL>|9417,9418
Tablet|9418,9424
(|9424,9425
s|9425,9426
)|9426,9427
sublingually|9428,9440
sl|9441,9443
as|9444,9446
needed|9447,9453
for|9454,9457
prn|9458,9461
chest|9462,9467
pain|9468,9472
may|9473,9476
use|9477,9480
3|9481,9482
<EOL>|9483,9484
doses|9484,9489
,|9489,9490
5|9491,9492
minutes|9493,9500
apart|9501,9506
;|9506,9507
if|9508,9510
no|9511,9513
relief|9514,9520
,|9520,9521
ED|9522,9524
visit|9525,9530
<EOL>|9531,9532
RANITIDINE|9532,9542
HCL|9543,9546
-|9547,9548
300|9549,9552
mg|9553,9555
Tablet|9556,9562
-|9563,9564
1|9565,9566
Tablet|9567,9573
(|9573,9574
s|9574,9575
)|9575,9576
by|9577,9579
mouth|9580,9585
once|9586,9590
a|9591,9592
day|9593,9596
<EOL>|9596,9597
SIMVASTATIN|9597,9608
-|9609,9610
80|9611,9613
mg|9614,9616
Tablet|9617,9623
-|9624,9625
1|9626,9627
Tablet|9628,9634
(|9634,9635
s|9635,9636
)|9636,9637
by|9638,9640
mouth|9641,9646
at|9647,9649
bedtime|9650,9657
<EOL>|9657,9658
<EOL>|9658,9659
Medications|9659,9670
-|9671,9672
OTC|9673,9676
<EOL>|9678,9679
ASPIRIN|9679,9686
[|9687,9688
ENTERIC|9688,9695
COATED|9696,9702
ASPIRIN|9703,9710
]|9710,9711
-|9712,9713
325|9714,9717
mg|9718,9720
Tablet|9721,9727
,|9727,9728
Delayed|9729,9736
<EOL>|9737,9738
Release|9738,9745
(|9746,9747
E.C|9747,9750
.|9750,9751
)|9751,9752
-|9753,9754
1|9755,9756
(|9757,9758
One|9758,9761
)|9761,9762
Tablet|9763,9769
(|9769,9770
s|9770,9771
)|9771,9772
by|9773,9775
mouth|9776,9781
once|9782,9786
a|9787,9788
day|9789,9792
<EOL>|9792,9793
INSULIN|9793,9800
NPH|9801,9804
&|9805,9806
REGULAR|9807,9814
HUMAN|9815,9820
[|9821,9822
HUMULIN|9822,9829
70|9830,9832
/|9832,9833
30|9833,9835
]|9835,9836
-|9837,9838
100|9839,9842
unit|9843,9847
/|9847,9848
mL|9848,9850
<EOL>|9851,9852
(|9852,9853
70|9853,9855
-|9855,9856
30|9856,9858
)|9858,9859
Suspension|9860,9870
-|9871,9872
30|9873,9875
units|9876,9881
at|9882,9884
dinner|9885,9891
at|9892,9894
dinner|9895,9901
<EOL>|9901,9902
MULTIVITAMIN|9902,9914
-|9915,9916
(|9917,9918
OTC|9918,9921
)|9921,9922
-|9923,9924
Tablet|9925,9931
-|9932,9933
1|9934,9935
Tablet|9936,9942
(|9942,9943
s|9943,9944
)|9944,9945
by|9946,9948
mouth|9949,9954
once|9955,9959
a|9960,9961
day|9962,9965
<EOL>|9965,9966
<EOL>|9967,9968
Discharge|9968,9977
Medications|9978,9989
:|9989,9990
<EOL>|9990,9991
1.|9991,9993
clopidogrel|9994,10005
75|10006,10008
mg|10009,10011
Tablet|10012,10018
Sig|10019,10022
:|10022,10023
One|10024,10027
(|10028,10029
1|10029,10030
)|10030,10031
Tablet|10032,10038
PO|10039,10041
DAILY|10042,10047
<EOL>|10048,10049
(|10049,10050
Daily|10050,10055
)|10055,10056
.|10056,10057
Disp|10058,10062
:|10062,10063
*|10063,10064
30|10064,10066
Tablet|10067,10073
(|10073,10074
s|10074,10075
)|10075,10076
*|10076,10077
Refills|10078,10085
:|10085,10086
*|10086,10087
2|10087,10088
*|10088,10089
<EOL>|10089,10090
2.|10090,10092
nitroglycerin|10093,10106
0.4|10107,10110
mg|10111,10113
Tablet|10114,10120
,|10120,10121
Sublingual|10122,10132
Sig|10133,10136
:|10136,10137
One|10138,10141
(|10142,10143
1|10143,10144
)|10144,10145
Tablet|10146,10152
,|10152,10153
<EOL>|10154,10155
Sublingual|10155,10165
Sublingual|10166,10176
PRN|10177,10180
(|10181,10182
as|10182,10184
needed|10185,10191
)|10191,10192
as|10193,10195
needed|10196,10202
for|10203,10206
chest|10207,10212
pain|10213,10217
:|10217,10218
<EOL>|10219,10220
may|10220,10223
take|10224,10228
up|10229,10231
to|10232,10234
3|10235,10236
over|10237,10241
15|10242,10244
minutes|10245,10252
.|10252,10253
Disp|10254,10258
:|10258,10259
*|10259,10260
30|10260,10262
Tablet|10263,10269
,|10269,10270
<EOL>|10271,10272
Sublingual|10272,10282
(|10282,10283
s|10283,10284
)|10284,10285
*|10285,10286
Refills|10287,10294
:|10294,10295
*|10295,10296
0|10296,10297
*|10297,10298
<EOL>|10298,10299
3.|10299,10301
multivitamin|10302,10314
Tablet|10319,10325
Sig|10326,10329
:|10329,10330
One|10331,10334
(|10335,10336
1|10336,10337
)|10337,10338
Tablet|10339,10345
PO|10346,10348
DAILY|10349,10354
(|10355,10356
Daily|10356,10361
)|10361,10362
.|10362,10363
<EOL>|10364,10365
Disp|10365,10369
:|10369,10370
*|10370,10371
30|10371,10373
Tablet|10374,10380
(|10380,10381
s|10381,10382
)|10382,10383
*|10383,10384
Refills|10385,10392
:|10392,10393
*|10393,10394
2|10394,10395
*|10395,10396
<EOL>|10396,10397
4.|10397,10399
ranitidine|10400,10410
HCl|10411,10414
150|10415,10418
mg|10419,10421
Tablet|10422,10428
Sig|10429,10432
:|10432,10433
Two|10434,10437
(|10438,10439
2|10439,10440
)|10440,10441
Tablet|10442,10448
PO|10449,10451
DAILY|10452,10457
<EOL>|10458,10459
(|10459,10460
Daily|10460,10465
)|10465,10466
.|10466,10467
Disp|10468,10472
:|10472,10473
*|10473,10474
60|10474,10476
Tablet|10477,10483
(|10483,10484
s|10484,10485
)|10485,10486
*|10486,10487
Refills|10488,10495
:|10495,10496
*|10496,10497
2|10497,10498
*|10498,10499
<EOL>|10499,10500
5.|10500,10502
pravastatin|10503,10514
80|10515,10517
mg|10518,10520
Tablet|10521,10527
Sig|10528,10531
:|10531,10532
One|10533,10536
(|10537,10538
1|10538,10539
)|10539,10540
Tablet|10541,10547
PO|10548,10550
DAILY|10551,10556
<EOL>|10557,10558
(|10558,10559
Daily|10559,10564
)|10564,10565
.|10565,10566
Disp|10567,10571
:|10571,10572
*|10572,10573
30|10573,10575
Tablet|10576,10582
(|10582,10583
s|10583,10584
)|10584,10585
*|10585,10586
Refills|10587,10594
:|10594,10595
*|10595,10596
2|10596,10597
*|10597,10598
<EOL>|10598,10599
6.|10599,10601
aspirin|10602,10609
81|10610,10612
mg|10613,10615
Tablet|10616,10622
,|10622,10623
Chewable|10624,10632
Sig|10633,10636
:|10636,10637
One|10638,10641
(|10642,10643
1|10643,10644
)|10644,10645
Tablet|10646,10652
,|10652,10653
Chewable|10654,10662
<EOL>|10663,10664
PO|10664,10666
DAILY|10667,10672
(|10673,10674
Daily|10674,10679
)|10679,10680
.|10680,10681
Disp|10682,10686
:|10686,10687
*|10687,10688
30|10688,10690
Tablet|10691,10697
,|10697,10698
Chewable|10699,10707
(|10707,10708
s|10708,10709
)|10709,10710
*|10710,10711
Refills|10712,10719
:|10719,10720
*|10720,10721
2|10721,10722
*|10722,10723
<EOL>|10723,10724
7.|10724,10726
lisinopril|10727,10737
20|10738,10740
mg|10741,10743
Tablet|10744,10750
Sig|10751,10754
:|10754,10755
One|10756,10759
(|10760,10761
1|10761,10762
)|10762,10763
Tablet|10764,10770
PO|10771,10773
DAILY|10774,10779
(|10780,10781
Daily|10781,10786
)|10786,10787
.|10787,10788
<EOL>|10789,10790
Disp|10790,10794
:|10794,10795
*|10795,10796
30|10796,10798
Tablet|10799,10805
(|10805,10806
s|10806,10807
)|10807,10808
*|10808,10809
Refills|10810,10817
:|10817,10818
*|10818,10819
2|10819,10820
*|10820,10821
<EOL>|10821,10822
8.|10822,10824
nifedipine|10825,10835
60|10836,10838
mg|10839,10841
Tablet|10842,10848
Extended|10849,10857
Release|10858,10865
Sig|10866,10869
:|10869,10870
Two|10871,10874
(|10875,10876
2|10876,10877
)|10877,10878
Tablet|10879,10885
<EOL>|10886,10887
Extended|10887,10895
Release|10896,10903
PO|10904,10906
DAILY|10907,10912
(|10913,10914
Daily|10914,10919
)|10919,10920
.|10920,10921
Disp|10922,10926
:|10926,10927
*|10927,10928
30|10928,10930
Tablet|10931,10937
Extended|10938,10946
<EOL>|10947,10948
Release|10948,10955
(|10955,10956
s|10956,10957
)|10957,10958
*|10958,10959
Refills|10960,10967
:|10967,10968
*|10968,10969
2|10969,10970
*|10970,10971
<EOL>|10971,10972
9.|10972,10974
furosemide|10975,10985
40|10986,10988
mg|10989,10991
Tablet|10992,10998
Sig|10999,11002
:|11002,11003
One|11004,11007
(|11008,11009
1|11009,11010
)|11010,11011
Tablet|11012,11018
PO|11019,11021
DAILY|11022,11027
(|11028,11029
Daily|11029,11034
)|11034,11035
.|11035,11036
<EOL>|11037,11038
Disp|11038,11042
:|11042,11043
*|11043,11044
30|11044,11046
Tablet|11047,11053
(|11053,11054
s|11054,11055
)|11055,11056
*|11056,11057
Refills|11058,11065
:|11065,11066
*|11066,11067
2|11067,11068
*|11068,11069
<EOL>|11069,11070
10.|11070,11073
insulin|11074,11081
NPH|11082,11085
&|11086,11087
regular|11088,11095
human|11096,11101
100|11102,11105
unit|11106,11110
/|11110,11111
mL|11111,11113
(|11114,11115
70|11115,11117
-|11117,11118
30|11118,11120
)|11120,11121
Insulin|11122,11129
Pen|11130,11133
<EOL>|11134,11135
Sig|11135,11138
:|11138,11139
Thirty|11140,11146
(|11147,11148
30|11148,11150
)|11150,11151
units|11152,11157
Subcutaneous|11158,11170
at|11171,11173
dinner.|11174,11181
Disp|11182,11186
:|11186,11187
*|11187,11188
900|11188,11191
units|11192,11197
*|11197,11198
<EOL>|11199,11200
Refills|11200,11207
:|11207,11208
*|11208,11209
2|11209,11210
*|11210,11211
<EOL>|11211,11212
11.|11212,11215
albuterol|11216,11225
sulfate|11226,11233
90|11234,11236
mcg|11237,11240
/|11240,11241
actuation|11241,11250
HFA|11251,11254
Aerosol|11255,11262
Inhaler|11263,11270
Sig|11271,11274
:|11274,11275
<EOL>|11276,11277
_|11277,11278
_|11278,11279
_|11279,11280
puffs|11281,11286
Inhalation|11287,11297
every|11298,11303
_|11304,11305
_|11305,11306
_|11306,11307
hours|11308,11313
as|11314,11316
needed|11317,11323
for|11324,11327
shortness|11328,11337
of|11338,11340
<EOL>|11341,11342
breath|11342,11348
or|11349,11351
wheezing|11352,11360
.|11360,11361
Disp|11362,11366
:|11366,11367
*|11367,11368
1|11368,11369
inhaler|11370,11377
*|11377,11378
Refills|11379,11386
:|11386,11387
*|11387,11388
1|11388,11389
*|11389,11390
<EOL>|11390,11391
<EOL>|11392,11393
Discharge|11393,11402
Disposition|11403,11414
:|11414,11415
<EOL>|11415,11416
Home|11416,11420
With|11421,11425
Service|11426,11433
<EOL>|11433,11434
<EOL>|11435,11436
Facility|11436,11444
:|11444,11445
<EOL>|11445,11446
_|11446,11447
_|11447,11448
_|11448,11449
<EOL>|11449,11450
<EOL>|11451,11452
Discharge|11452,11461
Diagnosis|11462,11471
:|11471,11472
<EOL>|11472,11473
-|11473,11474
Hypertension|11474,11486
with|11487,11491
hypertensive|11492,11504
urgency|11505,11512
<EOL>|11512,11513
-|11513,11514
Myocardial|11514,11524
infarction|11525,11535
attributed|11536,11546
to|11547,11549
demand|11550,11556
myonecrosis|11557,11568
<EOL>|11568,11569
-|11569,11570
Acute|11570,11575
on|11576,11578
chronic|11579,11586
left|11587,11591
ventricular|11592,11603
diastolic|11604,11613
heart|11614,11619
failure|11620,11627
<EOL>|11627,11628
-|11628,11629
Chronic|11629,11636
kidney|11637,11643
disease|11644,11651
,|11651,11652
stage|11653,11658
_|11659,11660
_|11660,11661
_|11661,11662
<EOL>|11662,11663
-|11663,11664
Chronic|11664,11671
obstructive|11672,11683
pulmonary|11684,11693
disease|11694,11701
<EOL>|11701,11702
-|11702,11703
Prior|11703,11708
cerebellar|11709,11719
-|11719,11720
medullary|11720,11729
stroke|11730,11736
<EOL>|11736,11737
-|11737,11738
Hyperlipidemia|11738,11752
<EOL>|11752,11753
-|11753,11754
Diabetes|11754,11762
mellitus|11763,11771
requiring|11772,11781
insulin|11782,11789
therapy|11790,11797
<EOL>|11797,11798
-|11798,11799
Medication|11799,11809
non-adherence|11810,11823
<EOL>|11823,11824
<EOL>|11825,11826
Mental|11847,11853
Status|11854,11860
:|11860,11861
Clear|11862,11867
and|11868,11871
coherent|11872,11880
.|11880,11881
<EOL>|11881,11882
Level|11882,11887
of|11888,11890
Consciousness|11891,11904
:|11904,11905
Alert|11906,11911
and|11912,11915
interactive|11916,11927
.|11927,11928
<EOL>|11928,11929
Activity|11929,11937
Status|11938,11944
:|11944,11945
Ambulatory|11946,11956
-|11957,11958
Independent|11959,11970
.|11970,11971
<EOL>|11971,11972
<EOL>|11973,11974
Dear|11998,12002
Ms.|12003,12006
_|12007,12008
_|12008,12009
_|12009,12010
,|12010,12011
<EOL>|12012,12013
<EOL>|12013,12014
You|12014,12017
were|12018,12022
admitted|12023,12031
for|12032,12035
shortness|12036,12045
of|12046,12048
breath|12049,12055
.|12055,12056
You|12057,12060
were|12061,12065
found|12066,12071
to|12072,12074
<EOL>|12075,12076
have|12076,12080
elevated|12081,12089
blood|12090,12095
pressure|12096,12104
on|12105,12107
admission|12108,12117
in|12118,12120
the|12121,12124
setting|12125,12132
of|12133,12135
not|12136,12139
<EOL>|12140,12141
taking|12141,12147
all|12148,12151
of|12152,12154
your|12155,12159
medications|12160,12171
regularly|12172,12181
.|12181,12182
We|12183,12185
obtained|12186,12194
an|12195,12197
<EOL>|12198,12199
echocargiogram|12199,12213
of|12214,12216
your|12217,12221
heart|12222,12227
which|12228,12233
showed|12234,12240
some|12241,12245
strain|12246,12252
on|12253,12255
your|12256,12260
<EOL>|12261,12262
heart|12262,12267
possibly|12268,12276
related|12277,12284
to|12285,12287
your|12288,12292
elevated|12293,12301
blood|12302,12307
pressures|12308,12317
.|12317,12318
<EOL>|12318,12319
<EOL>|12319,12320
You|12320,12323
will|12324,12328
be|12329,12331
contacted|12332,12341
about|12342,12347
an|12348,12350
outpatient|12351,12361
stress|12362,12368
test|12369,12373
.|12373,12374
This|12375,12379
will|12380,12384
<EOL>|12385,12386
be|12386,12388
completed|12389,12398
within|12399,12405
the|12406,12409
next|12410,12414
month|12415,12420
.|12420,12421
<EOL>|12421,12422
<EOL>|12422,12423
You|12423,12426
will|12427,12431
be|12432,12434
prescribed|12435,12445
several|12446,12453
new|12454,12457
medications|12458,12469
as|12470,12472
shown|12473,12478
below|12479,12484
.|12484,12485
A|12486,12487
<EOL>|12488,12489
visiting|12489,12497
nurse|12498,12503
_|12504,12505
_|12505,12506
_|12506,12507
come|12508,12512
to|12513,12515
your|12516,12520
home|12521,12525
to|12526,12528
help|12529,12533
with|12534,12538
managing|12539,12547
your|12548,12552
<EOL>|12553,12554
medications|12554,12565
.|12565,12566
You|12567,12570
should|12571,12577
dispose|12578,12585
of|12586,12588
all|12589,12592
your|12593,12597
home|12598,12602
medications|12603,12614
and|12615,12618
<EOL>|12619,12620
only|12620,12624
take|12625,12629
the|12630,12633
medications|12634,12645
shown|12646,12651
on|12652,12654
this|12655,12659
discharge|12660,12669
paperwork|12670,12679
.|12679,12680
<EOL>|12680,12681
<EOL>|12681,12682
STOP|12695,12699
Hydrochlorothiazide|12700,12719
<EOL>|12719,12720
STOP|12720,12724
Simvastatin|12725,12736
<EOL>|12736,12737
STOP|12737,12741
Clonidine|12742,12751
<EOL>|12751,12752
STOP|12752,12756
Atenolol|12757,12765
due|12766,12769
to|12770,12772
low|12773,12776
heart|12777,12782
rate|12783,12787
<EOL>|12787,12788
CHANGE|12788,12794
325mg|12795,12800
to|12801,12803
81mg|12804,12808
once|12809,12813
daily|12814,12819
<EOL>|12819,12820
START|12820,12825
Lisinopril|12826,12836
20mg|12837,12841
once|12842,12846
daily|12847,12852
<EOL>|12852,12853
START|12853,12858
Lasix|12859,12864
40mg|12865,12869
once|12870,12874
daily|12875,12880
<EOL>|12880,12881
START|12881,12886
Pravastin|12887,12896
80mg|12897,12901
once|12902,12906
daily|12907,12912
<EOL>|12912,12913
<EOL>|12913,12914
If|12914,12916
you|12917,12920
experience|12921,12931
any|12932,12935
chest|12936,12941
pain|12942,12946
,|12946,12947
excessive|12948,12957
shortness|12958,12967
of|12968,12970
breath|12971,12977
,|12977,12978
<EOL>|12979,12980
or|12980,12982
any|12983,12986
other|12987,12992
symptoms|12993,13001
concerning|13002,13012
to|13013,13015
you|13016,13019
,|13019,13020
please|13021,13027
call|13028,13032
or|13033,13035
come|13036,13040
<EOL>|13041,13042
into|13042,13046
the|13047,13050
emergency|13051,13060
department|13061,13071
for|13072,13075
further|13076,13083
evaluation|13084,13094
.|13094,13095
<EOL>|13095,13096
<EOL>|13096,13097
Thank|13097,13102
you|13103,13106
for|13107,13110
allowing|13111,13119
us|13120,13122
at|13123,13125
the|13126,13129
_|13130,13131
_|13131,13132
_|13132,13133
to|13134,13136
participate|13137,13148
in|13149,13151
your|13152,13156
care|13157,13161
.|13161,13162
<EOL>|13162,13163
<EOL>|13164,13165
Followup|13165,13173
Instructions|13174,13186
:|13186,13187
<EOL>|13187,13188
_|13188,13189
_|13189,13190
_|13190,13191
<EOL>|13191,13192

