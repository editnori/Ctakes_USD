 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
No|179,181
Known|182,187
Allergies|188,197
/|198,199
Adverse|200,207
Drug|208,212
Reactions|213,222
<EOL>|222,223
<EOL>|224,225
Attending|225,234
:|234,235
_|236,237
_|237,238
_|238,239
.|239,240
<EOL>|240,241
<EOL>|242,243
Chief|243,248
Complaint|249,258
:|258,259
<EOL>|259,260
Chest|260,265
pain|266,270
<EOL>|272,273
<EOL>|274,275
Major|275,280
Surgical|281,289
or|290,292
Invasive|293,301
Procedure|302,311
:|311,312
<EOL>|312,313
Cardiac|313,320
catheterization|321,336
with|337,341
stenting|342,350
with|351,355
drug|356,360
eluting|361,368
stent|369,374
to|375,377
<EOL>|378,379
the|379,382
left|383,387
circumflex|388,398
<EOL>|398,399
<EOL>|399,400
<EOL>|401,402
History|402,409
of|410,412
Present|413,420
Illness|421,428
:|428,429
<EOL>|429,430
_|430,431
_|431,432
_|432,433
year|434,438
old|439,442
woman|443,448
with|449,453
diastolic|454,463
CHF|464,467
,|467,468
COPD|469,473
,|473,474
DM|475,477
,|477,478
HTN|479,482
,|482,483
HLD|484,487
,|487,488
and|489,492
<EOL>|493,494
CAD|494,497
(|498,499
h|499,500
/|500,501
o|501,502
MI|503,505
in|506,508
_|509,510
_|510,511
_|511,512
with|513,517
LAD|518,521
stenting|522,530
,|530,531
repeat|532,538
stenting|539,547
with|548,552
DES|553,556
<EOL>|557,558
in|558,560
_|561,562
_|562,563
_|563,564
and|565,568
_|569,570
_|570,571
_|571,572
,|572,573
who|574,577
presents|578,586
with|587,591
chest|592,597
pain|598,602
.|602,603
She|604,607
has|608,611
been|612,616
<EOL>|617,618
having|618,624
chest|625,630
pain|631,635
episodes|636,644
over|645,649
the|650,653
past|654,658
2|659,660
weeks|661,666
.|666,667
A|668,669
tightness|670,679
<EOL>|680,681
located|681,688
in|689,691
the|692,695
_|696,697
_|697,698
_|698,699
her|700,703
chest|704,709
that|710,714
usually|715,722
occurs|723,729
with|730,734
<EOL>|735,736
exertion|736,744
or|745,747
when|748,752
lying|753,758
flat|759,763
at|764,766
night|767,772
,|772,773
but|774,777
she|778,781
has|782,785
also|786,790
<EOL>|791,792
experienced|792,803
at|804,806
rest|807,811
.|811,812
It|813,815
radiates|816,824
to|825,827
the|828,831
left|832,836
arm|837,840
,|840,841
and|842,845
is|846,848
<EOL>|849,850
relieved|850,858
with|859,863
NTG|864,867
.|867,868
It|869,871
is|872,874
not|875,878
pleuritic|879,888
,|888,889
but|890,893
is|894,896
reproducible|897,909
when|910,914
<EOL>|915,916
she|916,919
presses|920,927
over|928,932
the|933,936
_|937,938
_|938,939
_|939,940
her|941,944
chest|945,950
.|950,951
Somewhat|952,960
different|961,970
<EOL>|971,972
from|972,976
the|977,980
chest|981,986
pain|987,991
that|992,996
she|997,1000
had|1001,1004
prior|1005,1010
to|1011,1013
her|1014,1017
previous|1018,1026
PCIs|1027,1031
.|1031,1032
<EOL>|1033,1034
Associated|1034,1044
with|1045,1049
dsyspnea|1050,1058
and|1059,1062
lightheadedness|1063,1078
.|1078,1079
She|1080,1083
came|1084,1088
to|1089,1091
the|1092,1095
ED|1096,1098
<EOL>|1099,1100
today|1100,1105
after|1106,1111
having|1112,1118
a|1119,1120
more|1121,1125
severe|1126,1132
episode|1133,1140
yesterday|1141,1150
.|1150,1151
<EOL>|1153,1154
.|1154,1155
<EOL>|1157,1158
In|1158,1160
the|1161,1164
ED|1165,1167
initial|1168,1175
VS|1176,1178
were|1179,1183
:|1183,1184
97.5|1185,1189
,|1189,1190
67|1191,1193
,|1193,1194
127|1195,1198
/|1198,1199
73|1199,1201
,|1201,1202
16|1203,1205
,|1205,1206
100|1207,1210
%|1210,1211
RA|1211,1213
.|1213,1214
EKG|1215,1218
<EOL>|1219,1220
showed|1220,1226
SR|1227,1229
with|1230,1234
non-specific|1235,1247
ST|1248,1250
and|1251,1254
T|1255,1256
changes|1257,1264
.|1264,1265
CXR|1266,1269
negative|1270,1278
for|1279,1282
<EOL>|1283,1284
acute|1284,1289
process|1290,1297
.|1297,1298
Labs|1299,1303
notable|1304,1311
for|1312,1315
negative|1316,1324
troponin|1325,1333
but|1334,1337
Creat|1338,1343
1.7|1344,1347
<EOL>|1348,1349
(|1349,1350
was|1350,1353
1.4|1354,1357
in|1358,1360
_|1361,1362
_|1362,1363
_|1363,1364
and|1365,1368
normal|1369,1375
prior|1376,1381
to|1382,1384
that|1385,1389
)|1389,1390
.|1390,1391
She|1392,1395
received|1396,1404
ASA|1405,1408
<EOL>|1409,1410
325mg|1410,1415
.|1415,1416
VS|1417,1419
prior|1420,1425
to|1426,1428
transfer|1429,1437
were|1438,1442
:|1442,1443
97.6|1444,1448
,|1448,1449
70|1450,1452
,|1452,1453
119|1454,1457
/|1457,1458
60|1458,1460
,|1460,1461
16|1462,1464
,|1464,1465
99|1466,1468
%|1468,1469
RA|1469,1471
.|1471,1472
<EOL>|1474,1475
.|1475,1476
<EOL>|1478,1479
On|1479,1481
arrival|1482,1489
to|1490,1492
the|1493,1496
floor|1497,1502
,|1502,1503
patient|1504,1511
is|1512,1514
comfortable|1515,1526
and|1527,1530
denies|1531,1537
chest|1538,1543
<EOL>|1544,1545
pain|1545,1549
.|1549,1550
<EOL>|1552,1553
.|1553,1554
<EOL>|1556,1557
REVIEW|1557,1563
OF|1564,1566
SYSTEMS|1567,1574
:|1574,1575
As|1576,1578
noted|1579,1584
in|1585,1587
HPI|1588,1591
.|1591,1592
In|1593,1595
addition|1596,1604
,|1604,1605
denies|1606,1612
fevers|1613,1619
,|1619,1620
<EOL>|1621,1622
chills|1622,1628
,|1628,1629
sweats|1630,1636
,|1636,1637
presyncope|1638,1648
,|1648,1649
syncope|1650,1657
,|1657,1658
cough|1659,1664
,|1664,1665
PND|1666,1669
,|1669,1670
orthopnea|1671,1680
,|1680,1681
leg|1682,1685
<EOL>|1686,1687
swelling|1687,1695
,|1695,1696
abdominal|1697,1706
pain|1707,1711
,|1711,1712
nausea|1713,1719
,|1719,1720
vomiting|1721,1729
,|1729,1730
hematemesis|1731,1742
,|1742,1743
<EOL>|1744,1745
diarrhea|1745,1753
,|1753,1754
constipation|1755,1767
,|1767,1768
red|1769,1772
or|1773,1775
black|1776,1781
stools|1782,1788
,|1788,1789
dysuria|1790,1797
,|1797,1798
hematuria|1799,1808
,|1808,1809
<EOL>|1810,1811
myalgias|1811,1819
,|1819,1820
arthralgias|1821,1832
,|1832,1833
or|1834,1836
rash|1837,1841
.|1841,1842
No|1843,1845
history|1846,1853
of|1854,1856
DVT|1857,1860
or|1861,1863
PE|1864,1866
.|1866,1867
<EOL>|1869,1870
<EOL>|1870,1871
<EOL>|1872,1873
Past|1873,1877
Medical|1878,1885
History|1886,1893
:|1893,1894
<EOL>|1894,1895
-|1895,1896
CAD|1897,1900
:|1900,1901
MI|1902,1904
in|1905,1907
_|1908,1909
_|1909,1910
_|1910,1911
with|1912,1916
LAD|1917,1920
stenting|1921,1929
,|1929,1930
repeat|1931,1937
stenting|1938,1946
with|1947,1951
DES|1952,1955
in|1956,1958
<EOL>|1959,1960
<EOL>|1961,1962
_|1962,1963
_|1963,1964
_|1964,1965
and|1966,1969
_|1970,1971
_|1971,1972
_|1972,1973
<EOL>|1975,1976
-|1976,1977
Diastolic|1978,1987
CHF|1988,1991
<EOL>|1993,1994
-|1994,1995
DM|1996,1998
<EOL>|2000,2001
-|2001,2002
HTN|2003,2006
<EOL>|2008,2009
-|2009,2010
HLD|2011,2014
<EOL>|2016,2017
-|2017,2018
COPD|2019,2023
<EOL>|2025,2026
-|2026,2027
Depression|2028,2038
<EOL>|2040,2041
-|2041,2042
Right|2043,2048
shoulder|2049,2057
pain|2058,2062
(|2063,2064
bursitis|2064,2072
,|2072,2073
rotator|2074,2081
cuff|2082,2086
injury|2087,2093
)|2093,2094
<EOL>|2096,2097
<EOL>|2098,2099
Social|2099,2105
History|2106,2113
:|2113,2114
<EOL>|2114,2115
_|2115,2116
_|2116,2117
_|2117,2118
<EOL>|2118,2119
Family|2119,2125
History|2126,2133
:|2133,2134
<EOL>|2134,2135
She|2135,2138
was|2139,2142
a|2143,2144
ward|2145,2149
of|2150,2152
the|2153,2156
_|2157,2158
_|2158,2159
_|2159,2160
and|2161,2164
does|2165,2169
not|2170,2173
know|2174,2178
her|2179,2182
family|2183,2189
.|2189,2190
<EOL>|2192,2193
<EOL>|2193,2194
<EOL>|2195,2196
Physical|2196,2204
Exam|2205,2209
:|2209,2210
<EOL>|2210,2211
Admission|2211,2220
physical|2221,2229
exam|2230,2234
:|2234,2235
<EOL>|2235,2236
VS|2236,2238
:|2238,2239
98|2240,2242
,|2242,2243
139|2244,2247
/|2247,2248
76|2248,2250
,|2250,2251
71|2252,2254
,|2254,2255
18|2256,2258
,|2258,2259
100|2260,2263
%|2263,2264
RA|2265,2267
<EOL>|2269,2270
GENERAL|2270,2277
:|2277,2278
WDWN|2279,2283
woman|2284,2289
in|2290,2292
NAD|2293,2296
.|2296,2297
Oriented|2298,2306
x3|2307,2309
.|2309,2310
Mood|2311,2315
,|2315,2316
affect|2317,2323
<EOL>|2324,2325
appropriate|2325,2336
.|2336,2337
<EOL>|2339,2340
HEENT|2340,2345
:|2345,2346
NCAT|2347,2351
.|2351,2352
Sclera|2353,2359
anicteric|2360,2369
.|2369,2370
PERRL|2371,2376
,|2376,2377
EOMI|2378,2382
.|2382,2383
Conjunctiva|2384,2395
were|2396,2400
<EOL>|2401,2402
pink|2402,2406
,|2406,2407
no|2408,2410
pallor|2411,2417
or|2418,2420
cyanosis|2421,2429
of|2430,2432
the|2433,2436
oral|2437,2441
mucosa|2442,2448
.|2448,2449
No|2450,2452
xanthalesma|2453,2464
.|2464,2465
<EOL>|2467,2468
<EOL>|2468,2469
NECK|2469,2473
:|2473,2474
Supple|2475,2481
.|2481,2482
JVP|2483,2486
not|2487,2490
elevated|2491,2499
.|2499,2500
<EOL>|2502,2503
CARDIAC|2503,2510
:|2510,2511
RR|2512,2514
,|2514,2515
normal|2516,2522
S1|2523,2525
,|2525,2526
S2|2527,2529
.|2529,2530
No|2531,2533
m|2534,2535
/|2535,2536
r|2536,2537
/|2537,2538
g|2538,2539
.|2539,2540
No|2541,2543
S3|2544,2546
or|2547,2549
S4|2550,2552
.|2552,2553
Pain|2554,2558
<EOL>|2559,2560
reproducible|2560,2572
with|2573,2577
palpation|2578,2587
over|2588,2592
_|2593,2594
_|2594,2595
_|2595,2596
chest|2597,2602
and|2603,2606
left|2607,2611
<EOL>|2612,2613
breast|2613,2619
.|2619,2620
<EOL>|2622,2623
LUNGS|2623,2628
:|2628,2629
Resp|2630,2634
unlabored|2635,2644
,|2644,2645
no|2646,2648
accessory|2649,2658
muscle|2659,2665
use|2666,2669
.|2669,2670
CTAB|2671,2675
.|2675,2676
<EOL>|2678,2679
ABDOMEN|2679,2686
:|2686,2687
Soft|2688,2692
,|2692,2693
NTND|2694,2698
.|2698,2699
No|2700,2702
HSM|2703,2706
or|2707,2709
tenderness|2710,2720
.|2720,2721
Abd|2722,2725
aorta|2726,2731
not|2732,2735
<EOL>|2736,2737
enlarged|2737,2745
by|2746,2748
palpation|2749,2758
.|2758,2759
No|2760,2762
abdominial|2763,2773
bruits|2774,2780
.|2780,2781
<EOL>|2783,2784
EXTREMITIES|2784,2795
:|2795,2796
No|2797,2799
edema|2800,2805
.|2805,2806
WWP|2807,2810
.|2810,2811
<EOL>|2813,2814
SKIN|2814,2818
:|2818,2819
No|2820,2822
stasis|2823,2829
dermatitis|2830,2840
,|2840,2841
ulcers|2842,2848
,|2848,2849
scars|2850,2855
,|2855,2856
or|2857,2859
xanthomas|2860,2869
.|2869,2870
<EOL>|2872,2873
PULSES|2873,2879
:|2879,2880
<EOL>|2882,2883
Right|2883,2888
:|2888,2889
Carotid|2890,2897
2|2898,2899
+|2899,2900
Femoral|2901,2908
2|2909,2910
+|2910,2911
DP|2912,2914
2|2915,2916
+|2916,2917
_|2918,2919
_|2919,2920
_|2920,2921
2|2922,2923
+|2923,2924
<EOL>|2926,2927
Left|2927,2931
:|2931,2932
Carotid|2933,2940
2|2941,2942
+|2942,2943
Femoral|2944,2951
2|2952,2953
+|2953,2954
DP|2955,2957
2|2958,2959
+|2959,2960
_|2961,2962
_|2962,2963
_|2963,2964
2|2965,2966
+|2966,2967
<EOL>|2967,2968
.|2968,2969
<EOL>|2969,2970
Discharge|2970,2979
physical|2980,2988
exam|2989,2993
:|2993,2994
<EOL>|2995,2996
Vitals|2996,3002
:|3002,3003
Tc|3004,3006
98.1|3007,3011
BP|3012,3014
169|3015,3018
/|3018,3019
82|3019,3021
(|3022,3023
130|3023,3026
-|3026,3027
169|3027,3030
/|3030,3031
63|3031,3033
-|3033,3034
86|3034,3036
)|3036,3037
HR|3038,3040
71|3041,3043
(|3044,3045
70|3045,3047
-|3047,3048
77|3048,3050
)|3050,3051
RR|3052,3054
18|3055,3057
O2|3058,3060
<EOL>|3061,3062
Sat|3062,3065
98|3066,3068
%|3068,3069
RA|3070,3072
<EOL>|3073,3074
General|3074,3081
:|3081,3082
Patient|3083,3090
lying|3091,3096
in|3097,3099
bed|3100,3103
in|3104,3106
NAD|3107,3110
<EOL>|3110,3111
HEENT|3111,3116
:|3116,3117
EOMI|3118,3122
.|3122,3123
MMM|3124,3127
.|3127,3128
<EOL>|3128,3129
Neck|3129,3133
:|3133,3134
Supple|3135,3141
.|3141,3142
No|3143,3145
JVD|3146,3149
appreciated|3150,3161
.|3161,3162
<EOL>|3162,3163
CV|3163,3165
:|3165,3166
RRR|3167,3170
.|3170,3171
No|3172,3174
M|3175,3176
/|3176,3177
R|3177,3178
/|3178,3179
G|3179,3180
<EOL>|3180,3181
Lungs|3181,3186
:|3186,3187
Clear|3188,3193
to|3194,3196
auscultation|3197,3209
bilaterally|3210,3221
.|3221,3222
No|3223,3225
crackles|3226,3234
or|3235,3237
<EOL>|3238,3239
wheezes|3239,3246
.|3246,3247
Nml|3248,3251
work|3252,3256
of|3257,3259
breathing|3260,3269
.|3269,3270
<EOL>|3270,3271
Abd|3271,3274
:|3274,3275
Obese|3276,3281
.|3281,3282
NABS|3283,3287
+|3287,3288
.|3288,3289
Soft|3290,3294
.|3294,3295
NT|3296,3298
/|3298,3299
ND|3299,3301
.|3301,3302
<EOL>|3302,3303
Ext|3303,3306
:|3306,3307
WWP|3308,3311
.|3311,3312
2|3313,3314
+|3314,3315
DPs|3316,3319
bilaterally|3320,3331
.|3331,3332
No|3333,3335
clubbing|3336,3344
,|3344,3345
cyanosis|3346,3354
,|3354,3355
or|3356,3358
edema|3359,3364
.|3364,3365
<EOL>|3365,3366
<EOL>|3367,3368
Pertinent|3368,3377
Results|3378,3385
:|3385,3386
<EOL>|3386,3387
Admission|3387,3396
labs|3397,3401
:|3401,3402
<EOL>|3402,3403
_|3403,3404
_|3404,3405
_|3405,3406
10|3407,3409
:|3409,3410
10PM|3410,3414
BLOOD|3415,3420
WBC|3421,3424
-|3424,3425
10.9|3425,3429
RBC|3430,3433
-|3433,3434
3|3434,3435
.|3435,3436
78|3436,3438
*|3438,3439
Hgb|3440,3443
-|3443,3444
12.4|3444,3448
Hct|3449,3452
-|3452,3453
36.9|3453,3457
<EOL>|3458,3459
MCV|3459,3462
-|3462,3463
98|3463,3465
MCH|3466,3469
-|3469,3470
32|3470,3472
.|3472,3473
7|3473,3474
*|3474,3475
MCHC|3476,3480
-|3480,3481
33.6|3481,3485
RDW|3486,3489
-|3489,3490
12.5|3490,3494
Plt|3495,3498
_|3499,3500
_|3500,3501
_|3501,3502
<EOL>|3502,3503
_|3503,3504
_|3504,3505
_|3505,3506
10|3507,3509
:|3509,3510
10PM|3510,3514
BLOOD|3515,3520
Neuts|3521,3526
-|3526,3527
58.7|3527,3531
_|3532,3533
_|3533,3534
_|3534,3535
Monos|3536,3541
-|3541,3542
4.6|3542,3545
Eos|3546,3549
-|3549,3550
1.9|3550,3553
<EOL>|3554,3555
Baso|3555,3559
-|3559,3560
0.7|3560,3563
<EOL>|3563,3564
_|3564,3565
_|3565,3566
_|3566,3567
06|3568,3570
:|3570,3571
05AM|3571,3575
BLOOD|3576,3581
_|3582,3583
_|3583,3584
_|3584,3585
PTT|3586,3589
-|3589,3590
27.8|3590,3594
_|3595,3596
_|3596,3597
_|3597,3598
<EOL>|3598,3599
_|3599,3600
_|3600,3601
_|3601,3602
10|3603,3605
:|3605,3606
10PM|3606,3610
BLOOD|3611,3616
Glucose|3617,3624
-|3624,3625
338|3625,3628
*|3628,3629
UreaN|3630,3635
-|3635,3636
32|3636,3638
*|3638,3639
Creat|3640,3645
-|3645,3646
1|3646,3647
.|3647,3648
7|3648,3649
*|3649,3650
Na|3651,3653
-|3653,3654
134|3654,3657
<EOL>|3658,3659
K|3659,3660
-|3660,3661
4.3|3661,3664
Cl|3665,3667
-|3667,3668
100|3668,3671
HCO3|3672,3676
-|3676,3677
21|3677,3679
*|3679,3680
AnGap|3681,3686
-|3686,3687
17|3687,3689
<EOL>|3689,3690
_|3690,3691
_|3691,3692
_|3692,3693
10|3694,3696
:|3696,3697
10PM|3697,3701
BLOOD|3702,3707
cTropnT|3708,3715
-|3715,3716
<|3716,3717
0|3717,3718
.|3718,3719
01|3719,3721
<EOL>|3721,3722
<EOL>|3722,3723
Discharge|3723,3732
labs|3733,3737
:|3737,3738
<EOL>|3738,3739
_|3739,3740
_|3740,3741
_|3741,3742
06|3743,3745
:|3745,3746
05AM|3746,3750
BLOOD|3751,3756
WBC|3757,3760
-|3760,3761
10.1|3761,3765
RBC|3766,3769
-|3769,3770
3|3770,3771
.|3771,3772
74|3772,3774
*|3774,3775
Hgb|3776,3779
-|3779,3780
12.5|3780,3784
Hct|3785,3788
-|3788,3789
35|3789,3791
.|3791,3792
5|3792,3793
*|3793,3794
<EOL>|3795,3796
MCV|3796,3799
-|3799,3800
95|3800,3802
MCH|3803,3806
-|3806,3807
33|3807,3809
.|3809,3810
5|3810,3811
*|3811,3812
MCHC|3813,3817
-|3817,3818
35|3818,3820
.|3820,3821
2|3821,3822
*|3822,3823
RDW|3824,3827
-|3827,3828
12.8|3828,3832
Plt|3833,3836
_|3837,3838
_|3838,3839
_|3839,3840
<EOL>|3840,3841
_|3841,3842
_|3842,3843
_|3843,3844
06|3845,3847
:|3847,3848
05AM|3848,3852
BLOOD|3853,3858
Glucose|3859,3866
-|3866,3867
99|3867,3869
UreaN|3870,3875
-|3875,3876
29|3876,3878
*|3878,3879
Creat|3880,3885
-|3885,3886
1|3886,3887
.|3887,3888
4|3888,3889
*|3889,3890
Na|3891,3893
-|3893,3894
135|3894,3897
<EOL>|3898,3899
K|3899,3900
-|3900,3901
3.5|3901,3904
Cl|3905,3907
-|3907,3908
102|3908,3911
HCO3|3912,3916
-|3916,3917
26|3917,3919
AnGap|3920,3925
-|3925,3926
11|3926,3928
<EOL>|3928,3929
_|3929,3930
_|3930,3931
_|3931,3932
06|3933,3935
:|3935,3936
05AM|3936,3940
BLOOD|3941,3946
Calcium|3947,3954
-|3954,3955
9.0|3955,3958
Phos|3959,3963
-|3963,3964
4.3|3964,3967
Mg|3968,3970
-|3970,3971
2.0|3971,3974
<EOL>|3974,3975
<EOL>|3975,3976
Cardiac|3976,3983
enzymes|3984,3991
:|3991,3992
<EOL>|3992,3993
_|3993,3994
_|3994,3995
_|3995,3996
06|3997,3999
:|3999,4000
05AM|4000,4004
BLOOD|4005,4010
CK|4011,4013
(|4013,4014
CPK|4014,4017
)|4017,4018
-|4018,4019
61|4019,4021
<EOL>|4021,4022
_|4022,4023
_|4023,4024
_|4024,4025
06|4026,4028
:|4028,4029
05AM|4029,4033
BLOOD|4034,4039
CK|4040,4042
-|4042,4043
MB|4043,4045
-|4045,4046
2|4046,4047
cTropnT|4048,4055
-|4055,4056
<|4056,4057
0|4057,4058
.|4058,4059
01|4059,4061
<EOL>|4061,4062
_|4062,4063
_|4063,4064
_|4064,4065
10|4066,4068
:|4068,4069
10PM|4069,4073
BLOOD|4074,4079
cTropnT|4080,4087
-|4087,4088
<|4088,4089
0|4089,4090
.|4090,4091
01|4091,4093
<EOL>|4093,4094
<EOL>|4094,4095
EKG|4095,4098
:|4098,4099
<EOL>|4099,4100
Sinus|4100,4105
rhythm|4106,4112
at|4113,4115
a|4116,4117
rate|4118,4122
of|4123,4125
69|4126,4128
.|4128,4129
Normal|4130,4136
axis|4137,4141
.|4141,4142
The|4143,4146
PR|4147,4149
interval|4150,4158
is|4159,4161
<EOL>|4162,4163
prolonged|4163,4172
at|4173,4175
204ms|4176,4181
(|4182,4183
slightly|4183,4191
more|4192,4196
than|4197,4201
prior|4202,4207
ekg|4208,4211
)|4211,4212
.|4212,4213
Q|4214,4215
wave|4216,4220
in|4221,4223
<EOL>|4224,4225
III|4225,4228
.|4228,4229
Non-specific|4230,4242
ST|4243,4245
and|4246,4249
T|4250,4251
changes|4252,4259
.|4259,4260
<EOL>|4260,4261
<EOL>|4261,4262
Nuclear|4262,4269
Stress|4270,4276
Test|4277,4281
:|4281,4282
<EOL>|4283,4284
INTERPRETATION|4284,4298
:|4298,4299
<EOL>|4301,4302
The|4302,4305
image|4306,4311
quality|4312,4319
is|4320,4322
adequate|4323,4331
but|4332,4335
limited|4336,4343
due|4344,4347
to|4348,4350
soft|4351,4355
tissue|4356,4362
and|4363,4366
<EOL>|4367,4368
breast|4368,4374
attenuation|4375,4386
.|4386,4387
There|4388,4393
is|4394,4396
activity|4397,4405
adjacent|4406,4414
to|4415,4417
the|4418,4421
heart|4422,4427
in|4428,4430
<EOL>|4431,4432
the|4432,4435
rest|4436,4440
and|4441,4444
stress|4445,4451
images|4452,4458
.|4458,4459
<EOL>|4460,4461
Left|4461,4465
ventricular|4466,4477
cavity|4478,4484
size|4485,4489
is|4490,4492
increased|4493,4502
.|4502,4503
<EOL>|4504,4505
Rest|4505,4509
and|4510,4513
stress|4514,4520
perfusion|4521,4530
images|4531,4537
reveal|4538,4544
a|4545,4546
reversible|4547,4557
,|4557,4558
moderate|4559,4567
<EOL>|4568,4569
reduction|4569,4578
in|4579,4581
photon|4582,4588
counts|4589,4595
involving|4596,4605
the|4606,4609
mid|4610,4613
and|4614,4617
basal|4618,4623
<EOL>|4624,4625
inferolateral|4625,4638
walls|4639,4644
and|4645,4648
the|4649,4652
distal|4653,4659
lateral|4660,4667
wall|4668,4672
.|4672,4673
Gated|4674,4679
images|4680,4686
<EOL>|4687,4688
reveal|4688,4694
normal|4695,4701
wall|4702,4706
motion|4707,4713
.|4713,4714
<EOL>|4716,4717
The|4717,4720
calculated|4721,4731
left|4732,4736
ventricular|4737,4748
ejection|4749,4757
fraction|4758,4766
is|4767,4769
52|4770,4772
%|4772,4773
with|4774,4778
an|4779,4781
<EOL>|4782,4783
EDV|4783,4786
of|4787,4789
107|4790,4793
ml|4794,4796
(|4797,4798
reprocessed|4798,4809
at|4810,4812
workstation|4813,4824
)|4824,4825
.|4825,4826
<EOL>|4828,4829
IMPRESSION|4829,4839
:|4839,4840
<EOL>|4841,4842
1.|4842,4844
Reversible|4845,4855
,|4855,4856
medium|4857,4863
sized|4864,4869
,|4869,4870
moderate|4871,4879
severity|4880,4888
perfusion|4889,4898
defect|4899,4905
<EOL>|4906,4907
involving|4907,4916
the|4917,4920
LCx|4921,4924
territory|4925,4934
.|4934,4935
<EOL>|4936,4937
2.|4937,4939
Increased|4940,4949
left|4950,4954
ventricular|4955,4966
cavity|4967,4973
size|4974,4978
with|4979,4983
normal|4984,4990
systolic|4991,4999
<EOL>|5000,5001
function|5001,5009
.|5009,5010
<EOL>|5011,5012
Compared|5012,5020
to|5021,5023
the|5024,5027
prior|5028,5033
study|5034,5039
of|5040,5042
_|5043,5044
_|5044,5045
_|5045,5046
,|5046,5047
the|5048,5051
defect|5052,5058
is|5059,5061
new|5062,5065
.|5065,5066
<EOL>|5067,5068
.|5068,5069
<EOL>|5069,5070
Cardiac|5070,5077
catheterization|5078,5093
:|5093,5094
<EOL>|5094,5095
COMMENTS|5095,5103
:|5103,5104
<EOL>|5110,5111
1.|5111,5113
Selective|5114,5123
coronary|5124,5132
angiography|5133,5144
of|5145,5147
this|5148,5152
right|5153,5158
-|5158,5159
dominant|5159,5167
system|5168,5174
<EOL>|5175,5176
demonstrated|5176,5188
three|5189,5194
-|5194,5195
vessel|5195,5201
coronary|5202,5210
artery|5211,5217
disease|5218,5225
.|5225,5226
The|5228,5231
_|5232,5233
_|5233,5234
_|5234,5235
did|5236,5239
<EOL>|5240,5241
not|5241,5244
<EOL>|5245,5246
have|5246,5250
angiographically|5251,5267
-|5267,5268
apparent|5268,5276
flow|5277,5281
-|5281,5282
limiting|5282,5290
stenoses|5291,5299
.|5299,5300
The|5302,5305
LAD|5306,5309
<EOL>|5310,5311
had|5311,5314
60|5315,5317
%|5317,5318
<EOL>|5319,5320
in|5320,5322
-|5322,5323
stent|5323,5328
restenosis|5329,5339
at|5340,5342
the|5343,5346
junction|5347,5355
of|5356,5358
the|5359,5362
old|5363,5366
Cypher|5367,5373
stent|5374,5379
<EOL>|5380,5381
placed|5381,5387
in|5388,5390
<EOL>|5391,5392
_|5392,5393
_|5393,5394
_|5394,5395
and|5396,5399
the|5400,5403
new|5404,5407
Promus|5408,5414
stent|5415,5420
placed|5421,5427
in|5428,5430
_|5431,5432
_|5432,5433
_|5433,5434
the|5435,5438
D2|5439,5441
branch|5442,5448
was|5449,5452
<EOL>|5453,5454
jailed|5454,5460
<EOL>|5461,5462
with|5462,5466
60|5467,5469
%|5469,5470
origin|5471,5477
stenosis|5478,5486
.|5486,5487
The|5489,5492
LCx|5493,5496
had|5497,5500
a|5501,5502
50|5503,5505
%|5505,5506
stenosis|5507,5515
at|5516,5518
its|5519,5522
<EOL>|5523,5524
origin|5524,5530
;|5530,5531
<EOL>|5532,5533
there|5533,5538
was|5539,5542
a|5543,5544
90|5545,5547
%|5547,5548
stenosis|5549,5557
of|5558,5560
the|5561,5564
OM1|5565,5568
branch|5569,5575
.|5575,5576
The|5578,5581
mid-RCA|5582,5589
had|5590,5593
a|5594,5595
<EOL>|5596,5597
50|5597,5599
%|5599,5600
<EOL>|5601,5602
stenosis|5602,5610
.|5610,5611
<EOL>|5612,5613
2.|5613,5615
Limited|5616,5623
resting|5624,5631
hemodynamics|5632,5644
revealed|5645,5653
mild|5654,5658
systemic|5659,5667
arterial|5668,5676
<EOL>|5677,5678
hypertension|5678,5690
,|5690,5691
with|5692,5696
a|5697,5698
central|5699,5706
aortic|5707,5713
pressure|5714,5722
of|5723,5725
142|5726,5729
/|5729,5730
74|5730,5732
mmHg|5733,5737
.|5737,5738
<EOL>|5739,5740
3.|5740,5742
Successful|5743,5753
PTCA|5754,5758
and|5759,5762
stenting|5763,5771
of|5772,5774
OM1|5775,5778
with|5779,5783
a|5784,5785
3.0|5786,5789
x15mm|5789,5794
PROMUS|5795,5801
<EOL>|5802,5803
stent|5803,5808
<EOL>|5809,5810
which|5810,5815
was|5816,5819
postdilated|5820,5831
to|5832,5834
3.5|5835,5838
mm|5838,5840
.|5840,5841
Final|5842,5847
angiography|5848,5859
revealed|5860,5868
no|5869,5871
<EOL>|5872,5873
residual|5873,5881
<EOL>|5882,5883
stenosis|5883,5891
,|5891,5892
no|5893,5895
angiographically|5896,5912
apparent|5913,5921
dissection|5922,5932
and|5933,5936
TIMI|5937,5941
III|5942,5945
<EOL>|5946,5947
flow|5947,5951
(|5952,5953
see|5953,5956
<EOL>|5957,5958
PTCA|5958,5962
comments|5963,5971
)|5971,5972
.|5972,5973
<EOL>|5974,5975
FINAL|5975,5980
DIAGNOSIS|5981,5990
:|5990,5991
<EOL>|5996,5997
1.|5997,5999
Three|6000,6005
vessel|6006,6012
coronary|6013,6021
artery|6022,6028
disease|6029,6036
.|6036,6037
<EOL>|6038,6039
2.|6039,6041
Successful|6042,6052
PTCA|6053,6057
and|6058,6061
stenting|6062,6070
of|6071,6073
the|6074,6077
OM1|6078,6081
with|6082,6086
a|6087,6088
DES|6089,6092
.|6092,6093
<EOL>|6094,6095
.|6095,6096
<EOL>|6096,6097
<EOL>|6097,6098
<EOL>|6099,6100
Brief|6100,6105
Hospital|6106,6114
Course|6115,6121
:|6121,6122
<EOL>|6122,6123
#|6123,6124
Unstable|6125,6133
angina|6134,6140
:|6140,6141
Description|6142,6153
of|6154,6156
the|6157,6160
pain|6161,6165
was|6166,6169
somewhat|6170,6178
atypical|6179,6187
<EOL>|6188,6189
for|6189,6192
angina|6193,6199
in|6200,6202
that|6203,6207
she|6208,6211
experiences|6212,6223
in|6224,6226
when|6227,6231
she|6232,6235
lays|6236,6240
down|6241,6245
and|6246,6249
it|6250,6252
<EOL>|6253,6254
is|6254,6256
also|6257,6261
reproducible|6262,6274
.|6274,6275
However|6276,6283
,|6283,6284
given|6285,6290
her|6291,6294
history|6295,6302
of|6303,6305
CAD|6306,6309
status|6310,6316
<EOL>|6317,6318
post|6318,6322
multiple|6323,6331
PCIs|6332,6336
and|6337,6340
many|6341,6345
risk|6346,6350
factors|6351,6358
,|6358,6359
the|6360,6363
patient|6364,6371
underwent|6372,6381
<EOL>|6382,6383
stress|6383,6389
test|6390,6394
to|6395,6397
rule|6398,6402
out|6403,6406
CAD|6407,6410
.|6410,6411
Nuclear|6412,6419
stress|6420,6426
test|6427,6431
showed|6432,6438
a|6439,6440
<EOL>|6441,6442
reversible|6442,6452
,|6452,6453
medium|6454,6460
sized|6461,6466
,|6466,6467
moderate|6468,6476
severity|6477,6485
perfusion|6486,6495
defect|6496,6502
<EOL>|6503,6504
involving|6504,6513
the|6514,6517
left|6518,6522
circumflex|6523,6533
territory|6534,6543
.|6543,6544
In|6545,6547
light|6548,6553
of|6554,6556
these|6557,6562
<EOL>|6563,6564
stress|6564,6570
test|6571,6575
findings|6576,6584
,|6584,6585
the|6586,6589
patient|6590,6597
underwent|6598,6607
cardiac|6608,6615
<EOL>|6616,6617
catheterization|6617,6632
.|6632,6633
Prior|6634,6639
to|6640,6642
cardiac|6643,6650
catheterization|6651,6666
,|6666,6667
she|6668,6671
was|6672,6675
<EOL>|6676,6677
prehydrated|6677,6688
given|6689,6694
her|6695,6698
acute|6699,6704
kidney|6705,6711
injury|6712,6718
.|6718,6719
The|6720,6723
patient|6724,6731
had|6732,6735
a|6736,6737
<EOL>|6738,6739
drug|6739,6743
-|6743,6744
eluting|6744,6751
stent|6752,6757
placed|6758,6764
to|6765,6767
the|6768,6771
obtuse|6772,6778
marginal|6779,6787
branch|6788,6794
.|6794,6795
The|6796,6799
<EOL>|6800,6801
patient|6801,6808
became|6809,6815
acutely|6816,6823
hypertensive|6824,6836
during|6837,6843
cardiac|6844,6851
<EOL>|6852,6853
catheterization|6853,6868
and|6869,6872
was|6873,6876
started|6877,6884
on|6885,6887
a|6888,6889
nitroglycerin|6890,6903
drip|6904,6908
(|6909,6910
see|6910,6913
<EOL>|6914,6915
discussion|6915,6925
below|6926,6931
)|6931,6932
.|6932,6933
The|6934,6937
patient|6938,6945
was|6946,6949
weaned|6950,6956
from|6957,6961
this|6962,6966
quickly|6967,6974
.|6974,6975
The|6976,6979
<EOL>|6980,6981
patient|6981,6988
was|6989,6992
continued|6993,7002
on|7003,7005
aspirin|7006,7013
(|7014,7015
full|7015,7019
-|7019,7020
dose|7020,7024
)|7024,7025
,|7025,7026
plavix|7027,7033
,|7033,7034
<EOL>|7035,7036
metoprolol|7036,7046
,|7046,7047
and|7048,7051
imdur|7052,7057
.|7057,7058
Her|7059,7062
home|7063,7067
dose|7068,7072
of|7073,7075
atorvastatin|7076,7088
was|7089,7092
<EOL>|7093,7094
increased|7094,7103
given|7104,7109
evidence|7110,7118
of|7119,7121
coronary|7122,7130
artery|7131,7137
disease|7138,7145
.|7145,7146
Serial|7147,7153
<EOL>|7154,7155
cardiac|7155,7162
enzymes|7163,7170
were|7171,7175
negative|7176,7184
times|7185,7190
3|7191,7192
.|7192,7193
<EOL>|7193,7194
OUTPATIENT|7197,7207
ISSUES|7208,7214
:|7214,7215
Patient|7216,7223
is|7224,7226
to|7227,7229
continue|7230,7238
taking|7239,7245
aspirin|7246,7253
<EOL>|7254,7255
325mg|7255,7260
and|7261,7264
plavix|7265,7271
75mg|7272,7276
daily|7277,7282
for|7283,7286
the|7287,7290
next|7291,7295
year|7296,7300
.|7300,7301
Patient|7302,7309
will|7310,7314
have|7315,7319
<EOL>|7320,7321
cardiology|7321,7331
follow|7332,7338
-|7338,7339
up|7339,7341
as|7342,7344
an|7345,7347
outpatient|7348,7358
with|7359,7363
the|7364,7367
_|7368,7369
_|7369,7370
_|7370,7371
<EOL>|7372,7373
_|7373,7374
_|7374,7375
_|7375,7376
_|7377,7378
_|7378,7379
_|7379,7380
group|7381,7386
in|7387,7389
_|7390,7391
_|7391,7392
_|7392,7393
.|7393,7394
<EOL>|7395,7396
.|7396,7397
<EOL>|7399,7400
#|7400,7401
Acute|7402,7407
kidney|7408,7414
injury|7415,7421
:|7421,7422
Creatinine|7423,7433
currently|7434,7443
1.7|7444,7447
,|7447,7448
up|7449,7451
from|7452,7456
1.4|7457,7460
in|7461,7463
<EOL>|7464,7465
_|7465,7466
_|7466,7467
_|7467,7468
.|7468,7469
Renal|7470,7475
function|7476,7484
previously|7485,7495
was|7496,7499
normal|7500,7506
.|7506,7507
Upon|7508,7512
admission|7513,7522
,|7522,7523
<EOL>|7524,7525
the|7525,7528
patient|7529,7536
's|7536,7538
lisinopril|7539,7549
and|7550,7553
furosemide|7554,7564
were|7565,7569
discontinued|7570,7582
.|7582,7583
Of|7584,7586
<EOL>|7587,7588
note|7588,7592
,|7592,7593
hte|7594,7597
patient|7598,7605
was|7606,7609
started|7610,7617
on|7618,7620
furosemide|7621,7631
approximately|7632,7645
_|7646,7647
_|7647,7648
_|7648,7649
<EOL>|7650,7651
months|7651,7657
ago|7658,7661
,|7661,7662
which|7663,7668
coincides|7669,7678
with|7679,7683
the|7684,7687
development|7688,7699
of|7700,7702
the|7703,7706
<EOL>|7707,7708
patient|7708,7715
's|7715,7717
elevated|7718,7726
serum|7727,7732
creatinine|7733,7743
.|7743,7744
Serum|7745,7750
creatinine|7751,7761
was|7762,7765
<EOL>|7766,7767
trended|7767,7774
through|7775,7782
the|7783,7786
admission|7787,7796
and|7797,7800
improved|7801,7809
.|7809,7810
The|7811,7814
patient|7815,7822
was|7823,7826
<EOL>|7827,7828
restarted|7828,7837
on|7838,7840
her|7841,7844
home|7845,7849
lisinopril|7850,7860
,|7860,7861
though|7862,7868
her|7869,7872
serum|7873,7878
creatinine|7879,7889
<EOL>|7890,7891
was|7891,7894
noticed|7895,7902
to|7903,7905
be|7906,7908
increasing|7909,7919
so|7920,7922
was|7923,7926
discontinued|7927,7939
with|7940,7944
<EOL>|7945,7946
instructions|7946,7958
to|7959,7961
restart|7962,7969
this|7970,7974
medication|7975,7985
after|7986,7991
follow|7992,7998
-|7998,7999
up|7999,8001
with|8002,8006
her|8007,8010
<EOL>|8011,8012
primary|8012,8019
care|8020,8024
physician|8025,8034
.|8034,8035
The|8036,8039
patient|8040,8047
was|8048,8051
instructed|8052,8062
to|8063,8065
have|8066,8070
a|8071,8072
<EOL>|8073,8074
basic|8074,8079
metabolic|8080,8089
panel|8090,8095
drawn|8096,8101
_|8102,8103
_|8103,8104
_|8104,8105
.|8105,8106
<EOL>|8107,8108
.|8108,8109
<EOL>|8111,8112
#|8112,8113
Diastolic|8114,8123
heart|8124,8129
failure|8130,8137
:|8137,8138
Patient|8139,8146
was|8147,8150
euvolemic|8151,8160
through|8161,8168
her|8169,8172
<EOL>|8173,8174
admission|8174,8183
.|8183,8184
Her|8185,8188
home|8189,8193
lasix|8194,8199
was|8200,8203
discontinued|8204,8216
during|8217,8223
this|8224,8228
admission|8229,8238
<EOL>|8239,8240
given|8240,8245
her|8246,8249
acute|8250,8255
kidney|8256,8262
injury|8263,8269
.|8269,8270
The|8271,8274
patient|8275,8282
will|8283,8287
follow|8288,8294
-|8294,8295
up|8295,8297
with|8298,8302
<EOL>|8303,8304
her|8304,8307
primary|8308,8315
care|8316,8320
physician|8321,8330
regarding|8331,8340
_|8341,8342
_|8342,8343
_|8343,8344
of|8345,8347
lasix|8348,8353
.|8353,8354
<EOL>|8355,8356
OUTPATIENT|8359,8369
ISSUES|8370,8376
:|8376,8377
Outpatient|8378,8388
BMP|8389,8392
for|8393,8396
monitoring|8397,8407
of|8408,8410
serum|8411,8416
<EOL>|8417,8418
creatinine|8418,8428
and|8429,8432
reinitiation|8433,8445
of|8446,8448
lasix|8449,8454
by|8455,8457
the|8458,8461
primary|8462,8469
care|8470,8474
<EOL>|8475,8476
physician|8476,8485
.|8485,8486
<EOL>|8487,8488
.|8488,8489
<EOL>|8491,8492
#|8492,8493
Type|8494,8498
2|8499,8500
Diabetes|8501,8509
Melltius|8510,8518
,|8518,8519
insulin|8520,8527
dependent|8528,8537
:|8537,8538
Moderately|8539,8549
<EOL>|8550,8551
controlled|8551,8561
with|8562,8566
last|8567,8571
A1c|8572,8575
7.9|8576,8579
%|8579,8580
in|8581,8583
_|8584,8585
_|8585,8586
_|8586,8587
.|8587,8588
Lantus|8589,8595
and|8596,8599
sliding|8600,8607
<EOL>|8608,8609
scale|8609,8614
was|8615,8618
continued|8619,8628
through|8629,8636
the|8637,8640
hospitalization|8641,8656
.|8656,8657
She|8658,8661
was|8662,8665
<EOL>|8666,8667
discharged|8667,8677
home|8678,8682
on|8683,8685
her|8686,8689
home|8690,8694
doses|8695,8700
of|8701,8703
lantus|8704,8710
and|8711,8714
her|8715,8718
home|8719,8723
insulin|8724,8731
<EOL>|8732,8733
sliding|8733,8740
scale|8741,8746
.|8746,8747
<EOL>|8750,8751
.|8751,8752
<EOL>|8752,8753
#|8753,8754
Hypertension|8755,8767
:|8767,8768
Through|8769,8776
most|8777,8781
of|8782,8784
the|8785,8788
patient|8789,8796
's|8796,8798
admission|8799,8808
,|8808,8809
her|8810,8813
<EOL>|8814,8815
blood|8815,8820
pressure|8821,8829
was|8830,8833
well|8835,8839
controlled|8840,8850
(|8851,8852
goal|8852,8856
<|8857,8858
130|8858,8861
/|8861,8862
80|8862,8864
)|8864,8865
.|8865,8866
She|8867,8870
was|8871,8874
<EOL>|8875,8876
continued|8876,8885
on|8886,8888
metoprolol|8889,8899
and|8900,8903
imdur|8904,8909
,|8909,8910
though|8911,8917
furosemide|8918,8928
and|8929,8932
<EOL>|8933,8934
lisinopril|8934,8944
were|8945,8949
discontinued|8950,8962
in|8963,8965
light|8966,8971
of|8972,8974
the|8975,8978
patient|8979,8986
's|8986,8988
elevated|8989,8997
<EOL>|8998,8999
serum|8999,9004
creatinine|9005,9015
.|9015,9016
However|9017,9024
,|9024,9025
during|9026,9032
the|9033,9036
patient|9037,9044
's|9044,9046
cardiac|9047,9054
<EOL>|9055,9056
catheterization|9056,9071
,|9071,9072
she|9073,9076
was|9077,9080
noted|9081,9086
to|9087,9089
have|9090,9094
elevated|9095,9103
systolic|9104,9112
blood|9113,9118
<EOL>|9119,9120
pressures|9120,9129
and|9130,9133
was|9134,9137
started|9138,9145
on|9146,9148
a|9149,9150
nitroglycerin|9151,9164
drip|9165,9169
for|9170,9173
control|9174,9181
of|9182,9184
<EOL>|9185,9186
blood|9186,9191
pressures|9192,9201
.|9201,9202
The|9203,9206
patient|9207,9214
was|9215,9218
weaned|9219,9225
from|9226,9230
the|9231,9234
nitroglycerin|9235,9248
<EOL>|9249,9250
drip|9250,9254
with|9255,9259
in|9260,9262
4|9263,9264
hours|9265,9270
after|9271,9276
cardiac|9277,9284
catheterization|9285,9300
.|9300,9301
The|9302,9305
patient|9306,9313
<EOL>|9314,9315
received|9315,9323
a|9324,9325
dose|9326,9330
of|9331,9333
lisinopril|9334,9344
,|9344,9345
but|9346,9349
because|9350,9357
of|9358,9360
rising|9361,9367
serum|9368,9373
<EOL>|9374,9375
creatinine|9375,9385
,|9385,9386
the|9387,9390
patient|9391,9398
's|9398,9400
next|9401,9405
dose|9406,9410
was|9411,9414
held|9415,9419
.|9419,9420
<EOL>|9421,9422
OUTPATIENT|9425,9435
ISSUES|9436,9442
:|9442,9443
Follow|9444,9450
-|9450,9451
up|9451,9453
with|9454,9458
primary|9459,9466
care|9467,9471
physician|9472,9481
<EOL>|9482,9483
regarding|9483,9492
recent|9493,9499
hospitalization|9500,9515
and|9516,9519
anti-hypertensive|9520,9537
regimen|9538,9545
<EOL>|9546,9547
in|9547,9549
light|9550,9555
of|9556,9558
elevated|9559,9567
serum|9568,9573
creatinine|9574,9584
.|9584,9585
<EOL>|9587,9588
.|9588,9589
<EOL>|9589,9590
#|9590,9591
Hyperlipidemia|9592,9606
:|9606,9607
Well|9608,9612
controlled|9613,9623
with|9624,9628
last|9629,9633
LDL|9634,9637
50|9638,9640
in|9641,9643
_|9644,9645
_|9645,9646
_|9646,9647
<EOL>|9648,9649
(|9649,9650
goal|9650,9654
LDL|9655,9658
<|9658,9659
70|9659,9661
)|9661,9662
,|9662,9663
though|9664,9670
triglycerides|9671,9684
mildly|9685,9691
elevated|9692,9700
.|9700,9701
<EOL>|9703,9704
Atorvastatin|9704,9716
was|9717,9720
increased|9721,9730
to|9731,9733
80mg|9734,9738
daily|9739,9744
given|9745,9750
the|9751,9754
new|9755,9758
CAD|9759,9762
<EOL>|9763,9764
lesions|9764,9771
.|9771,9772
Patient|9773,9780
also|9781,9785
had|9786,9789
a|9790,9791
fasting|9792,9799
lipid|9800,9805
panel|9806,9811
that|9812,9816
was|9817,9820
drawn|9821,9826
,|9826,9827
<EOL>|9828,9829
which|9829,9834
was|9835,9838
pending|9839,9846
at|9847,9849
time|9850,9854
of|9855,9857
discharge|9858,9867
.|9867,9868
<EOL>|9868,9869
OUTPATIENT|9872,9882
ISSUES|9883,9889
:|9889,9890
Follow|9891,9897
-|9897,9898
up|9898,9900
of|9901,9903
pending|9904,9911
fasting|9912,9919
lipid|9920,9925
panel|9926,9931
.|9931,9932
<EOL>|9934,9935
<EOL>|9935,9936
.|9936,9937
<EOL>|9938,9939
#|9939,9940
COPD|9941,9945
:|9945,9946
Currently|9947,9956
asymptomatic|9957,9969
.|9969,9970
Patient|9971,9978
was|9979,9982
continue|9983,9991
fluticasone|9992,10003
<EOL>|10004,10005
and|10005,10008
albuterol|10009,10018
as|10019,10021
needed|10022,10028
.|10028,10029
<EOL>|10032,10033
<EOL>|10033,10034
<EOL>|10035,10036
Medications|10036,10047
on|10048,10050
Admission|10051,10060
:|10060,10061
<EOL>|10061,10062
-|10062,10063
Clopidogrel|10064,10075
75|10076,10078
mg|10079,10081
daily|10082,10087
<EOL>|10089,10090
-|10090,10091
Asprin|10092,10098
325|10099,10102
mg|10103,10105
daily|10106,10111
<EOL>|10113,10114
-|10114,10115
Atorvastatin|10116,10128
40|10129,10131
mg|10132,10134
daily|10135,10140
<EOL>|10142,10143
-|10143,10144
Lisinopril|10145,10155
10|10156,10158
mg|10159,10161
daily|10162,10167
<EOL>|10169,10170
-|10170,10171
Metoprolol|10172,10182
succinate|10183,10192
100|10193,10196
mg|10197,10199
daily|10200,10205
<EOL>|10207,10208
-|10208,10209
Isosorbide|10210,10220
mononitrate|10221,10232
30|10233,10235
mg|10236,10238
daily|10239,10244
<EOL>|10246,10247
-|10247,10248
Furosemide|10249,10259
20|10260,10262
mg|10263,10265
daily|10266,10271
<EOL>|10273,10274
-|10274,10275
Nitroglycerin|10276,10289
0.4|10290,10293
mg|10294,10296
SL|10297,10299
prn|10300,10303
<EOL>|10305,10306
-|10306,10307
Glargine|10308,10316
insulin|10317,10324
80|10325,10327
units|10328,10333
QHS|10334,10337
<EOL>|10339,10340
-|10340,10341
Lispro|10342,10348
insulin|10349,10356
sliding|10357,10364
scale|10365,10370
<EOL>|10372,10373
-|10373,10374
Albuterol|10375,10384
90|10385,10387
mcg|10388,10391
,|10391,10392
2|10393,10394
puffs|10395,10400
Q4|10401,10403
-|10403,10404
6|10404,10405
hrs|10406,10409
prn|10410,10413
<EOL>|10415,10416
-|10416,10417
Fluticasone|10418,10429
110|10430,10433
mcg|10434,10437
,|10437,10438
2|10439,10440
puffs|10441,10446
BID|10447,10450
<EOL>|10452,10453
-|10453,10454
Pantoprazole|10455,10467
40|10468,10470
mg|10471,10473
BID|10474,10477
<EOL>|10479,10480
-|10480,10481
Oxycode|10482,10489
-|10489,10490
Acetaminophen|10490,10503
5|10504,10505
mg|10506,10508
-|10508,10509
325|10509,10512
mg|10513,10515
Q8h|10516,10519
prn|10520,10523
pain|10524,10528
<EOL>|10530,10531
-|10531,10532
Potassium|10533,10542
chloride|10543,10551
20|10552,10554
mEq|10555,10558
BID|10559,10562
<EOL>|10564,10565
-|10565,10566
Cholecalciferol|10567,10582
1,000|10583,10588
unit|10589,10593
daily|10594,10599
<EOL>|10601,10602
-|10602,10603
Metronidazole|10604,10617
0.75|10618,10622
%|10622,10623
lotion|10624,10630
for|10631,10634
_|10635,10636
_|10636,10637
_|10637,10638
<EOL>|10640,10641
<EOL>|10641,10642
<EOL>|10643,10644
Discharge|10644,10653
Medications|10654,10665
:|10665,10666
<EOL>|10666,10667
1.|10667,10669
clopidogrel|10670,10681
75|10682,10684
mg|10685,10687
Tablet|10688,10694
Sig|10695,10698
:|10698,10699
One|10700,10703
(|10704,10705
1|10705,10706
)|10706,10707
Tablet|10708,10714
PO|10715,10717
DAILY|10718,10723
<EOL>|10724,10725
(|10725,10726
Daily|10726,10731
)|10731,10732
.|10732,10733
<EOL>|10735,10736
2.|10736,10738
aspirin|10739,10746
325|10747,10750
mg|10751,10753
Tablet|10754,10760
Sig|10761,10764
:|10764,10765
One|10766,10769
(|10770,10771
1|10771,10772
)|10772,10773
Tablet|10774,10780
PO|10781,10783
DAILY|10784,10789
(|10790,10791
Daily|10791,10796
)|10796,10797
.|10797,10798
<EOL>|10800,10801
3.|10801,10803
atorvastatin|10804,10816
40|10817,10819
mg|10820,10822
Tablet|10823,10829
Sig|10830,10833
:|10833,10834
One|10835,10838
(|10839,10840
1|10840,10841
)|10841,10842
Tablet|10843,10849
PO|10850,10852
DAILY|10853,10858
<EOL>|10859,10860
(|10860,10861
Daily|10861,10866
)|10866,10867
.|10867,10868
<EOL>|10870,10871
4.|10871,10873
metoprolol|10874,10884
succinate|10885,10894
100|10895,10898
mg|10899,10901
Tablet|10902,10908
Extended|10909,10917
Release|10918,10925
24|10926,10928
hr|10929,10931
<EOL>|10932,10933
Sig|10933,10936
:|10936,10937
One|10938,10941
(|10942,10943
1|10943,10944
)|10944,10945
Tablet|10946,10952
Extended|10953,10961
Release|10962,10969
24|10970,10972
hr|10973,10975
PO|10976,10978
once|10979,10983
a|10984,10985
day|10986,10989
.|10989,10990
<EOL>|10992,10993
5.|10993,10995
isosorbide|10996,11006
mononitrate|11007,11018
30|11019,11021
mg|11022,11024
Tablet|11025,11031
Extended|11032,11040
Release|11041,11048
24|11049,11051
hr|11052,11054
<EOL>|11055,11056
Sig|11056,11059
:|11059,11060
One|11061,11064
(|11065,11066
1|11066,11067
)|11067,11068
Tablet|11069,11075
Extended|11076,11084
Release|11085,11092
24|11093,11095
hr|11096,11098
PO|11099,11101
DAILY|11102,11107
(|11108,11109
Daily|11109,11114
)|11114,11115
.|11115,11116
<EOL>|11118,11119
6.|11119,11121
nitroglycerin|11122,11135
0.4|11136,11139
mg|11140,11142
Tablet|11143,11149
,|11149,11150
Sublingual|11151,11161
Sig|11162,11165
:|11165,11166
One|11167,11170
(|11171,11172
1|11172,11173
)|11173,11174
tablet|11175,11181
<EOL>|11183,11184
Sublingual|11184,11194
PRN|11195,11198
as|11200,11202
needed|11203,11209
for|11210,11213
chest|11214,11219
pain|11220,11224
.|11224,11225
<EOL>|11227,11228
7.|11228,11230
insulin|11231,11238
glargine|11239,11247
100|11248,11251
unit|11252,11256
/|11256,11257
mL|11257,11259
Solution|11260,11268
Sig|11269,11272
:|11272,11273
Eighty|11274,11280
(|11281,11282
80|11282,11284
)|11284,11285
units|11286,11291
<EOL>|11292,11293
Subcutaneous|11293,11305
at|11306,11308
bedtime|11309,11316
.|11316,11317
<EOL>|11319,11320
8.|11320,11322
insulin|11323,11330
lispro|11331,11337
100|11338,11341
unit|11342,11346
/|11346,11347
mL|11347,11349
Solution|11350,11358
Sig|11359,11362
:|11362,11363
Sliding|11364,11371
scale|11372,11377
units|11378,11383
<EOL>|11384,11385
of|11385,11387
insulin|11388,11395
Subcutaneous|11396,11408
three|11409,11414
times|11415,11420
a|11421,11422
day|11423,11426
:|11426,11427
As|11428,11430
directed|11431,11439
by|11440,11442
<EOL>|11443,11444
outpatient|11444,11454
provider|11455,11463
.|11464,11465
<EOL>|11467,11468
9.|11468,11470
albuterol|11471,11480
sulfate|11481,11488
90|11489,11491
mcg|11492,11495
/|11495,11496
actuation|11496,11505
HFA|11506,11509
Aerosol|11510,11517
Inhaler|11518,11525
Sig|11526,11529
:|11529,11530
<EOL>|11531,11532
Two|11532,11535
(|11536,11537
2|11537,11538
)|11538,11539
Puff|11540,11544
Inhalation|11545,11555
every|11556,11561
_|11562,11563
_|11563,11564
_|11564,11565
hours|11566,11571
as|11572,11574
needed|11575,11581
for|11582,11585
SOB|11586,11589
,|11589,11590
<EOL>|11591,11592
wheezing|11592,11600
.|11600,11601
<EOL>|11603,11604
10.|11604,11607
fluticasone|11608,11619
110|11620,11623
mcg|11624,11627
/|11627,11628
actuation|11628,11637
Aerosol|11638,11645
Sig|11646,11649
:|11649,11650
Two|11651,11654
(|11655,11656
2|11656,11657
)|11657,11658
Puff|11659,11663
<EOL>|11664,11665
Inhalation|11665,11675
BID|11676,11679
(|11680,11681
2|11681,11682
times|11683,11688
a|11689,11690
day|11691,11694
)|11694,11695
.|11695,11696
<EOL>|11698,11699
11.|11699,11702
pantoprazole|11703,11715
40|11716,11718
mg|11719,11721
Tablet|11722,11728
,|11728,11729
Delayed|11730,11737
Release|11738,11745
(|11746,11747
E.C|11747,11750
.|11750,11751
)|11751,11752
Sig|11753,11756
:|11756,11757
One|11758,11761
<EOL>|11762,11763
(|11763,11764
1|11764,11765
)|11765,11766
Tablet|11767,11773
,|11773,11774
Delayed|11775,11782
Release|11783,11790
(|11791,11792
E.C|11792,11795
.|11795,11796
)|11796,11797
PO|11798,11800
Q12H|11801,11805
(|11806,11807
every|11807,11812
12|11813,11815
hours|11816,11821
)|11821,11822
.|11822,11823
<EOL>|11825,11826
12.|11826,11829
oxycodone|11830,11839
-|11839,11840
acetaminophen|11840,11853
_|11854,11855
_|11855,11856
_|11856,11857
mg|11858,11860
Tablet|11861,11867
Sig|11868,11871
:|11871,11872
One|11873,11876
(|11877,11878
1|11878,11879
)|11879,11880
Tablet|11881,11887
<EOL>|11888,11889
PO|11889,11891
Q8H|11892,11895
(|11896,11897
every|11897,11902
8|11903,11904
hours|11905,11910
)|11910,11911
as|11912,11914
needed|11915,11921
for|11922,11925
pain|11926,11930
.|11930,11931
<EOL>|11933,11934
13.|11934,11937
cholecalciferol|11938,11953
(|11954,11955
vitamin|11955,11962
D3|11963,11965
)|11965,11966
1,000|11967,11972
unit|11973,11977
Capsule|11978,11985
Sig|11986,11989
:|11989,11990
One|11991,11994
(|11995,11996
1|11996,11997
)|11997,11998
<EOL>|11999,12000
Capsule|12000,12007
PO|12008,12010
once|12011,12015
a|12016,12017
day|12018,12021
.|12021,12022
<EOL>|12024,12025
14.|12025,12028
metronidazole|12029,12042
0.75|12043,12047
%|12048,12049
Lotion|12050,12056
Sig|12057,12060
:|12060,12061
One|12062,12065
(|12066,12067
1|12067,12068
)|12068,12069
application|12070,12081
<EOL>|12083,12084
Topical|12084,12091
as|12092,12094
directed|12095,12103
.|12104,12105
<EOL>|12107,12108
<EOL>|12108,12109
<EOL>|12110,12111
Discharge|12111,12120
Disposition|12121,12132
:|12132,12133
<EOL>|12133,12134
Home|12134,12138
<EOL>|12138,12139
<EOL>|12140,12141
Discharge|12141,12150
Diagnosis|12151,12160
:|12160,12161
<EOL>|12161,12162
Primary|12162,12169
diagnosis|12170,12179
:|12179,12180
<EOL>|12180,12181
Atypical|12181,12189
chest|12190,12195
pain|12196,12200
<EOL>|12200,12201
<EOL>|12201,12202
Secondary|12202,12211
diagnosis|12212,12221
:|12221,12222
<EOL>|12222,12223
Coronary|12223,12231
artery|12232,12238
disease|12239,12246
<EOL>|12247,12248
Hypertension|12248,12260
<EOL>|12260,12261
Hyperlipidemia|12261,12275
<EOL>|12275,12276
Type|12276,12280
2|12281,12282
Diabetes|12283,12291
Mellitus|12292,12300
<EOL>|12300,12301
<EOL>|12301,12302
<EOL>|12303,12304
Discharge|12304,12313
Condition|12314,12323
:|12323,12324
<EOL>|12324,12325
Mental|12325,12331
Status|12332,12338
:|12338,12339
Clear|12340,12345
and|12346,12349
coherent|12350,12358
.|12358,12359
<EOL>|12359,12360
Level|12360,12365
of|12366,12368
Consciousness|12369,12382
:|12382,12383
Alert|12384,12389
and|12390,12393
interactive|12394,12405
.|12405,12406
<EOL>|12406,12407
Activity|12407,12415
Status|12416,12422
:|12422,12423
Ambulatory|12424,12434
-|12435,12436
Independent|12437,12448
.|12448,12449
<EOL>|12449,12450
<EOL>|12450,12451
<EOL>|12452,12453
Discharge|12453,12462
Instructions|12463,12475
:|12475,12476
<EOL>|12476,12477
It|12477,12479
was|12480,12483
a|12484,12485
pleasure|12486,12494
taking|12495,12501
care|12502,12506
of|12507,12509
you|12510,12513
during|12514,12520
your|12521,12525
hospitalization|12526,12541
<EOL>|12542,12543
at|12543,12545
_|12546,12547
_|12547,12548
_|12548,12549
.|12549,12550
<EOL>|12551,12552
<EOL>|12552,12553
You|12553,12556
were|12557,12561
hospitalized|12562,12574
with|12575,12579
chest|12580,12585
pain|12586,12590
and|12591,12594
had|12595,12598
a|12599,12600
nuclear|12601,12608
stress|12609,12615
<EOL>|12616,12617
test|12617,12621
that|12622,12626
was|12627,12630
abnormal|12631,12639
.|12639,12640
You|12641,12644
subsequently|12645,12657
had|12658,12661
a|12662,12663
cardiac|12664,12671
<EOL>|12672,12673
catheterization|12673,12688
and|12689,12692
you|12693,12696
were|12697,12701
found|12702,12707
to|12708,12710
have|12711,12715
a|12716,12717
blockage|12718,12726
in|12727,12729
the|12730,12733
<EOL>|12734,12735
left|12735,12739
circumflex|12740,12750
coronary|12751,12759
artery|12760,12766
(|12767,12768
one|12768,12771
of|12772,12774
the|12775,12778
heart|12779,12784
vessels|12785,12792
)|12792,12793
.|12793,12794
<EOL>|12795,12796
<EOL>|12796,12797
Take|12797,12801
all|12802,12805
medication|12806,12816
as|12817,12819
instructed|12820,12830
.|12830,12831
Please|12832,12838
note|12839,12843
the|12844,12847
following|12848,12857
<EOL>|12858,12859
medication|12859,12869
changes|12870,12877
:|12877,12878
<EOL>|12878,12879
1|12879,12880
.|12880,12881
Stop|12882,12886
taking|12887,12893
your|12894,12898
potassium|12899,12908
supplement|12909,12919
for|12920,12923
now|12924,12927
,|12927,12928
as|12929,12931
your|12932,12936
<EOL>|12937,12938
potassium|12938,12947
levels|12948,12954
were|12955,12959
normal|12960,12966
in|12967,12969
the|12970,12973
hospital|12974,12982
.|12982,12983
<EOL>|12983,12984
2.|12984,12986
Increase|12987,12995
your|12996,13000
atorvastatin|13001,13013
(|13014,13015
lipitor|13015,13022
)|13022,13023
dose|13024,13028
from|13029,13033
40mg|13034,13038
to|13039,13041
80mg|13042,13046
<EOL>|13047,13048
daily|13048,13053
.|13053,13054
<EOL>|13054,13055
3|13055,13056
.|13056,13057
Stop|13058,13062
your|13063,13067
lisinopril|13068,13078
and|13079,13082
lasix|13083,13088
(|13089,13090
furosemide|13090,13100
)|13100,13101
until|13102,13107
otherwise|13108,13117
<EOL>|13118,13119
instructed|13119,13129
by|13130,13132
your|13133,13137
primary|13138,13145
care|13146,13150
physician|13151,13160
.|13160,13161
You|13162,13165
will|13166,13170
need|13171,13175
repeat|13176,13182
<EOL>|13183,13184
bloodwork|13184,13193
on|13194,13196
_|13197,13198
_|13198,13199
_|13199,13200
,|13200,13201
which|13202,13207
should|13208,13214
be|13215,13217
sent|13218,13222
to|13223,13225
your|13226,13230
<EOL>|13231,13232
primary|13232,13239
care|13240,13244
physician|13245,13254
,|13254,13255
_|13256,13257
_|13257,13258
_|13258,13259
.|13259,13260
<EOL>|13260,13261
<EOL>|13261,13262
Keep|13262,13266
all|13267,13270
hospital|13271,13279
follow|13280,13286
-|13286,13287
up|13287,13289
appointments|13290,13302
.|13302,13303
Your|13304,13308
up|13309,13311
-|13311,13312
coming|13312,13318
<EOL>|13319,13320
appointments|13320,13332
are|13333,13336
listed|13337,13343
below|13344,13349
.|13349,13350
<EOL>|13351,13352
<EOL>|13353,13354
Followup|13354,13362
Instructions|13363,13375
:|13375,13376
<EOL>|13376,13377
_|13377,13378
_|13378,13379
_|13379,13380
<EOL>|13380,13381

