 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
.|206,207
<EOL>|207,208
<EOL>|209,210
Chest|227,232
Pain|233,237
<EOL>|237,238
<EOL>|239,240
Major|240,245
Surgical|246,254
or|255,257
Invasive|258,266
Procedure|267,276
:|276,277
<EOL>|277,278
Exercise|278,286
Echocardiography|287,303
<EOL>|303,304
<EOL>|304,305
<EOL>|306,307
_|335,336
_|336,337
_|337,338
pmh|339,342
severe|343,349
known|350,355
CAD|356,359
s|360,361
/|361,362
p|362,363
CABG|364,368
and|369,372
multiple|373,381
caths|382,387
with|388,392
<EOL>|393,394
chronic|394,401
medicaly|402,410
managed|411,418
angina|419,425
,|425,426
_|427,428
_|428,429
_|429,430
,|430,431
HTN|432,435
,|435,436
DM|437,439
who|440,443
presents|444,452
with|453,457
<EOL>|458,459
atypical|459,467
chest|468,473
pain|474,478
.|478,479
<EOL>|481,482
.|482,483
<EOL>|485,486
Patient|486,493
has|494,497
history|498,505
of|506,508
CAD|509,512
and|513,516
is|517,519
s|520,521
/|521,522
p|522,523
3|524,525
vessel|526,532
CABG|533,537
(|538,539
LIMA|539,543
-|543,544
LAD|544,547
,|547,548
<EOL>|550,551
SVG|551,554
-|554,555
OM1|555,558
,|558,559
SVG|560,563
-|563,564
D1|564,566
)|566,567
by|568,570
Dr.|571,574
_|575,576
_|576,577
_|577,578
on|579,581
_|582,583
_|583,584
_|584,585
.|585,586
On|587,589
_|590,591
_|591,592
_|592,593
<EOL>|594,595
_|595,596
_|596,597
_|597,598
admitted|599,607
to|608,610
_|611,612
_|612,613
_|613,614
for|615,618
NSTEMI|619,625
and|626,629
had|630,633
cath|634,638
which|639,644
showed|645,651
<EOL>|652,653
occluded|653,661
graft|662,667
to|668,670
a|671,672
small|673,678
diagonal|679,687
branch|688,694
,|694,695
as|696,698
well|699,703
as|704,706
a|707,708
70|709,711
%|711,712
<EOL>|713,714
stenosis|714,722
in|723,725
the|726,729
LAD|730,733
stent|734,739
and|740,743
a|744,745
70|746,748
-|748,749
80|749,751
%|751,752
stenosis|753,761
at|762,764
the|765,768
LCx|769,772
<EOL>|773,774
origin|774,780
.|780,781
She|782,785
was|786,789
medically|790,799
managed|800,807
with|808,812
uptitration|813,824
of|825,827
her|828,831
BB|832,834
and|835,838
<EOL>|839,840
Imdur|840,845
and|846,849
initiation|850,860
of|861,863
losartan|864,872
for|873,876
better|877,883
BP|884,886
control|887,894
.|894,895
She|896,899
<EOL>|900,901
often|901,906
has|907,910
angina|911,917
at|918,920
rest|921,925
and|926,929
at|930,932
her|933,936
recent|937,943
baseline|944,952
takes|953,958
<EOL>|959,960
nitroglycerin|960,973
SL|974,976
approximately|977,990
twice|991,996
weekly|997,1003
.|1003,1004
<EOL>|1006,1007
.|1007,1008
<EOL>|1010,1011
Since|1011,1016
_|1017,1018
_|1018,1019
_|1019,1020
she|1021,1024
complains|1025,1034
of|1035,1037
frequent|1038,1046
chest|1047,1052
pains|1053,1058
which|1059,1064
are|1065,1068
<EOL>|1069,1070
different|1070,1079
from|1080,1084
her|1085,1088
chronic|1089,1096
angina|1097,1103
as|1104,1106
she|1107,1110
usually|1111,1118
ahs|1119,1122
chest|1123,1128
<EOL>|1129,1130
pressire|1130,1138
but|1139,1142
currently|1143,1152
feels|1153,1158
more|1159,1163
like|1164,1168
"|1169,1170
needle|1170,1176
pricks|1177,1183
"|1183,1184
,|1184,1185
pain|1186,1190
is|1191,1193
<EOL>|1194,1195
also|1195,1199
more|1200,1204
persistent|1205,1215
and|1216,1219
she|1220,1223
does|1224,1228
not|1229,1232
have|1233,1237
significant|1238,1249
relief|1250,1256
<EOL>|1257,1258
with|1258,1262
nitro|1263,1268
.|1268,1269
It|1270,1272
is|1273,1275
also|1276,1280
worse|1281,1286
with|1287,1291
deep|1292,1296
breathing|1297,1306
and|1307,1310
with|1311,1315
<EOL>|1316,1317
pressure|1317,1325
on|1326,1328
anterior|1329,1337
chest|1338,1343
.|1343,1344
She|1345,1348
states|1349,1355
it|1356,1358
does|1359,1363
not|1364,1367
feel|1368,1372
like|1373,1377
the|1378,1381
<EOL>|1382,1383
pain|1383,1387
she|1388,1391
had|1392,1395
before|1396,1402
her|1403,1406
CABG|1407,1411
.|1411,1412
Today|1413,1418
pain|1419,1423
was|1424,1427
_|1428,1429
_|1429,1430
_|1430,1431
and|1432,1435
remained|1436,1444
<EOL>|1445,1446
continous|1446,1455
.|1455,1456
It|1457,1459
was|1460,1463
accompanied|1464,1475
by|1476,1478
some|1479,1483
SOB|1484,1487
w|1488,1489
/|1489,1490
o|1490,1491
diaphoresis|1492,1503
,|1503,1504
<EOL>|1505,1506
lighthededness|1506,1520
,|1520,1521
nausea|1522,1528
,|1528,1529
v|1530,1531
or|1532,1534
palpitations|1535,1547
.|1547,1548
She|1549,1552
denies|1553,1559
paroxysmal|1560,1570
<EOL>|1571,1572
nocturnal|1572,1581
dyspnea|1582,1589
,|1589,1590
orthopnea|1591,1600
,|1600,1601
ankle|1602,1607
edema|1608,1613
,|1613,1614
palpitations|1615,1627
,|1627,1628
syncope|1629,1636
<EOL>|1637,1638
or|1638,1640
presyncope|1641,1651
.|1651,1652
<EOL>|1654,1655
.|1655,1656
<EOL>|1658,1659
She|1659,1662
says|1663,1667
that|1668,1672
she|1673,1676
has|1677,1680
been|1681,1685
feeling|1686,1693
more|1694,1698
cold|1699,1703
than|1704,1708
usual|1709,1714
recently|1715,1723
<EOL>|1724,1725
nut|1725,1728
denies|1729,1735
any|1736,1739
fevers|1740,1746
or|1747,1749
chills|1750,1756
.|1756,1757
She|1758,1761
has|1762,1765
a|1766,1767
chronic|1768,1775
productive|1776,1786
<EOL>|1787,1788
cough|1788,1793
.|1793,1794
She|1795,1798
denies|1799,1805
any|1806,1809
GI|1810,1812
,|1812,1813
GU|1814,1816
complaints|1817,1827
.|1827,1828
<EOL>|1830,1831
.|1831,1832
<EOL>|1834,1835
Of|1835,1837
note|1838,1842
patient|1843,1850
currently|1851,1860
being|1861,1866
work|1867,1871
up|1872,1874
for|1875,1878
memeory|1879,1886
loss|1887,1891
and|1892,1895
<EOL>|1896,1897
cognitive|1897,1906
impairment|1907,1917
.|1917,1918
<EOL>|1920,1921
.|1921,1922
<EOL>|1924,1925
ED|1925,1927
Course|1928,1934
19|1935,1937
:|1937,1938
33|1938,1940
4|1941,1942
97.9|1943,1947
69|1948,1950
117|1951,1954
/|1954,1955
76|1955,1957
16|1958,1960
96|1961,1963
%|1963,1964
ra|1965,1967
<EOL>|1969,1970
-|1970,1971
EKG|1972,1975
:|1975,1976
sinus|1977,1982
@|1983,1984
68|1985,1987
,|1987,1988
lateral|1989,1996
depressions|1997,2008
similar|2009,2016
to|2017,2019
prior|2020,2025
,|2025,2026
no|2027,2029
new|2030,2033
<EOL>|2034,2035
ischemic|2035,2043
chgs|2044,2048
.|2048,2049
Labs|2050,2054
unremarkable|2055,2067
,|2067,2068
trop|2069,2073
neg|2074,2077
X1|2078,2080
,|2080,2081
CXR|2082,2085
non|2086,2089
acute|2090,2095
.|2095,2096
<EOL>|2098,2099
<EOL>|2100,2101
1.|2123,2125
CARDIAC|2126,2133
RISK|2134,2138
FACTORS|2139,2146
:|2146,2147
(|2148,2149
-|2149,2150
)|2150,2151
Diabetes|2151,2159
,|2159,2160
(|2161,2162
+|2162,2163
)|2163,2164
Dyslipidemia|2164,2176
,|2176,2177
(|2178,2179
+|2179,2180
)|2180,2181
HTN|2181,2184
<EOL>|2186,2187
2.|2187,2189
CARDIAC|2190,2197
-|2209,2210
Coronary|2210,2218
artery|2219,2225
disease|2226,2233
<EOL>|2235,2236
-|2236,2237
Diastolic|2237,2246
congestive|2247,2257
heart|2258,2263
failure|2264,2271
<EOL>|2273,2274
-|2274,2275
CABG|2275,2279
:|2279,2280
CABG|2281,2285
x|2286,2287
3|2288,2289
(|2290,2291
Off|2291,2294
pump|2295,2299
coronary|2300,2308
artery|2309,2315
bypass|2316,2322
graft|2323,2328
x3|2329,2331
,|2331,2332
left|2333,2337
<EOL>|2339,2340
<EOL>|2340,2341
internal|2341,2349
mammary|2350,2357
artery|2358,2364
to|2365,2367
left|2368,2372
anterior|2373,2381
descending|2382,2392
artery|2393,2399
and|2400,2403
<EOL>|2405,2406
saphenous|2406,2415
vein|2416,2420
grafts|2421,2427
to|2428,2430
diagonal|2431,2439
,|2439,2440
and|2441,2444
obtuse|2445,2451
marginal|2452,2460
arteries|2461,2469
)|2469,2470
<EOL>|2471,2472
<EOL>|2473,2474
-|2474,2475
PERCUTANEOUS|2475,2487
CORONARY|2488,2496
INTERVENTIONS|2497,2510
:|2510,2511
BMS|2512,2515
to|2516,2518
proximal|2519,2527
LAD|2528,2531
<EOL>|2533,2534
_|2534,2535
_|2535,2536
_|2536,2537
,|2537,2538
DES|2539,2542
to|2543,2545
mid|2546,2549
LAD|2550,2553
_|2554,2555
_|2555,2556
_|2556,2557
,|2557,2558
DES|2559,2562
to|2563,2565
edge|2566,2570
ISR|2571,2574
of|2575,2577
mid|2578,2581
LAD|2582,2585
DES|2586,2589
and|2590,2593
<EOL>|2595,2596
stenosis|2596,2604
distal|2605,2611
to|2612,2614
stent|2615,2620
_|2621,2622
_|2622,2623
_|2623,2624
,|2624,2625
DES|2626,2629
to|2630,2632
OM1|2633,2636
,|2636,2637
_|2638,2639
_|2639,2640
_|2640,2641
<EOL>|2643,2644
-|2644,2645
PACING|2645,2651
/|2651,2652
ICD|2652,2655
:|2655,2656
none|2656,2660
<EOL>|2662,2663
Morbid|2663,2669
obesity|2670,2677
.|2677,2678
<EOL>|2680,2681
COPD|2681,2685
<EOL>|2687,2688
GERD|2688,2692
<EOL>|2694,2695
Right|2695,2700
rotator|2701,2708
cuff|2709,2713
injury|2714,2720
/|2720,2721
bursitis|2721,2729
<EOL>|2731,2732
Migraines|2732,2741
<EOL>|2743,2744
Depression|2744,2754
<EOL>|2756,2757
DJD|2757,2760
<EOL>|2762,2763
Hemorrhoids|2763,2774
<EOL>|2776,2777
Rosacea|2777,2784
<EOL>|2786,2787
<EOL>|2787,2788
<EOL>|2789,2790
:|2804,2805
<EOL>|2805,2806
_|2806,2807
_|2807,2808
_|2808,2809
<EOL>|2809,2810
:|2824,2825
<EOL>|2825,2826
She|2826,2829
was|2830,2833
a|2834,2835
ward|2836,2840
of|2841,2843
the|2844,2847
_|2848,2849
_|2849,2850
_|2850,2851
and|2852,2855
does|2856,2860
not|2861,2864
know|2865,2869
her|2870,2873
family|2874,2880
.|2880,2881
<EOL>|2883,2884
<EOL>|2884,2885
<EOL>|2886,2887
ADMISSION|2902,2911
EXAM|2912,2916
:|2916,2917
<EOL>|2917,2918
VS|2918,2920
:|2920,2921
T|2922,2923
=|2923,2924
98.1|2924,2928
BP|2929,2931
=|2931,2932
150|2932,2935
/|2935,2936
69|2936,2938
HR|2939,2941
=|2941,2942
71|2942,2944
RR|2945,2947
=|2947,2948
18|2948,2950
O2|2951,2953
sat|2954,2957
=|2957,2958
97RA|2958,2962
<EOL>|2964,2965
GENERAL|2965,2972
:|2972,2973
Oriented|2974,2982
x3|2983,2985
.|2985,2986
Mood|2987,2991
,|2991,2992
affect|2993,2999
appropriate|3000,3011
.|3011,3012
<EOL>|3014,3015
HEENT|3015,3020
:|3020,3021
NCAT|3022,3026
.|3026,3027
Sclera|3028,3034
anicteric|3035,3044
.|3044,3045
PERRL|3046,3051
,|3051,3052
EOMI|3053,3057
.|3057,3058
Conjunctiva|3059,3070
were|3071,3075
<EOL>|3076,3077
pink|3077,3081
,|3081,3082
no|3083,3085
pallor|3086,3092
or|3093,3095
cyanosis|3096,3104
of|3105,3107
the|3108,3111
oral|3112,3116
mucosa|3117,3123
.|3123,3124
No|3125,3127
xanthelasma|3128,3139
.|3139,3140
<EOL>|3142,3143
<EOL>|3143,3144
NECK|3144,3148
:|3148,3149
Supple|3150,3156
with|3157,3161
JVP|3162,3165
of|3166,3168
5|3169,3170
cm|3171,3173
.|3173,3174
<EOL>|3176,3177
Chest|3177,3182
:|3182,3183
significant|3184,3195
diffuse|3196,3203
TTP|3204,3207
over|3208,3212
anterior|3213,3221
chest|3222,3227
wall|3228,3232
.|3232,3233
<EOL>|3235,3236
CARDIAC|3236,3243
:|3243,3244
s|3245,3246
/|3246,3247
p|3247,3248
CABG|3249,3253
RRR|3254,3257
No|3258,3260
m|3261,3262
/|3262,3263
r|3263,3264
/|3264,3265
g|3265,3266
.|3266,3267
No|3268,3270
thrills|3271,3278
,|3278,3279
lifts|3280,3285
.|3285,3286
No|3287,3289
S3|3290,3292
or|3293,3295
S4|3296,3298
.|3298,3299
<EOL>|3301,3302
<EOL>|3302,3303
LUNGS|3303,3308
:|3308,3309
coarse|3310,3316
left|3317,3321
basilar|3322,3329
crackles|3330,3338
which|3339,3344
may|3345,3348
be|3349,3351
consistent|3352,3362
with|3363,3367
<EOL>|3368,3369
pleural|3369,3376
process|3377,3384
seen|3385,3389
on|3390,3392
CXR|3393,3396
,|3396,3397
otherwise|3398,3407
good|3408,3412
air|3413,3416
movement|3417,3425
with|3426,3430
no|3431,3433
<EOL>|3434,3435
wheezes|3435,3442
or|3443,3445
rhonchi|3446,3453
.|3453,3454
<EOL>|3456,3457
ABDOMEN|3457,3464
:|3464,3465
Soft|3466,3470
,|3470,3471
NTND|3472,3476
.|3476,3477
No|3478,3480
HSM|3481,3484
or|3485,3487
tenderness|3488,3498
.|3498,3499
Abd|3500,3503
aorta|3504,3509
not|3510,3513
<EOL>|3514,3515
enlarged|3515,3523
by|3524,3526
palpation|3527,3536
.|3536,3537
No|3538,3540
abdominal|3541,3550
bruits|3551,3557
.|3557,3558
<EOL>|3560,3561
EXTREMITIES|3561,3572
:|3572,3573
No|3574,3576
c|3577,3578
/|3578,3579
c|3579,3580
/|3580,3581
e|3581,3582
.|3582,3583
No|3584,3586
femoral|3587,3594
bruits|3595,3601
.|3601,3602
<EOL>|3604,3605
SKIN|3605,3609
:|3609,3610
No|3611,3613
stasis|3614,3620
dermatitis|3621,3631
,|3631,3632
ulcers|3633,3639
,|3639,3640
scars|3641,3646
,|3646,3647
or|3648,3650
xanthomas|3651,3660
.|3660,3661
<EOL>|3663,3664
PULSES|3664,3670
:|3670,3671
papable|3672,3679
throughout|3680,3690
<EOL>|3692,3693
Neuro|3693,3698
:|3698,3699
no|3700,3702
gross|3703,3708
deficits|3709,3717
.|3717,3718
<EOL>|3720,3721
<EOL>|3721,3722
DISCHARGE|3722,3731
EXAM|3732,3736
:|3736,3737
<EOL>|3737,3738
VS|3738,3740
:|3740,3741
T|3742,3743
=|3743,3744
98.6|3744,3748
BP|3749,3751
=|3751,3752
113|3752,3755
-|3755,3756
180|3756,3759
/|3759,3760
60|3760,3762
-|3762,3763
82|3763,3765
_|3766,3767
_|3767,3768
_|3768,3769
RR|3770,3772
=|3772,3773
20|3773,3775
O2|3776,3778
sat|3779,3782
=|3782,3783
99RA|3783,3787
<EOL>|3789,3790
GENERAL|3790,3797
:|3797,3798
Oriented|3799,3807
x3|3808,3810
.|3810,3811
Mood|3812,3816
appropriate|3817,3828
with|3829,3833
flat|3834,3838
affect|3839,3845
.|3845,3846
NAD|3848,3851
<EOL>|3853,3854
HEENT|3854,3859
:|3859,3860
NCAT|3861,3865
.|3865,3866
Sclera|3867,3873
anicteric|3874,3883
.|3883,3884
PERRL|3885,3890
,|3890,3891
EOMI|3892,3896
.|3896,3897
Conjunctiva|3898,3909
were|3910,3914
<EOL>|3915,3916
pink|3916,3920
,|3920,3921
no|3922,3924
pallor|3925,3931
or|3932,3934
cyanosis|3935,3943
of|3944,3946
the|3947,3950
oral|3951,3955
mucosa|3956,3962
.|3962,3963
No|3964,3966
xanthelasma|3967,3978
.|3978,3979
<EOL>|3981,3982
Left|3982,3986
cornea|3987,3993
with|3994,3998
scar|3999,4003
tissue|4004,4010
medial|4011,4017
to|4018,4020
_|4021,4022
_|4022,4023
_|4023,4024
.|4024,4025
<EOL>|4025,4026
NECK|4026,4030
:|4030,4031
Supple|4032,4038
with|4039,4043
flat|4044,4048
JVP|4049,4052
.|4052,4053
No|4055,4057
thyromegaly|4058,4069
.|4069,4070
<EOL>|4070,4071
CHEST|4071,4076
:|4076,4077
TTP|4078,4081
over|4082,4086
sternum|4087,4094
<EOL>|4094,4095
CARDIAC|4095,4102
:|4102,4103
Distant|4104,4111
heart|4112,4117
sounds|4118,4124
.|4124,4125
No|4126,4128
m|4129,4130
/|4130,4131
r|4131,4132
/|4132,4133
g|4133,4134
.|4134,4135
No|4136,4138
thrills|4139,4146
,|4146,4147
lifts|4148,4153
.|4153,4154
No|4155,4157
<EOL>|4158,4159
S3|4159,4161
or|4162,4164
S4|4165,4167
.|4167,4168
<EOL>|4170,4171
LUNGS|4171,4176
:|4176,4177
CTAB|4178,4182
no|4183,4185
wheezing|4186,4194
,|4194,4195
rales|4196,4201
,|4201,4202
rhonchi|4203,4210
<EOL>|4212,4213
ABDOMEN|4213,4220
:|4220,4221
Obese|4222,4227
,|4227,4228
soft|4229,4233
,|4233,4234
NTND|4235,4239
.|4239,4240
No|4241,4243
HSM|4244,4247
or|4248,4250
tenderness|4251,4261
.|4261,4262
Abd|4263,4266
aorta|4267,4272
not|4273,4276
<EOL>|4277,4278
enlarged|4278,4286
by|4287,4289
palpation|4290,4299
.|4299,4300
No|4301,4303
abdominal|4304,4313
bruits|4314,4320
.|4320,4321
<EOL>|4323,4324
EXTREMITIES|4324,4335
:|4335,4336
No|4337,4339
c|4340,4341
/|4341,4342
c|4342,4343
/|4343,4344
e|4344,4345
.|4345,4346
No|4347,4349
femoral|4350,4357
bruits|4358,4364
.|4364,4365
<EOL>|4367,4368
SKIN|4368,4372
:|4372,4373
No|4374,4376
stasis|4377,4383
dermatitis|4384,4394
,|4394,4395
ulcers|4396,4402
,|4402,4403
scars|4404,4409
,|4409,4410
or|4411,4413
xanthomas|4414,4423
.|4423,4424
<EOL>|4426,4427
PULSES|4427,4433
:|4433,4434
2|4435,4436
+|4436,4437
radial|4438,4444
/|4444,4445
DPP|4445,4448
<EOL>|4448,4449
Neuro|4449,4454
:|4454,4455
AOX3|4456,4460
.|4460,4461
non-focal|4462,4471
exam|4472,4476
.|4476,4477
<EOL>|4477,4478
<EOL>|4479,4480
Pertinent|4480,4489
Results|4490,4497
:|4497,4498
<EOL>|4498,4499
ADMISSION|4499,4508
LABS|4509,4513
:|4513,4514
<EOL>|4514,4515
<EOL>|4515,4516
_|4516,4517
_|4517,4518
_|4518,4519
09|4520,4522
:|4522,4523
03PM|4523,4527
BLOOD|4528,4533
WBC|4534,4537
-|4537,4538
7.7|4538,4541
RBC|4542,4545
-|4545,4546
3|4546,4547
.|4547,4548
89|4548,4550
*|4550,4551
Hgb|4552,4555
-|4555,4556
12.6|4556,4560
Hct|4561,4564
-|4564,4565
36.1|4565,4569
<EOL>|4570,4571
MCV|4571,4574
-|4574,4575
93|4575,4577
MCH|4578,4581
-|4581,4582
32|4582,4584
.|4584,4585
5|4585,4586
*|4586,4587
MCHC|4588,4592
-|4592,4593
34.9|4593,4597
RDW|4598,4601
-|4601,4602
12.3|4602,4606
Plt|4607,4610
_|4611,4612
_|4612,4613
_|4613,4614
<EOL>|4614,4615
_|4615,4616
_|4616,4617
_|4617,4618
10|4619,4621
:|4621,4622
47PM|4622,4626
BLOOD|4627,4632
_|4633,4634
_|4634,4635
_|4635,4636
PTT|4637,4640
-|4640,4641
28.2|4641,4645
_|4646,4647
_|4647,4648
_|4648,4649
<EOL>|4649,4650
_|4650,4651
_|4651,4652
_|4652,4653
09|4654,4656
:|4656,4657
03PM|4657,4661
BLOOD|4662,4667
Glucose|4668,4675
-|4675,4676
413|4676,4679
*|4679,4680
UreaN|4681,4686
-|4686,4687
19|4687,4689
Creat|4690,4695
-|4695,4696
1.1|4696,4699
Na|4700,4702
-|4702,4703
136|4703,4706
<EOL>|4707,4708
K|4708,4709
-|4709,4710
3.6|4710,4713
Cl|4714,4716
-|4716,4717
95|4717,4719
*|4719,4720
HCO3|4721,4725
-|4725,4726
28|4726,4728
AnGap|4729,4734
-|4734,4735
17|4735,4737
<EOL>|4737,4738
_|4738,4739
_|4739,4740
_|4740,4741
09|4742,4744
:|4744,4745
03PM|4745,4749
BLOOD|4750,4755
ALT|4756,4759
-|4759,4760
12|4760,4762
AST|4763,4766
-|4766,4767
12|4767,4769
AlkPhos|4770,4777
-|4777,4778
62|4778,4780
TotBili|4781,4788
-|4788,4789
0.5|4789,4792
<EOL>|4792,4793
_|4793,4794
_|4794,4795
_|4795,4796
09|4797,4799
:|4799,4800
03PM|4800,4804
BLOOD|4805,4810
Lipase|4811,4817
-|4817,4818
80|4818,4820
*|4820,4821
<EOL>|4821,4822
_|4822,4823
_|4823,4824
_|4824,4825
09|4826,4828
:|4828,4829
03PM|4829,4833
BLOOD|4834,4839
cTropnT|4840,4847
-|4847,4848
<|4848,4849
0|4849,4850
.|4850,4851
01|4851,4853
<EOL>|4853,4854
_|4854,4855
_|4855,4856
_|4856,4857
07|4858,4860
:|4860,4861
50AM|4861,4865
BLOOD|4866,4871
CK|4872,4874
-|4874,4875
MB|4875,4877
-|4877,4878
1|4878,4879
cTropnT|4880,4887
-|4887,4888
<|4888,4889
0|4889,4890
.|4890,4891
01|4891,4893
<EOL>|4893,4894
_|4894,4895
_|4895,4896
_|4896,4897
07|4898,4900
:|4900,4901
50AM|4901,4905
BLOOD|4906,4911
Calcium|4912,4919
-|4919,4920
8.7|4920,4923
Phos|4924,4928
-|4928,4929
3.7|4929,4932
Mg|4933,4935
-|4935,4936
1.8|4936,4939
<EOL>|4939,4940
<EOL>|4940,4941
CXR|4941,4944
_|4945,4946
_|4946,4947
_|4947,4948
:|4948,4949
<EOL>|4949,4950
:|4958,4959
<EOL>|4959,4960
<EOL>|4961,4962
Frontal|4962,4969
and|4970,4973
lateral|4974,4981
views|4982,4987
of|4988,4990
the|4991,4994
chest|4995,5000
.|5000,5001
There|5003,5008
is|5009,5011
persistent|5012,5022
<EOL>|5023,5024
blunting|5024,5032
of|5033,5035
left|5036,5040
costophrenic|5041,5053
angle|5054,5059
laterally|5060,5069
suggestive|5070,5080
of|5081,5083
<EOL>|5084,5085
underlying|5085,5095
scarring|5096,5104
or|5105,5107
pleural|5108,5115
thickening|5116,5126
.|5126,5127
The|5129,5132
lungs|5133,5138
are|5139,5142
<EOL>|5143,5144
otherwise|5144,5153
clear|5154,5159
.|5159,5160
Cardiomediastinal|5162,5179
silhouette|5180,5190
is|5191,5193
within|5194,5200
normal|5201,5207
<EOL>|5208,5209
limits|5209,5215
.|5215,5216
Median|5218,5224
sternotomy|5225,5235
wires|5236,5241
and|5242,5245
mediastinal|5246,5257
clips|5258,5263
again|5264,5269
<EOL>|5270,5271
noted|5271,5276
.|5276,5277
<EOL>|5277,5278
<EOL>|5279,5280
No|5294,5296
acute|5297,5302
cardiopulmonary|5303,5318
process|5319,5326
.|5326,5327
<EOL>|5327,5328
<EOL>|5328,5329
Exercise|5329,5337
Stress|5338,5344
_|5345,5346
_|5346,5347
_|5347,5348
:|5348,5349
<EOL>|5349,5350
IMPRESSION|5350,5360
:|5360,5361
Atypical|5362,5370
sudden|5371,5377
onset|5378,5383
of|5384,5386
chest|5387,5392
tightness|5393,5402
with|5403,5407
<EOL>|5408,5409
non-specific|5409,5421
ST|5422,5424
segment|5425,5432
changes|5433,5440
to|5441,5443
achieved|5444,5452
low|5453,5456
workload|5457,5465
.|5465,5466
<EOL>|5467,5468
Resting|5468,5475
mild|5476,5480
systolic|5481,5489
hypertension|5490,5502
with|5503,5507
a|5508,5509
blunted|5510,5517
hemodynamic|5518,5529
<EOL>|5530,5531
response|5531,5539
to|5540,5542
exercise|5543,5551
.|5551,5552
Echo|5553,5557
report|5558,5564
sent|5565,5569
separately|5570,5580
.|5580,5581
<EOL>|5581,5582
<EOL>|5582,5583
Exercise|5583,5591
Echo|5592,5596
_|5597,5598
_|5598,5599
_|5599,5600
:|5600,5601
<EOL>|5601,5602
IMPRESSION|5602,5612
:|5612,5613
Poor|5614,5618
functional|5619,5629
exercise|5630,5638
capacity|5639,5647
.|5647,5648
Non-specific|5649,5661
ECG|5662,5665
<EOL>|5666,5667
changes|5667,5674
in|5675,5677
the|5678,5681
absence|5682,5689
of|5690,5692
2D|5693,5695
echocardiographic|5696,5713
evidence|5714,5722
of|5723,5725
<EOL>|5726,5727
inducible|5727,5736
ischemia|5737,5745
to|5746,5748
achieved|5749,5757
low|5758,5761
workload|5762,5770
.|5770,5771
Resting|5772,5779
mild|5780,5784
<EOL>|5785,5786
systolic|5786,5794
hypertension|5795,5807
with|5808,5812
a|5813,5814
blunted|5815,5822
hemodynamic|5823,5834
response|5835,5843
to|5844,5846
<EOL>|5847,5848
physiologic|5848,5859
stress|5860,5866
.|5866,5867
<EOL>|5868,5869
<EOL>|5869,5870
DISCHARGE|5870,5879
LABS|5880,5884
:|5884,5885
<EOL>|5885,5886
<EOL>|5886,5887
_|5887,5888
_|5888,5889
_|5889,5890
07|5891,5893
:|5893,5894
50AM|5894,5898
BLOOD|5899,5904
WBC|5905,5908
-|5908,5909
7.0|5909,5912
RBC|5913,5916
-|5916,5917
3|5917,5918
.|5918,5919
80|5919,5921
*|5921,5922
Hgb|5923,5926
-|5926,5927
12.2|5927,5931
Hct|5932,5935
-|5935,5936
35|5936,5938
.|5938,5939
5|5939,5940
*|5940,5941
<EOL>|5942,5943
MCV|5943,5946
-|5946,5947
94|5947,5949
MCH|5950,5953
-|5953,5954
32|5954,5956
.|5956,5957
2|5957,5958
*|5958,5959
MCHC|5960,5964
-|5964,5965
34.5|5965,5969
RDW|5970,5973
-|5973,5974
11.9|5974,5978
Plt|5979,5982
_|5983,5984
_|5984,5985
_|5985,5986
<EOL>|5986,5987
_|5987,5988
_|5988,5989
_|5989,5990
07|5991,5993
:|5993,5994
25AM|5994,5998
BLOOD|5999,6004
Creat|6005,6010
-|6010,6011
0.9|6011,6014
Na|6015,6017
-|6017,6018
135|6018,6021
K|6022,6023
-|6023,6024
3.9|6024,6027
Cl|6028,6030
-|6030,6031
99|6031,6033
HCO3|6034,6038
-|6038,6039
26|6039,6041
<EOL>|6042,6043
AnGap|6043,6048
-|6048,6049
14|6049,6051
<EOL>|6051,6052
_|6052,6053
_|6053,6054
_|6054,6055
07|6056,6058
:|6058,6059
25AM|6059,6063
BLOOD|6064,6069
Phos|6070,6074
-|6074,6075
4.3|6075,6078
Mg|6079,6081
-|6081,6082
1|6082,6083
.|6083,6084
_|6084,6085
_|6085,6086
_|6086,6087
SSESSMENT|6087,6096
AND|6097,6100
PLAN|6101,6105
:|6105,6106
_|6107,6108
_|6108,6109
_|6109,6110
pmh|6111,6114
severe|6115,6121
known|6122,6127
CAD|6128,6131
s|6132,6133
/|6133,6134
p|6134,6135
CABG|6136,6140
with|6141,6145
<EOL>|6146,6147
chronic|6147,6154
angina|6156,6162
,|6162,6163
dCHF|6164,6168
,|6168,6169
HTN|6170,6173
,|6173,6174
DM|6175,6177
who|6178,6181
presents|6182,6190
with|6191,6195
chest|6196,6201
pain|6202,6206
<EOL>|6207,6208
concerning|6208,6218
for|6219,6222
crescendo|6223,6232
angina|6233,6239
.|6239,6240
<EOL>|6240,6241
<EOL>|6241,6242
ACTIVE|6242,6248
ISSUES|6249,6255
:|6255,6256
<EOL>|6256,6257
<EOL>|6259,6260
Chest|6260,6265
pain|6266,6270
:|6270,6271
patient|6272,6279
with|6280,6284
high|6285,6289
coronary|6290,6298
risk|6299,6303
,|6303,6304
however|6305,6312
recent|6313,6319
cat|6320,6323
<EOL>|6324,6325
6|6325,6326
months|6327,6333
ago|6334,6337
did|6338,6341
not|6342,6345
reveal|6346,6352
interveneable|6353,6366
disease|6367,6374
.|6374,6375
Fact|6377,6381
that|6382,6386
<EOL>|6387,6388
she|6388,6391
is|6392,6394
having|6395,6401
reproducability|6402,6417
on|6418,6420
physical|6421,6429
exam|6430,6434
suggests|6435,6443
non|6444,6447
<EOL>|6448,6449
cardiac|6449,6456
cause|6457,6462
,|6462,6463
however|6464,6471
symptoms|6472,6480
are|6481,6484
complicated|6485,6496
by|6497,6499
patient|6500,6507
's|6507,6509
<EOL>|6510,6511
history|6511,6518
of|6519,6521
cognitive|6522,6531
impairment|6532,6542
.|6542,6543
Given|6545,6550
known|6551,6556
CAD|6557,6560
with|6561,6565
70|6566,6568
%|6568,6569
<EOL>|6570,6571
stenosis|6571,6579
stress|6580,6586
echo|6587,6591
was|6592,6595
performed|6596,6605
to|6606,6608
assess|6609,6615
for|6616,6619
functional|6620,6630
<EOL>|6631,6632
abnormality|6632,6643
with|6644,6648
exertion|6649,6657
.|6657,6658
No|6660,6662
ECHO|6663,6667
abnormalities|6668,6681
were|6682,6686
noted|6687,6692
<EOL>|6693,6694
although|6694,6702
pt|6703,6705
reported|6706,6714
atypical|6715,6723
chest|6724,6729
pain|6730,6734
with|6735,6739
stress|6740,6746
.|6746,6747
She|6749,6752
was|6753,6756
<EOL>|6757,6758
continued|6758,6767
on|6768,6770
home|6771,6775
ASA|6776,6779
,|6779,6780
plavix|6781,6787
,|6787,6788
statin|6789,6795
,|6795,6796
nitrate|6797,6804
and|6805,6808
metoprolol|6809,6819
<EOL>|6820,6821
while|6821,6826
in|6827,6829
-|6829,6830
house|6830,6835
.|6835,6836
She|6838,6841
was|6842,6845
monitored|6846,6855
on|6856,6858
tele|6859,6863
without|6864,6871
any|6872,6875
alarms|6876,6882
.|6882,6883
<EOL>|6885,6886
She|6886,6889
was|6890,6893
discharged|6894,6904
home|6905,6909
after|6910,6915
a|6916,6917
negative|6918,6926
stress|6927,6933
to|6934,6936
follow|6937,6943
-|6943,6944
up|6944,6946
<EOL>|6947,6948
with|6948,6952
her|6953,6956
PCP|6957,6960
and|6961,6964
_|6965,6966
_|6966,6967
_|6967,6968
.|6968,6969
<EOL>|6969,6970
<EOL>|6970,6971
CHRONIC|6971,6978
ISSUES|6979,6985
:|6985,6986
<EOL>|6987,6988
<EOL>|6989,6990
#|6990,6991
Diastolic|6992,7001
CHF|7002,7005
(|7006,7007
EF|7007,7009
>|7009,7010
50|7010,7012
%|7012,7013
)|7013,7014
:|7014,7015
No|7016,7018
signs|7019,7024
of|7025,7027
fluid|7028,7033
overload|7034,7042
currently|7043,7052
.|7052,7053
<EOL>|7055,7056
Not|7056,7059
on|7060,7062
baseline|7063,7071
diuresis|7072,7080
.|7080,7081
She|7083,7086
was|7087,7090
continued|7091,7100
on|7101,7103
home|7104,7108
BB|7109,7111
and|7112,7115
_|7116,7117
_|7117,7118
_|7118,7119
<EOL>|7120,7121
and|7121,7124
monitored|7125,7134
daily|7135,7140
for|7141,7144
signs|7145,7150
of|7151,7153
decompensation|7154,7168
and|7169,7172
required|7173,7181
no|7182,7184
<EOL>|7185,7186
diuresis|7186,7194
.|7194,7195
<EOL>|7195,7196
<EOL>|7197,7198
#|7198,7199
Diabetes|7200,7208
:|7208,7209
HISS|7211,7215
in|7216,7218
-|7218,7219
house|7219,7224
,|7224,7225
she|7226,7229
was|7230,7233
also|7234,7238
continued|7239,7248
on|7249,7251
home|7252,7256
<EOL>|7257,7258
insulin|7258,7265
regimen|7266,7273
with|7274,7278
80|7279,7281
lantus|7282,7288
QHS|7289,7292
<EOL>|7294,7295
<EOL>|7296,7297
Medications|7297,7308
on|7309,7311
Admission|7312,7321
:|7321,7322
<EOL>|7322,7323
The|7323,7326
Preadmission|7327,7339
Medication|7340,7350
list|7351,7355
is|7356,7358
accurate|7359,7367
and|7368,7371
complete|7372,7380
.|7380,7381
<EOL>|7381,7382
1.|7382,7384
Losartan|7385,7393
Potassium|7394,7403
25|7404,7406
mg|7407,7409
PO|7410,7412
DAILY|7413,7418
<EOL>|7419,7420
2.|7420,7422
Aspirin|7423,7430
81|7431,7433
mg|7434,7436
PO|7437,7439
DAILY|7440,7445
<EOL>|7446,7447
3.|7447,7449
carisoprodol|7450,7462
*|7463,7464
NF|7464,7466
*|7466,7467
250|7468,7471
mg|7472,7474
Oral|7475,7479
qhs|7480,7483
spasm|7484,7489
<EOL>|7490,7491
Take|7491,7495
1|7496,7497
tablet|7498,7504
po|7505,7507
at|7508,7510
bedtime|7511,7518
PRN|7519,7522
muscle|7523,7529
spasm|7530,7535
<EOL>|7536,7537
4.|7537,7539
Pantoprazole|7540,7552
40|7553,7555
mg|7556,7558
PO|7559,7561
Q24H|7562,7566
<EOL>|7567,7568
5.|7568,7570
traZODONE|7571,7580
50|7581,7583
mg|7584,7586
PO|7587,7589
HS|7590,7592
<EOL>|7593,7594
6.|7594,7596
Oxycodone|7597,7606
-|7606,7607
Acetaminophen|7607,7620
(|7621,7622
5mg|7622,7625
-|7625,7626
325mg|7626,7631
)|7631,7632
1|7633,7634
TAB|7635,7638
PO|7639,7641
Q8H|7642,7645
:|7645,7646
PRN|7646,7649
pain|7650,7654
<EOL>|7655,7656
7.|7656,7658
Atorvastatin|7659,7671
40|7672,7674
mg|7675,7677
PO|7678,7680
DAILY|7681,7686
<EOL>|7687,7688
8.|7688,7690
Nitroglycerin|7691,7704
SL|7705,7707
0.4|7708,7711
mg|7712,7714
SL|7715,7717
PRN|7718,7721
chest|7722,7727
pain|7728,7732
<EOL>|7733,7734
9.|7734,7736
Metoprolol|7737,7747
Succinate|7748,7757
XL|7758,7760
200|7761,7764
mg|7765,7767
PO|7768,7770
DAILY|7771,7776
<EOL>|7777,7778
10.|7778,7781
Isosorbide|7782,7792
Mononitrate|7793,7804
(|7805,7806
Extended|7806,7814
Release|7815,7822
)|7822,7823
120|7824,7827
mg|7828,7830
PO|7831,7833
DAILY|7834,7839
<EOL>|7840,7841
11.|7841,7844
Clopidogrel|7845,7856
75|7857,7859
mg|7860,7862
PO|7863,7865
DAILY|7866,7871
<EOL>|7872,7873
12.|7873,7876
Fluticasone|7877,7888
Propionate|7889,7899
110mcg|7900,7906
2|7907,7908
PUFF|7909,7913
IH|7914,7916
BID|7917,7920
<EOL>|7921,7922
13|7922,7924
.|7924,7925
Other|7926,7931
90|7932,7934
Units|7935,7940
Bedtime|7941,7948
<EOL>|7948,7949
Insulin|7949,7956
SC|7957,7959
Sliding|7960,7967
Scale|7968,7973
using|7974,7979
HUM|7980,7983
InsulinMax|7984,7994
Dose|7995,7999
Override|8000,8008
<EOL>|8009,8010
Reason|8010,8016
:|8016,8017
Levemir|8018,8025
-|8025,8026
90|8027,8029
U|8030,8031
QHS|8032,8035
per|8036,8039
pharmacy|8040,8048
list|8049,8053
<EOL>|8053,8054
<EOL>|8054,8055
<EOL>|8056,8057
Discharge|8057,8066
Medications|8067,8078
:|8078,8079
<EOL>|8079,8080
1.|8080,8082
Aspirin|8083,8090
81|8091,8093
mg|8094,8096
PO|8097,8099
DAILY|8100,8105
<EOL>|8106,8107
2.|8107,8109
Atorvastatin|8110,8122
40|8123,8125
mg|8126,8128
PO|8129,8131
DAILY|8132,8137
<EOL>|8138,8139
3.|8139,8141
Clopidogrel|8142,8153
75|8154,8156
mg|8157,8159
PO|8160,8162
DAILY|8163,8168
<EOL>|8169,8170
4.|8170,8172
Fluticasone|8173,8184
Propionate|8185,8195
110mcg|8196,8202
2|8203,8204
PUFF|8205,8209
IH|8210,8212
BID|8213,8216
<EOL>|8217,8218
5.|8218,8220
Other|8221,8226
90|8227,8229
Units|8230,8235
Bedtime|8236,8243
<EOL>|8243,8244
Insulin|8244,8251
SC|8252,8254
Sliding|8255,8262
Scale|8263,8268
using|8269,8274
HUM|8275,8278
InsulinMax|8279,8289
Dose|8290,8294
Override|8295,8303
<EOL>|8304,8305
Reason|8305,8311
:|8311,8312
Levemir|8313,8320
-|8320,8321
90|8322,8324
U|8325,8326
QHS|8327,8330
per|8331,8334
pharmacy|8335,8343
list|8344,8348
<EOL>|8348,8349
<EOL>|8349,8350
6.|8350,8352
Losartan|8353,8361
Potassium|8362,8371
25|8372,8374
mg|8375,8377
PO|8378,8380
DAILY|8381,8386
<EOL>|8387,8388
7.|8388,8390
Nitroglycerin|8391,8404
SL|8405,8407
0.4|8408,8411
mg|8412,8414
SL|8415,8417
PRN|8418,8421
chest|8422,8427
pain|8428,8432
<EOL>|8433,8434
8.|8434,8436
Pantoprazole|8437,8449
40|8450,8452
mg|8453,8455
PO|8456,8458
Q24H|8459,8463
<EOL>|8464,8465
9.|8465,8467
traZODONE|8468,8477
50|8478,8480
mg|8481,8483
PO|8484,8486
HS|8487,8489
<EOL>|8490,8491
10.|8491,8494
carisoprodol|8495,8507
*|8508,8509
NF|8509,8511
*|8511,8512
250|8513,8516
mg|8517,8519
Oral|8520,8524
qhs|8525,8528
spasm|8529,8534
<EOL>|8535,8536
11|8536,8538
.|8538,8539
Metoprolol|8540,8550
Succinate|8551,8560
XL|8561,8563
200|8564,8567
mg|8568,8570
PO|8571,8573
DAILY|8574,8579
<EOL>|8580,8581
12.|8581,8584
Oxycodone|8585,8594
-|8594,8595
Acetaminophen|8595,8608
(|8609,8610
5mg|8610,8613
-|8613,8614
325mg|8614,8619
)|8619,8620
1|8621,8622
TAB|8623,8626
PO|8627,8629
Q8H|8630,8633
:|8633,8634
PRN|8634,8637
pain|8638,8642
<EOL>|8643,8644
13|8644,8646
.|8646,8647
Isosorbide|8648,8658
Mononitrate|8659,8670
(|8671,8672
Extended|8672,8680
Release|8681,8688
)|8688,8689
90|8690,8692
mg|8693,8695
PO|8696,8698
DAILY|8699,8704
<EOL>|8705,8706
<EOL>|8706,8707
<EOL>|8708,8709
Discharge|8709,8718
Disposition|8719,8730
:|8730,8731
<EOL>|8731,8732
Home|8732,8736
<EOL>|8736,8737
<EOL>|8738,8739
Discharge|8739,8748
Diagnosis|8749,8758
:|8758,8759
<EOL>|8759,8760
Atypical|8760,8768
Chest|8769,8774
Pain|8775,8779
<EOL>|8779,8780
<EOL>|8780,8781
<EOL>|8782,8783
Level|8804,8809
of|8810,8812
Consciousness|8813,8826
:|8826,8827
Alert|8828,8833
and|8834,8837
interactive|8838,8849
.|8849,8850
<EOL>|8850,8851
Mental|8851,8857
Status|8858,8864
:|8864,8865
Confused|8866,8874
-|8875,8876
sometimes|8877,8886
.|8886,8887
<EOL>|8887,8888
Activity|8888,8896
Status|8897,8903
:|8903,8904
Ambulatory|8905,8915
-|8916,8917
Independent|8918,8929
.|8929,8930
<EOL>|8930,8931
<EOL>|8931,8932
<EOL>|8933,8934
Ms.|8958,8961
_|8962,8963
_|8963,8964
_|8964,8965
-|8965,8966
<EOL>|8966,8967
<EOL>|8967,8968
You|8968,8971
came|8972,8976
to|8977,8979
the|8980,8983
hospital|8984,8992
with|8993,8997
chest|8998,9003
pain|9004,9008
.|9008,9009
You|9011,9014
had|9015,9018
lab|9019,9022
chests|9023,9029
<EOL>|9030,9031
and|9031,9034
EKG|9035,9038
's|9038,9040
that|9041,9045
were|9046,9050
reassuring|9051,9061
that|9062,9066
you|9067,9070
were|9071,9075
not|9076,9079
having|9080,9086
a|9087,9088
heart|9089,9094
<EOL>|9095,9096
attack|9096,9102
.|9102,9103
While|9105,9110
you|9111,9114
were|9115,9119
here|9120,9124
,|9124,9125
you|9126,9129
had|9130,9133
a|9134,9135
stress|9136,9142
test|9143,9147
which|9148,9153
did|9154,9157
<EOL>|9158,9159
not|9159,9162
suggest|9163,9170
any|9171,9174
evidence|9175,9183
of|9184,9186
worsening|9187,9196
coronary|9197,9205
artery|9206,9212
disease|9213,9220
.|9220,9221
<EOL>|9223,9224
Your|9224,9228
chest|9229,9234
pain|9235,9239
was|9240,9243
reproducible|9244,9256
with|9257,9261
touching|9262,9270
your|9271,9275
chest|9276,9281
,|9281,9282
which|9283,9288
<EOL>|9289,9290
is|9290,9292
not|9293,9296
typical|9297,9304
of|9305,9307
coronary|9308,9316
artery|9317,9323
disease|9324,9331
pain|9332,9336
.|9336,9337
This|9339,9343
likely|9344,9350
is|9351,9353
<EOL>|9354,9355
related|9355,9362
to|9363,9365
musculoskeletal|9366,9381
pain|9382,9386
.|9386,9387
<EOL>|9389,9390
Some|9390,9394
changes|9395,9402
have|9403,9407
been|9408,9412
made|9413,9417
to|9418,9420
your|9421,9425
medication|9426,9436
list|9437,9441
.|9441,9442
Please|9444,9450
<EOL>|9451,9452
followup|9452,9460
with|9461,9465
your|9466,9470
cardiologist|9471,9483
for|9484,9487
further|9488,9495
medication|9496,9506
changes|9507,9514
.|9514,9515
<EOL>|9515,9516
<EOL>|9517,9518
Followup|9518,9526
Instructions|9527,9539
:|9539,9540
<EOL>|9540,9541
_|9541,9542
_|9542,9543
_|9543,9544
<EOL>|9544,9545

