 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|184,193|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|184,193|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|196,218|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|204,208|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|204,208|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|204,218|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|221,230|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|Chief Complaint|256,261|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Chief Complaint|256,261|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Chief Complaint|278,283|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Chief Complaint|278,283|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Chief Complaint|278,283|false|false|false|C0010200|Coughing|cough
Finding|Classification|Chief Complaint|286,291|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|292,300|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|292,300|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|304,322|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|313,322|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|313,322|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|313,322|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|313,322|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|372,375|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|History of Present Illness|377,380|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|377,380|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|377,380|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|377,380|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|377,380|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|377,380|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|377,380|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|382,386|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|382,386|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|382,386|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Sign or Symptom|History of Present Illness|391,397|false|false|false|C0015967|Fever|fevers
Drug|Organic Chemical|History of Present Illness|414,419|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|414,419|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|414,419|false|false|false|C0010200|Coughing|cough
Finding|Functional Concept|History of Present Illness|462,467|false|false|false|C1442792|State|state
Finding|Finding|History of Present Illness|462,477|false|false|false|C0683314|personal health|state of health
Finding|Idea or Concept|History of Present Illness|471,477|false|false|false|C0018684|Health|health
Drug|Organic Chemical|History of Present Illness|518,523|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|518,523|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|518,523|false|false|false|C0010200|Coughing|cough
Finding|Body Substance|History of Present Illness|539,545|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|History of Present Illness|539,545|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Drug|Organic Chemical|History of Present Illness|562,572|false|false|false|C0723110|Robitussin|robitussin
Drug|Pharmacologic Substance|History of Present Illness|562,572|false|false|false|C0723110|Robitussin|robitussin
Disorder|Disease or Syndrome|History of Present Illness|585,588|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|History of Present Illness|585,588|false|false|false|C2346952|Bachelor of Education|bed
Finding|Idea or Concept|History of Present Illness|608,612|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Classification|History of Present Illness|629,636|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|general
Procedure|Health Care Activity|History of Present Illness|629,636|false|false|false|C3812897|General medical service|general
Finding|Sign or Symptom|History of Present Illness|629,644|false|false|false|C0231218|Malaise|general malaise
Finding|Sign or Symptom|History of Present Illness|637,644|false|false|false|C0231218|Malaise|malaise
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|646,651|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|646,651|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|646,651|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|646,651|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|646,651|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|646,651|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|History of Present Illness|646,662|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Finding|Pathologic Function|History of Present Illness|652,662|false|false|false|C0700148|Congestion|congestion
Finding|Finding|History of Present Illness|680,696|false|false|false|C0239134|Productive Cough|productive cough
Drug|Organic Chemical|History of Present Illness|691,696|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|691,696|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|691,696|false|false|false|C0010200|Coughing|cough
Drug|Inorganic Chemical|History of Present Illness|746,751|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|History of Present Illness|746,751|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|History of Present Illness|746,751|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|746,751|false|false|false|C0020311|Hydrotherapy|water
Finding|Finding|History of Present Illness|752,760|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|752,760|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|780,788|false|false|false|C0042963|Vomiting|vomiting
Attribute|Clinical Attribute|History of Present Illness|798,804|true|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|798,804|true|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|818,824|true|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|History of Present Illness|826,832|false|false|false|C0085593|Chills|chills
Finding|Body Substance|History of Present Illness|836,842|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|836,842|true|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|852,856|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|852,856|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|852,856|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|History of Present Illness|874,877|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|874,877|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|874,877|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|874,877|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|874,877|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|874,877|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|874,877|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|874,877|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|History of Present Illness|874,877|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|874,877|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Drug|Biomedical or Dental Material|History of Present Illness|899,903|false|false|false|C1999262|Pack|pack
Event|Activity|History of Present Illness|899,903|false|false|false|C2828395|Packing (action)|pack
Finding|Functional Concept|History of Present Illness|910,918|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|910,918|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Attribute|Clinical Attribute|History of Present Illness|948,952|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|948,952|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|948,952|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|958,966|false|false|false|C0010200|Coughing|coughing
Anatomy|Body Location or Region|History of Present Illness|985,992|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|History of Present Illness|985,992|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|History of Present Illness|985,992|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Location or Region|History of Present Illness|985,996|false|false|false|C0000726|Abdomen|abdomen and
Anatomy|Body Location or Region|History of Present Illness|997,1002|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|997,1002|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Location or Region|History of Present Illness|997,1008|false|false|false|C0446470|Surface region of lower chest|lower chest
Anatomy|Body Location or Region|History of Present Illness|1003,1008|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1003,1008|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Space or Junction|History of Present Illness|1024,1029|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|History of Present Illness|1024,1029|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|History of Present Illness|1024,1029|false|false|false|C0575044|Joint problem|joint
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1033,1039|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|History of Present Illness|1033,1039|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Sign or Symptom|History of Present Illness|1033,1044|false|false|false|C0231528|Myalgia|muscle pain
Attribute|Clinical Attribute|History of Present Illness|1040,1044|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1040,1044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1040,1044|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|1068,1071|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1068,1071|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1068,1071|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1068,1071|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1068,1071|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1068,1071|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1068,1071|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1068,1071|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|History of Present Illness|1068,1071|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1068,1071|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|History of Present Illness|1079,1082|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1079,1082|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Procedure|Health Care Activity|History of Present Illness|1086,1095|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|History of Present Illness|1105,1108|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1105,1108|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1105,1108|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1105,1108|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1105,1108|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1105,1108|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1105,1108|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1105,1108|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|History of Present Illness|1105,1108|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1105,1108|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|History of Present Illness|1112,1118|false|false|false|C1549636|Address type - Office|office
Finding|Pathologic Function|History of Present Illness|1123,1130|false|false|false|C0242184|Hypoxia|hypoxic
Disorder|Disease or Syndrome|History of Present Illness|1165,1168|false|false|false|C0021400|Influenza|flu
Finding|Gene or Genome|History of Present Illness|1165,1168|false|false|false|C3811318|ZMYND10 wt Allele|flu
Drug|Immunologic Factor|History of Present Illness|1165,1176|false|false|false|C0021403|Influenza virus vaccine|flu vaccine
Drug|Pharmacologic Substance|History of Present Illness|1165,1176|false|false|false|C0021403|Influenza virus vaccine|flu vaccine
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1169,1176|false|false|false|C0042210;C5399710|Vaccine [APC];Vaccines|vaccine
Drug|Immunologic Factor|History of Present Illness|1169,1176|false|false|false|C0042210;C5399710|Vaccine [APC];Vaccines|vaccine
Drug|Pharmacologic Substance|History of Present Illness|1169,1176|false|false|false|C0042210;C5399710|Vaccine [APC];Vaccines|vaccine
Finding|Idea or Concept|History of Present Illness|1183,1187|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|1183,1187|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Drug|Immunologic Factor|History of Present Illness|1192,1201|false|false|false|C0071315|Pneumovax|pneumovax
Drug|Pharmacologic Substance|History of Present Illness|1192,1201|false|false|false|C0071315|Pneumovax|pneumovax
Finding|Idea or Concept|History of Present Illness|1207,1211|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|1207,1211|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Sign or Symptom|History of Present Illness|1213,1219|false|false|false|C0043144|Wheezing|wheezy
Finding|Functional Concept|History of Present Illness|1223,1227|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1223,1227|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|History of Present Illness|1275,1283|false|false|false|C0277797|Apyrexial|afebrile
Finding|Functional Concept|History of Present Illness|1304,1308|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|1304,1308|false|false|false|C0582103|Medical Examination|exam
Finding|Sign or Symptom|History of Present Illness|1313,1320|false|false|false|C0043144|Wheezing|wheezes
Finding|Finding|History of Present Illness|1327,1336|false|false|false|C0857465|Peak flow|peak flow
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1332,1336|false|false|false|C0806140|Flow|flow
Drug|Biomedical or Dental Material|History of Present Illness|1348,1356|true|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|1348,1356|true|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Intellectual Product|History of Present Illness|1376,1385|false|false|false|C0876929|Sentence|sentences
Disorder|Congenital Abnormality|History of Present Illness|1394,1410|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|History of Present Illness|1394,1414|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1404,1410|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|History of Present Illness|1404,1410|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|History of Present Illness|1411,1414|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|History of Present Illness|1411,1414|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Attribute|Clinical Attribute|History of Present Illness|1437,1442|false|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|1437,1442|false|false|false|C0013604|Edema|edema
Disorder|Disease or Syndrome|History of Present Illness|1445,1448|false|false|false|C0021400|Influenza|Flu
Finding|Gene or Genome|History of Present Illness|1445,1448|false|false|false|C3811318|ZMYND10 wt Allele|Flu
Procedure|Diagnostic Procedure|History of Present Illness|1449,1455|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Procedure|Laboratory Procedure|History of Present Illness|1449,1455|false|false|false|C0199230;C0220908;C0430054;C1710031|Disease Screening;Screening for cancer;Screening procedure;Toxicology screen, general (procedure)|screen
Procedure|Diagnostic Procedure|History of Present Illness|1472,1475|false|false|false|C0039985|Plain chest X-ray|CXR
Drug|Biomedical or Dental Material|History of Present Illness|1526,1530|false|false|false|C1300458|Nebulizer solution|nebs
Drug|Hormone|History of Present Illness|1532,1536|false|false|false|C0032952;C0044955|prednisone;prednylidene|pred
Drug|Organic Chemical|History of Present Illness|1532,1536|false|false|false|C0032952;C0044955|prednisone;prednylidene|pred
Drug|Pharmacologic Substance|History of Present Illness|1532,1536|false|false|false|C0032952;C0044955|prednisone;prednylidene|pred
Disorder|Disease or Syndrome|Past Medical History|1569,1575|false|false|false|C0004096|Asthma|ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1579,1591|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|1595,1609|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Finding|Finding|Past Medical History|1595,1609|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Finding|Sign or Symptom|Past Medical History|1613,1621|false|false|false|C0018681|Headache|HEADACHE
Disorder|Disease or Syndrome|Past Medical History|1625,1639|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Finding|Finding|Past Medical History|1643,1651|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|1643,1662|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|1652,1657|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1652,1657|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|1652,1662|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|1652,1662|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|1658,1662|false|true|false|C2598155||PAIN
Finding|Functional Concept|Past Medical History|1658,1662|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|1658,1662|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Drug|Hazardous or Poisonous Substance|Past Medical History|1666,1673|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Past Medical History|1666,1673|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Past Medical History|1666,1673|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Past Medical History|1666,1673|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1666,1679|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1674,1679|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Past Medical History|1674,1679|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Past Medical History|1674,1679|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Finding|Past Medical History|1683,1691|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Idea or Concept|Past Medical History|1683,1691|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Finding|Past Medical History|1683,1697|false|false|false|C0742257|chest abnormal|ABNORMAL CHEST
Finding|Finding|Past Medical History|1683,1702|false|false|false|C0436503|Standard chest X-ray abnormal|ABNORMAL CHEST XRAY
Anatomy|Body Location or Region|Past Medical History|1692,1697|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1692,1697|false|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|Past Medical History|1692,1702|false|false|false|C0039985|Plain chest X-ray|CHEST XRAY
Phenomenon|Natural Phenomenon or Process|Past Medical History|1698,1702|false|false|false|C0043309|Roentgen Rays|XRAY
Procedure|Diagnostic Procedure|Past Medical History|1698,1702|false|false|false|C0043299|Diagnostic radiologic examination|XRAY
Disorder|Disease or Syndrome|Past Medical History|1706,1710|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1706,1710|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Past Medical History|1706,1710|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|Family Medical History|1751,1757|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|1764,1767|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Conceptual Entity|Family Medical History|1770,1776|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1770,1776|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Conceptual Entity|Family Medical History|1787,1794|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1787,1794|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Conceptual Entity|Family Medical History|1802,1809|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1802,1809|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Finding|Family Medical History|1820,1828|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|1820,1828|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|1820,1828|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|1837,1846|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1925,1930|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Family Medical History|1925,1930|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Family Medical History|1925,1930|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Family Medical History|1925,1930|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Family Medical History|1925,1930|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Family Medical History|1925,1930|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1931,1938|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|Family Medical History|1931,1938|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Family Medical History|1931,1938|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Attribute|Clinical Attribute|Family Medical History|1948,1959|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Family Medical History|1948,1959|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Family Medical History|1948,1959|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Family Medical History|1948,1959|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|Family Medical History|1948,1968|true|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|Family Medical History|1960,1968|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|1960,1968|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|1969,1974|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1977,1980|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|1977,1980|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1985,1988|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|1985,1988|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Family Medical History|1985,1988|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|Family Medical History|1993,1996|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|Family Medical History|1998,2002|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Family Medical History|1998,2002|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Family Medical History|1998,2002|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|Family Medical History|1998,2009|false|false|false|C2230237|Supple neck|neck supple
Finding|Functional Concept|Family Medical History|2003,2009|false|false|false|C0332254|Supple|supple
Finding|Finding|Family Medical History|2039,2046|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|Family Medical History|2055,2059|true|false|false|C0232267|Pericardial friction rub|rubs
Procedure|Health Care Activity|Family Medical History|2061,2065|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Drug|Organic Chemical|Family Medical History|2067,2071|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Finding|Family Medical History|2075,2083|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Sign or Symptom|Family Medical History|2087,2094|true|false|false|C0043144|Wheezing|wheezes
Finding|Idea or Concept|Family Medical History|2096,2100|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Organism Function|Family Medical History|2101,2112|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|Family Medical History|2113,2119|false|false|false|C0015264|Exertion|effort
Finding|Gene or Genome|Family Medical History|2130,2135|false|false|false|C1424898|RXFP2 gene|great
Drug|Inorganic Chemical|Family Medical History|2136,2139|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|2136,2139|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|2136,2139|false|true|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Family Medical History|2136,2139|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|2136,2139|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|2136,2139|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Family Medical History|2136,2148|false|true|false|C0001868|Air Movements|air movement
Finding|Organism Function|Family Medical History|2140,2148|false|true|false|C0026649|Movement|movement
Finding|Organism Function|Family Medical History|2169,2179|false|false|false|C0231800|Expiration, Respiratory|expiratory
Anatomy|Body Location or Region|Family Medical History|2187,2190|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|Family Medical History|2187,2190|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|Family Medical History|2192,2196|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|Family Medical History|2216,2219|false|false|false|C5848551|Neg - answer|neg
Finding|Gene or Genome|Family Medical History|2220,2223|false|false|false|C1537594|LRRC4B gene|HSM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2225,2236|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|Family Medical History|2246,2251|true|false|false|C1717255||edema
Finding|Pathologic Function|Family Medical History|2246,2251|true|false|false|C0013604|Edema|edema
Finding|Gene or Genome|Family Medical History|2253,2256|false|false|false|C1843919|PDSS1 gene|DPs
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2258,2261|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Enzyme|Family Medical History|2258,2261|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Organic Chemical|Family Medical History|2258,2261|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Pharmacologic Substance|Family Medical History|2258,2261|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Finding|Gene or Genome|Family Medical History|2258,2261|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Finding|Intellectual Product|Family Medical History|2258,2261|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Anatomy|Body System|Family Medical History|2266,2270|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|Family Medical History|2266,2270|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|Family Medical History|2266,2270|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|Family Medical History|2266,2270|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|Family Medical History|2266,2270|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Sign or Symptom|Family Medical History|2286,2292|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2299,2304|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Anatomy|Body System|Family Medical History|2306,2309|false|false|false|C3714787|Central Nervous System|CNs
Finding|Finding|Family Medical History|2317,2323|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Body Substance|Family Medical History|2329,2338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|2329,2338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|2329,2338|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|2329,2338|false|false|false|C0030685|Patient Discharge|DISCHARGE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2417,2422|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Family Medical History|2417,2422|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Family Medical History|2417,2422|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Family Medical History|2417,2422|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Family Medical History|2417,2422|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Family Medical History|2417,2422|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2423,2430|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|Family Medical History|2423,2430|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Family Medical History|2423,2430|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Attribute|Clinical Attribute|Family Medical History|2440,2451|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Family Medical History|2440,2451|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Family Medical History|2440,2451|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Family Medical History|2440,2451|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|Family Medical History|2440,2460|true|false|false|C0476273|Respiratory distress|respiratory distress
Finding|Finding|Family Medical History|2452,2460|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|Family Medical History|2452,2460|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|Family Medical History|2461,2466|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2469,2472|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|2469,2472|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2477,2480|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|2477,2480|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Family Medical History|2477,2480|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|Family Medical History|2485,2488|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|Family Medical History|2490,2494|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Family Medical History|2490,2494|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Family Medical History|2490,2494|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|Family Medical History|2490,2501|false|false|false|C2230237|Supple neck|neck supple
Finding|Functional Concept|Family Medical History|2495,2501|false|false|false|C0332254|Supple|supple
Finding|Finding|Family Medical History|2531,2538|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|Family Medical History|2547,2551|true|false|false|C0232267|Pericardial friction rub|rubs
Procedure|Health Care Activity|Family Medical History|2553,2557|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Drug|Organic Chemical|Family Medical History|2559,2563|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Finding|Family Medical History|2567,2575|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Sign or Symptom|Family Medical History|2579,2586|true|false|false|C0043144|Wheezing|wheezes
Finding|Idea or Concept|Family Medical History|2588,2592|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Finding|Organism Function|Family Medical History|2593,2604|false|false|false|C0004048|Inspiration (function)|inspiratory
Finding|Organism Function|Family Medical History|2605,2611|false|false|false|C0015264|Exertion|effort
Finding|Gene or Genome|Family Medical History|2622,2627|false|false|false|C1424898|RXFP2 gene|great
Drug|Inorganic Chemical|Family Medical History|2628,2631|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|2628,2631|false|true|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|2628,2631|false|true|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Family Medical History|2628,2631|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|2628,2631|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|2628,2631|false|true|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Family Medical History|2628,2640|false|true|false|C0001868|Air Movements|air movement
Finding|Organism Function|Family Medical History|2632,2640|false|true|false|C0026649|Movement|movement
Finding|Organism Function|Family Medical History|2661,2671|false|false|false|C0231800|Expiration, Respiratory|expiratory
Anatomy|Body Location or Region|Family Medical History|2679,2682|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|Family Medical History|2679,2682|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|Family Medical History|2684,2688|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|Family Medical History|2708,2711|false|false|false|C5848551|Neg - answer|neg
Finding|Gene or Genome|Family Medical History|2712,2715|false|false|false|C1537594|LRRC4B gene|HSM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2717,2728|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|Family Medical History|2738,2743|true|false|false|C1717255||edema
Finding|Pathologic Function|Family Medical History|2738,2743|true|false|false|C0013604|Edema|edema
Finding|Gene or Genome|Family Medical History|2745,2748|false|false|false|C1843919|PDSS1 gene|DPs
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2750,2753|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Enzyme|Family Medical History|2750,2753|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Organic Chemical|Family Medical History|2750,2753|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Pharmacologic Substance|Family Medical History|2750,2753|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Finding|Gene or Genome|Family Medical History|2750,2753|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Finding|Intellectual Product|Family Medical History|2750,2753|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Anatomy|Body System|Family Medical History|2758,2762|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|Family Medical History|2758,2762|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|Family Medical History|2758,2762|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|Family Medical History|2758,2762|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|Family Medical History|2758,2762|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Sign or Symptom|Family Medical History|2778,2784|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2791,2796|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Anatomy|Body System|Family Medical History|2798,2801|false|false|false|C3714787|Central Nervous System|CNs
Finding|Finding|Family Medical History|2809,2815|false|false|false|C1554187|Gender Status - Intact|intact
Lab|Laboratory or Test Result|Family Medical History|2837,2841|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Family Medical History|2855,2860|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|2855,2860|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2861,2864|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2869,2872|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2869,2872|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2869,2872|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2878,2881|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2878,2881|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2878,2881|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2878,2881|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2887,2890|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2887,2890|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2896,2899|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Family Medical History|2896,2899|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2896,2899|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2896,2899|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2904,2907|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2904,2907|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Family Medical History|2904,2907|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2904,2907|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2904,2907|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|2913,2917|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|2932,2935|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2952,2957|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|2952,2957|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2958,2961|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2967,2970|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2967,2970|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2967,2970|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2977,2980|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2977,2980|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2977,2980|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2977,2980|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2986,2989|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2986,2989|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2997,3000|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Family Medical History|2997,3000|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2997,3000|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2997,3000|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3004,3007|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3004,3007|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Family Medical History|3004,3007|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3004,3007|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3004,3007|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|3013,3017|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Family Medical History|3033,3036|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|3053,3058|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3053,3058|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3053,3066|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3053,3066|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3053,3066|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3059,3066|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3059,3066|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3059,3066|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Family Medical History|3059,3066|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3059,3066|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3111,3115|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3111,3115|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3111,3115|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|3137,3142|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Family Medical History|3137,3142|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|3137,3150|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|3137,3150|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|3137,3150|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|3143,3150|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|3143,3150|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|3143,3150|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Family Medical History|3143,3150|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|3143,3150|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|3193,3197|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|3193,3197|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|3193,3197|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Conceptual Entity|Family Medical History|3212,3217|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Finding|Intellectual Product|Family Medical History|3212,3217|false|false|false|C3811161;C4049106|Micro (prefix);Microbiology - Laboratory Class|MICRO
Procedure|Laboratory Procedure|Family Medical History|3212,3217|false|false|false|C0085672|Microbiology procedure|MICRO
Finding|Idea or Concept|Family Medical History|3225,3230|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|Family Medical History|3225,3237|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|Family Medical History|3231,3237|false|false|false|C4255046||REPORT
Finding|Intellectual Product|Family Medical History|3231,3237|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|Family Medical History|3231,3237|false|false|false|C0700287|Reporting|REPORT
Finding|Intellectual Product|Family Medical History|3246,3252|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|DIRECT
Disorder|Disease or Syndrome|Family Medical History|3253,3262|false|false|false|C0021400|Influenza|INFLUENZA
Drug|Immunologic Factor|Family Medical History|3253,3262|false|false|false|C0021403|Influenza virus vaccine|INFLUENZA
Drug|Pharmacologic Substance|Family Medical History|3253,3262|false|false|false|C0021403|Influenza virus vaccine|INFLUENZA
Disorder|Disease or Syndrome|Family Medical History|3253,3264|false|false|false|C2062441|influenza A|INFLUENZA A
Drug|Immunologic Factor|Family Medical History|3263,3272|false|false|false|C0348042|Blood group antigen A|A ANTIGEN
Drug|Immunologic Factor|Family Medical History|3265,3272|false|false|false|C0003320|Antigens|ANTIGEN
Procedure|Laboratory Procedure|Family Medical History|3265,3277|false|false|false|C0729856|Antigen test|ANTIGEN TEST
Anatomy|Body Location or Region|Family Medical History|3273,3277|false|false|false|C4318744|Test - temporal region|TEST
Finding|Functional Concept|Family Medical History|3273,3277|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Finding|Intellectual Product|Family Medical History|3273,3277|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TEST
Lab|Laboratory or Test Result|Family Medical History|3273,3277|false|false|false|C0456984|Test Result|TEST
Procedure|Laboratory Procedure|Family Medical History|3273,3277|false|false|false|C0022885|Laboratory Procedures|TEST
Finding|Idea or Concept|Family Medical History|3279,3284|false|false|false|C1546485|Diagnosis Type - Final|Final
Disorder|Cell or Molecular Dysfunction|Family Medical History|3297,3305|false|false|false|C4727483|BRAF Gene Rearrangement|POSITIVE
Finding|Classification|Family Medical History|3297,3305|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|Family Medical History|3297,3305|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|POSITIVE
Finding|Finding|Family Medical History|3297,3309|false|false|false|C1446409|Positive|POSITIVE FOR
Disorder|Disease or Syndrome|Family Medical History|3310,3319|false|false|false|C0021400|Influenza|INFLUENZA
Drug|Immunologic Factor|Family Medical History|3310,3319|false|false|false|C0021403|Influenza virus vaccine|INFLUENZA
Drug|Pharmacologic Substance|Family Medical History|3310,3319|false|false|false|C0021403|Influenza virus vaccine|INFLUENZA
Disorder|Disease or Syndrome|Family Medical History|3310,3321|false|false|false|C2062441|influenza A|INFLUENZA A
Finding|Functional Concept|Family Medical History|3322,3327|false|false|false|C0521026|Viral|VIRAL
Drug|Immunologic Factor|Family Medical History|3322,3335|false|false|false|C0003342|Antigens, Viral|VIRAL ANTIGEN
Drug|Immunologic Factor|Family Medical History|3328,3335|false|false|false|C0003320|Antigens|ANTIGEN
Finding|Idea or Concept|Family Medical History|3359,3364|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|PHONE
Finding|Intellectual Product|Family Medical History|3359,3364|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|PHONE
Finding|Finding|Family Medical History|3388,3395|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|Family Medical History|3388,3395|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Procedure|Diagnostic Procedure|Family Medical History|3397,3400|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Impression|3425,3430|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|3431,3436|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|3431,3436|false|false|false|C0741025|Chest problem|chest
Disorder|Disease or Syndrome|Impression|3431,3446|true|false|false|C0742323|CHEST PATHOLOGY|chest pathology
Finding|Functional Concept|Impression|3437,3446|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Impression|3437,3446|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Impression|3437,3446|false|false|false|C0919386|Pathology procedure|pathology
Finding|Intellectual Product|Impression|3452,3458|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Tissue|Impression|3459,3466|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|Impression|3459,3466|false|false|false|C0032226|Pleural Diseases|pleural
Finding|Finding|Impression|3480,3484|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Gene or Genome|Impression|3480,3484|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Pathologic Function|Impression|3480,3484|false|false|false|C0241158;C1419736;C2004491|Cicatrix;RPS4X gene;Scar Tissue|scar
Finding|Functional Concept|Impression|3490,3500|false|false|false|C0016203|Flattened|Flattening
Anatomy|Body Part, Organ, or Organ Component|Impression|3508,3522|false|false|false|C1269845|Structure of hemidiaphragm|hemidiaphragms
Finding|Idea or Concept|Impression|3523,3533|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|3523,3538|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Impression|3539,3543|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Impression|3539,3543|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Impression|3539,3543|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|Hospital Course|3581,3585|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|3581,3585|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Sign or Symptom|Hospital Course|3617,3623|false|false|false|C0015967|Fever|fevers
Drug|Organic Chemical|Hospital Course|3637,3642|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|3637,3642|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|3637,3642|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|Hospital Course|3665,3679|false|false|false|C0008033|Pleuritic pain|pleuritic pain
Attribute|Clinical Attribute|Hospital Course|3675,3679|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3675,3679|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3675,3679|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Cell or Molecular Dysfunction|Hospital Course|3691,3699|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|3691,3699|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|3691,3699|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|Hospital Course|3705,3714|false|false|false|C0021400|Influenza|influenza
Drug|Immunologic Factor|Hospital Course|3705,3714|false|false|false|C0021403|Influenza virus vaccine|influenza
Drug|Pharmacologic Substance|Hospital Course|3705,3714|false|false|false|C0021403|Influenza virus vaccine|influenza
Disorder|Disease or Syndrome|Hospital Course|3705,3716|false|false|false|C2062441|influenza A|influenza A
Finding|Sign or Symptom|Hospital Course|3722,3728|false|false|false|C0015967|Fever|Fevers
Finding|Sign or Symptom|Hospital Course|3730,3737|false|false|false|C0231218|Malaise|malaise
Drug|Organic Chemical|Hospital Course|3739,3744|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|3739,3744|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|3739,3744|false|false|false|C0010200|Coughing|cough
Finding|Functional Concept|Hospital Course|3773,3781|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|3773,3781|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Idea or Concept|Hospital Course|3783,3793|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|3783,3798|false|false|false|C0332290|Consistent with|consistent with
Finding|Functional Concept|Hospital Course|3799,3804|false|false|false|C0521026|Viral|viral
Disorder|Disease or Syndrome|Hospital Course|3799,3814|false|false|false|C0042769|Virus Diseases|viral infection
Disorder|Disease or Syndrome|Hospital Course|3805,3814|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|3805,3814|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|Hospital Course|3842,3850|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3865,3884|false|false|false|C1443870|Respiratory secretion precautions|droplet precautions
Finding|Conceptual Entity|Hospital Course|3873,3884|false|false|false|C1882442|Precaution|precautions
Finding|Idea or Concept|Hospital Course|3904,3911|false|false|false|C2699424|Concern|concern
Disorder|Disease or Syndrome|Hospital Course|3929,3932|false|false|false|C0021400|Influenza|flu
Finding|Gene or Genome|Hospital Course|3929,3932|false|false|false|C3811318|ZMYND10 wt Allele|flu
Drug|Organic Chemical|Hospital Course|3967,3978|false|false|false|C0874161|oseltamivir|Oseltamivir
Drug|Pharmacologic Substance|Hospital Course|3967,3978|false|false|false|C0874161|oseltamivir|Oseltamivir
Disorder|Mental or Behavioral Dysfunction|Hospital Course|3987,3990|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3987,3990|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|3987,3990|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|3987,3990|false|false|false|C1332410|BID gene|BID
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3993,4007|false|false|false|C0027442|Nasopharynx|nasopharyngeal
Finding|Body Substance|Hospital Course|3993,4012|false|false|false|C0444192|Nasopharyngeal swab (specimen)|nasopharyngeal swab
Procedure|Laboratory Procedure|Hospital Course|3993,4012|false|false|false|C2266655;C4318939|Nasal Swab Test;nasopharyngeal swab (lab test)|nasopharyngeal swab
Drug|Biomedical or Dental Material|Hospital Course|4008,4012|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Drug|Substance|Hospital Course|4008,4012|false|false|false|C0183753;C1706069|Swab Dosage Form;Swab specimen|swab
Procedure|Diagnostic Procedure|Hospital Course|4008,4012|false|false|false|C0563454|Taking of swab|swab
Disorder|Cell or Molecular Dysfunction|Hospital Course|4017,4025|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|4017,4025|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|4017,4025|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|4017,4029|false|false|false|C1446409|Positive|positive for
Disorder|Disease or Syndrome|Hospital Course|4031,4040|false|false|false|C0021400|Influenza|influenza
Drug|Immunologic Factor|Hospital Course|4031,4040|false|false|false|C0021403|Influenza virus vaccine|influenza
Drug|Pharmacologic Substance|Hospital Course|4031,4040|false|false|false|C0021403|Influenza virus vaccine|influenza
Finding|Idea or Concept|Hospital Course|4073,4076|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4073,4076|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|4090,4101|false|false|false|C0874161|oseltamivir|oseltamivir
Drug|Pharmacologic Substance|Hospital Course|4090,4101|false|false|false|C0874161|oseltamivir|oseltamivir
Disorder|Disease or Syndrome|Hospital Course|4110,4113|false|false|false|C0021400|Influenza|flu
Finding|Gene or Genome|Hospital Course|4110,4113|false|false|false|C3811318|ZMYND10 wt Allele|flu
Finding|Classification|Hospital Course|4154,4164|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4154,4164|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Mental Process|Hospital Course|4165,4172|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|4178,4182|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4178,4182|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4178,4182|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4178,4195|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|4183,4195|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Cell or Molecular Dysfunction|Hospital Course|4208,4216|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|4208,4216|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|4208,4216|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|4208,4220|false|false|false|C1446409|Positive|positive for
Disorder|Disease or Syndrome|Hospital Course|4225,4228|false|false|false|C0021400|Influenza|flu
Finding|Gene or Genome|Hospital Course|4225,4228|false|false|false|C3811318|ZMYND10 wt Allele|flu
Disorder|Disease or Syndrome|Hospital Course|4262,4266|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|4262,4266|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|4262,4266|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|4262,4279|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Hospital Course|4267,4279|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Finding|Hospital Course|4295,4302|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|4295,4302|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Body Substance|Hospital Course|4308,4314|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|Hospital Course|4308,4314|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Organ or Tissue Function|Hospital Course|4308,4325|false|false|false|C0242104|Sputum production|sputum production
Event|Occupational Activity|Hospital Course|4315,4325|false|false|false|C0033268|production|production
Finding|Intellectual Product|Hospital Course|4315,4325|false|false|false|C1548180|Production Processing ID|production
Drug|Hormone|Hospital Course|4347,4357|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|4347,4357|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|4347,4357|false|false|false|C0032952|prednisone|prednisone
Drug|Antibiotic|Hospital Course|4374,4386|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Hospital Course|4374,4386|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|4374,4386|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4398,4403|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|4398,4403|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|4398,4403|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|4398,4403|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|4398,4403|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|4398,4403|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4404,4411|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|Hospital Course|4404,4411|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Hospital Course|4404,4411|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Daily or Recreational Activity|Hospital Course|4418,4425|false|false|false|C0035253|Rest|resting
Finding|Finding|Hospital Course|4464,4468|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4464,4468|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4464,4468|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|4472,4481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4472,4481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4472,4481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4472,4481|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|4584,4587|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4584,4587|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Antibiotic|Hospital Course|4598,4610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|4598,4610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|4598,4610|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Hormone|Hospital Course|4623,4633|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|4623,4633|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|4623,4633|false|false|false|C0032952|prednisone|prednisone
Finding|Intellectual Product|Hospital Course|4655,4659|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|4662,4666|false|false|false|C1561540|Transaction counts and value totals - week|week
Procedure|Health Care Activity|Hospital Course|4672,4677|false|false|false|C0441640||taper
Finding|Idea or Concept|Hospital Course|4697,4701|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|4697,4701|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|4697,4701|false|false|false|C1553498|home health encounter|home
Finding|Functional Concept|Hospital Course|4715,4723|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|4715,4723|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Body Substance|Hospital Course|4739,4746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4739,4746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4739,4746|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|4794,4798|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|4806,4810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4806,4810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4806,4810|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Body Substance|Hospital Course|4815,4824|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4815,4824|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4815,4824|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4815,4824|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|4862,4866|false|false|false|C5575035|Well (answer to question)|well
Finding|Classification|Hospital Course|4886,4896|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|4886,4896|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Mental Process|Hospital Course|4897,4904|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|4910,4916|false|false|false|C0004096|Asthma|ASTHMA
Finding|Sign or Symptom|Hospital Course|4926,4934|false|false|false|C0043144|Wheezing|wheezing
Disorder|Disease or Syndrome|Hospital Course|4952,4955|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4952,4955|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|4952,4955|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4952,4955|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|4952,4955|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|4952,4955|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|4952,4955|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|4952,4955|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|4952,4955|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|4952,4955|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|Hospital Course|4956,4962|false|false|false|C1549636|Address type - Office|office
Finding|Finding|Hospital Course|4973,4980|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Hospital Course|4973,4980|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|Hospital Course|5041,5045|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|5041,5045|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|Hospital Course|5048,5054|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|5048,5054|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Disorder|Disease or Syndrome|Hospital Course|5062,5068|false|true|false|C0004096|Asthma|asthma
Finding|Functional Concept|Hospital Course|5069,5077|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5069,5077|false|true|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Mental Process|Hospital Course|5081,5088|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|Hospital Course|5092,5096|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5092,5096|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Hospital Course|5092,5096|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|Hospital Course|5139,5143|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5139,5143|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5139,5143|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|Hospital Course|5175,5185|false|false|false|C2064916|nebulizers (medication)|nebulizers
Finding|Finding|Hospital Course|5237,5241|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|Hospital Course|5249,5253|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5249,5253|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5249,5253|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|5254,5265|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5254,5265|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|5254,5265|false|false|false|C4284232|Medications|medications
Attribute|Clinical Attribute|Hospital Course|5268,5279|false|false|false|C0231832|Respiratory rate|Respiratory
Finding|Body Substance|Hospital Course|5268,5279|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Functional Concept|Hospital Course|5268,5279|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Finding|Intellectual Product|Hospital Course|5268,5279|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|Respiratory
Attribute|Clinical Attribute|Hospital Course|5268,5286|false|false|false|C2598168||Respiratory status
Finding|Finding|Hospital Course|5268,5286|false|false|false|C1998827|Respiratory Status|Respiratory status
Attribute|Clinical Attribute|Hospital Course|5280,5286|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|5280,5286|false|false|false|C1546481|What subject filter - Status|status
Finding|Idea or Concept|Hospital Course|5302,5307|false|false|false|C1552828|Table Frame - above|above
Disorder|Disease or Syndrome|Hospital Course|5311,5323|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Finding|Finding|Hospital Course|5337,5349|false|false|false|C0857121|Hypertensive (finding)|hypertensive
Finding|Idea or Concept|Hospital Course|5371,5379|false|false|false|C0549178|Continuous|continue
Disorder|Disease or Syndrome|Hospital Course|5380,5384|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Finding|Intellectual Product|Hospital Course|5380,5384|false|false|false|C4284232|Medications|meds
Phenomenon|Natural Phenomenon or Process|Hospital Course|5388,5395|false|false|false|C1705970|Electrical Current|current
Disorder|Disease or Syndrome|Hospital Course|5443,5447|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|meds
Finding|Intellectual Product|Hospital Course|5443,5447|false|false|false|C4284232|Medications|meds
Finding|Classification|Hospital Course|5485,5495|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|5485,5495|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Mental Process|Hospital Course|5497,5504|false|false|false|C0542559|contextual factors|setting
Finding|Idea or Concept|Hospital Course|5544,5552|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Anatomical Structure|Hospital Course|5566,5571|false|false|false|C3714591|Floor (anatomic)|floor
Drug|Organic Chemical|Hospital Course|5587,5596|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|5587,5596|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Organic Chemical|Hospital Course|5615,5619|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Hospital Course|5615,5619|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Organic Chemical|Hospital Course|5638,5643|false|false|false|C0590690|Imdur|IMDUR
Drug|Pharmacologic Substance|Hospital Course|5638,5643|false|false|false|C0590690|Imdur|IMDUR
Disorder|Disease or Syndrome|Hospital Course|5667,5671|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Finding|Hospital Course|5683,5695|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Drug|Organic Chemical|Hospital Course|5711,5721|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|5711,5721|false|false|false|C0028978|omeprazole|omeprazole
Disorder|Disease or Syndrome|Hospital Course|5740,5743|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5740,5743|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5740,5743|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|5740,5743|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5740,5743|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5740,5743|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5740,5743|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Finding|Hospital Course|5776,5782|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Disorder|Disease or Syndrome|Hospital Course|5776,5797|false|false|false|C0856737|Single vessel disease|single vessel disease
Anatomy|Body Location or Region|Hospital Course|5783,5789|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5783,5789|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Hospital Course|5790,5797|false|false|false|C0012634|Disease|disease
Finding|Finding|Hospital Course|5808,5820|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Finding|Hospital Course|5829,5833|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|5829,5833|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|5829,5833|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Hazardous or Poisonous Substance|Hospital Course|5859,5866|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|5859,5866|false|false|false|C0728873|Monitor brand of insecticide|monitor
Finding|Functional Concept|Hospital Course|5876,5884|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5876,5884|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Procedure|Health Care Activity|Hospital Course|5897,5906|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|5922,5929|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|5922,5929|false|false|false|C0004057|aspirin|aspirin
Drug|Hazardous or Poisonous Substance|Hospital Course|5946,5953|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Hospital Course|5946,5953|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Hospital Course|5946,5953|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Hospital Course|5946,5953|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5946,5959|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5954,5959|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Hospital Course|5954,5959|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Hospital Course|5954,5959|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Functional Concept|Hospital Course|6042,6046|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Hospital Course|6042,6050|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Drug|Hazardous or Poisonous Substance|Hospital Course|6053,6061|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|Hospital Course|6053,6061|false|false|false|C0028040|nicotine|nicotine
Drug|Clinical Drug|Hospital Course|6053,6067|false|false|false|C0358855|Nicotine Transdermal Patch|nicotine patch
Drug|Biomedical or Dental Material|Hospital Course|6062,6067|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Hospital Course|6062,6067|false|false|false|C0332461|Plaque (lesion)|patch
Anatomy|Tissue|Hospital Course|6071,6074|false|false|false|C0017562|Gingiva|gum
Drug|Biomedical or Dental Material|Hospital Course|6071,6074|false|false|false|C0812395;C1378701|Gum Dose Form;Gum as an ingredient|gum
Finding|Gene or Genome|Hospital Course|6071,6074|false|false|false|C1825233;C5444202|OTULIN gene;OTULIN wt Allele|gum
Finding|Finding|Hospital Course|6084,6088|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|6084,6088|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|6084,6088|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|Hospital Course|6097,6108|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6097,6108|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|6097,6108|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|6097,6121|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|6112,6121|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6126,6136|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|6126,6136|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|6153,6162|false|false|false|C0939261|B-Complex|B complex
Drug|Pharmacologic Substance|Hospital Course|6153,6162|false|false|false|C0939261|B-Complex|B complex
Drug|Vitamin|Hospital Course|6153,6162|false|false|false|C0939261|B-Complex|B complex
Drug|Chemical Viewed Structurally|Hospital Course|6155,6162|false|false|false|C1704241|complex (molecular entity)|complex
Drug|Organic Chemical|Hospital Course|6163,6170|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|6163,6170|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|6163,6170|false|false|false|C0042890|Vitamins|vitamin
Drug|Organic Chemical|Hospital Course|6163,6172|false|false|false|C0003968;C2349136;C3714687;C4522080|Vitamin C Drug Class;Vitamin C Vitamins;Vitamin C [EPC];ascorbic acid|vitamin C
Drug|Pharmacologic Substance|Hospital Course|6163,6172|false|false|false|C0003968;C2349136;C3714687;C4522080|Vitamin C Drug Class;Vitamin C Vitamins;Vitamin C [EPC];ascorbic acid|vitamin C
Drug|Vitamin|Hospital Course|6163,6172|false|false|false|C0003968;C2349136;C3714687;C4522080|Vitamin C Drug Class;Vitamin C Vitamins;Vitamin C [EPC];ascorbic acid|vitamin C
Procedure|Laboratory Procedure|Hospital Course|6163,6172|false|false|false|C0201898|Ascorbic acid measurement|vitamin C
Drug|Organic Chemical|Hospital Course|6173,6183|false|false|false|C0016410|folic acid|folic acid
Drug|Pharmacologic Substance|Hospital Course|6173,6183|false|false|false|C0016410|folic acid|folic acid
Drug|Vitamin|Hospital Course|6173,6183|false|false|false|C0016410|folic acid|folic acid
Procedure|Laboratory Procedure|Hospital Course|6173,6183|false|false|false|C0523631|Folic acid measurement|folic acid
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6189,6196|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6189,6196|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6189,6196|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Congenital Abnormality|Hospital Course|6210,6213|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|6210,6213|false|false|false|C0006935|capsule (pharmacologic)|Cap
Finding|Gene or Genome|Hospital Course|6210,6213|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6210,6213|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Drug|Organic Chemical|Hospital Course|6240,6250|false|false|false|C1337242|cinacalcet|cinacalcet
Drug|Pharmacologic Substance|Hospital Course|6240,6250|false|false|false|C1337242|cinacalcet|cinacalcet
Drug|Biomedical or Dental Material|Hospital Course|6257,6263|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6277,6283|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6308,6319|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|6308,6319|false|false|false|C0074554|simvastatin|simvastatin
Drug|Biomedical or Dental Material|Hospital Course|6326,6332|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6346,6352|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6378,6388|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|6378,6388|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|6378,6398|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Pharmacologic Substance|Hospital Course|6378,6398|false|false|false|C0724633|metoprolol succinate|metoprolol succinate
Drug|Organic Chemical|Hospital Course|6389,6398|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Drug|Biomedical or Dental Material|Hospital Course|6406,6412|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|6423,6430|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6423,6430|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6423,6430|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|6452,6458|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|6469,6476|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6469,6476|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6469,6476|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|Hospital Course|6486,6490|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6486,6496|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6493,6496|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6493,6496|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6503,6512|false|false|false|C0114873|doxazosin|doxazosin
Drug|Pharmacologic Substance|Hospital Course|6503,6512|false|false|false|C0114873|doxazosin|doxazosin
Drug|Biomedical or Dental Material|Hospital Course|6518,6524|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6538,6544|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6571,6578|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|6571,6578|false|false|false|C0004057|aspirin|aspirin
Drug|Biomedical or Dental Material|Hospital Course|6585,6591|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6585,6601|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6602,6605|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6602,6605|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6602,6605|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6602,6605|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|6615,6621|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6615,6631|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Organic Chemical|Hospital Course|6658,6669|false|false|false|C0078569|venlafaxine|venlafaxine
Drug|Pharmacologic Substance|Hospital Course|6658,6669|false|false|false|C0078569|venlafaxine|venlafaxine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6676,6683|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6676,6683|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6676,6683|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6691,6698|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6691,6698|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6691,6698|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6720,6727|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6720,6727|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6720,6727|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6735,6742|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6735,6742|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6735,6742|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|6772,6783|false|false|false|C0078569|venlafaxine|venlafaxine
Drug|Pharmacologic Substance|Hospital Course|6772,6783|false|false|false|C0078569|venlafaxine|venlafaxine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6792,6799|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6792,6799|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6792,6799|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6807,6814|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6807,6814|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6807,6814|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6837,6844|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6837,6844|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6837,6844|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|6852,6859|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6852,6859|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6852,6859|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|6890,6899|false|false|false|C0718050|sevelamer|sevelamer
Drug|Pharmacologic Substance|Hospital Course|6890,6899|false|false|false|C0718050|sevelamer|sevelamer
Drug|Organic Chemical|Hospital Course|6890,6903|false|false|false|C0772463|sevelamer hydrochloride|sevelamer HCl
Drug|Pharmacologic Substance|Hospital Course|6890,6903|false|false|false|C0772463|sevelamer hydrochloride|sevelamer HCl
Disorder|Neoplastic Process|Hospital Course|6900,6903|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|6900,6903|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|6900,6903|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|6900,6903|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Biomedical or Dental Material|Hospital Course|6911,6917|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6931,6937|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Daily or Recreational Activity|Hospital Course|6949,6954|false|false|false|C1998602|Meal (occasion for eating)|MEALS
Finding|Finding|Hospital Course|6956,6963|false|false|false|C4035626|3 times|3 TIMES
Disorder|Disease or Syndrome|Hospital Course|6958,6963|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|TIMES
Finding|Idea or Concept|Hospital Course|6966,6969|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|6966,6969|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Daily or Recreational Activity|Hospital Course|6975,6980|false|false|false|C1998602|Meal (occasion for eating)|MEALS
Drug|Biomedical or Dental Material|Hospital Course|6995,7001|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|7006,7013|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|7024,7034|false|false|false|C0009011|clonazepam|clonazepam
Drug|Pharmacologic Substance|Hospital Course|7024,7034|false|false|false|C0009011|clonazepam|clonazepam
Drug|Biomedical or Dental Material|Hospital Course|7040,7046|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7060,7066|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Body Substance|Hospital Course|7087,7096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7087,7096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7087,7096|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7087,7096|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|7087,7108|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|7097,7108|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7097,7108|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|7097,7108|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|7113,7126|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|7113,7126|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|Hospital Course|7113,7126|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|7134,7140|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7154,7160|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|Hospital Course|7200,7204|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7200,7204|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7200,7204|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|7211,7220|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|7211,7220|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|7211,7228|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|7211,7228|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|7221,7228|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|7221,7228|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|7221,7228|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Disorder|Disease or Syndrome|Hospital Course|7246,7249|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|7246,7249|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|7250,7257|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Functional Concept|Hospital Course|7258,7265|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Hospital Course|7281,7291|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|7281,7291|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Drug|Antibiotic|Hospital Course|7314,7326|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|7314,7326|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|7314,7326|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Biomedical or Dental Material|Hospital Course|7334,7340|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7354,7360|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|7370,7375|false|false|false|C1720374|Every - dosing instruction fragment|every
Drug|Biomedical or Dental Material|Hospital Course|7407,7413|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|7418,7425|false|false|false|C0807726|refill|Refills
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7451,7458|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7451,7458|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7451,7458|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7472,7479|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7472,7479|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7472,7479|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7483,7486|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7483,7486|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|7483,7486|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|7483,7486|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|7491,7496|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|7499,7502|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7499,7502|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7524,7531|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7524,7531|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7524,7531|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|7536,7543|false|false|false|C0807726|refill|Refills
Drug|Hormone|Hospital Course|7551,7561|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|7551,7561|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|7551,7561|false|false|false|C0032952|prednisone|prednisone
Drug|Biomedical or Dental Material|Hospital Course|7568,7574|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7589,7595|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|7599,7603|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7599,7609|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7606,7609|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7606,7609|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7647,7651|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|7671,7675|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Hospital Course|7696,7700|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Biomedical or Dental Material|Hospital Course|7703,7706|false|false|false|C0039225|Tablet Dosage Form|tab
Drug|Biomedical or Dental Material|Hospital Course|7728,7734|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|7739,7746|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|7754,7763|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|7754,7763|false|false|false|C0012373|diltiazem|diltiazem
Drug|Organic Chemical|Hospital Course|7754,7767|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Hospital Course|7754,7767|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Hospital Course|7764,7767|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|7764,7767|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|7764,7767|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|7764,7767|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7775,7782|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7775,7782|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7775,7782|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7775,7800|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Hospital Course|7784,7792|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7784,7792|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7793,7800|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7793,7800|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7793,7800|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7815,7822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7815,7822|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7815,7822|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7815,7840|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Hospital Course|7824,7832|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7824,7832|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|7833,7840|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7833,7840|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7833,7840|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|7864,7875|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|7864,7875|false|false|false|C0082607|fluticasone|fluticasone
Drug|Biomedical or Dental Material|Hospital Course|7893,7898|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|7893,7898|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|7893,7898|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|7893,7910|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Hospital Course|7900,7910|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|7900,7910|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Finding|Functional Concept|Hospital Course|7900,7910|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|Hospital Course|7925,7930|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|7925,7930|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|7925,7930|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7931,7936|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|7931,7936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|7931,7936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|7931,7936|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|7931,7936|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|7931,7936|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Drug|Organic Chemical|Hospital Course|7957,7968|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|7957,7968|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|7957,7979|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|7969,7979|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|7969,7979|false|false|false|C0073992|salmeterol|salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7996,8000|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|7996,8000|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|8006,8012|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8013,8016|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8013,8016|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|8013,8016|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|8013,8016|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8027,8031|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|8027,8031|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|8037,8043|false|false|false|C1550509|Participation Type - device|Device
Finding|Functional Concept|Hospital Course|8044,8054|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|8044,8054|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8055,8058|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8055,8058|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8055,8058|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|8055,8058|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|8060,8067|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|8062,8067|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|8070,8073|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8070,8073|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|8081,8100|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|8081,8100|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8109,8116|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8109,8116|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8109,8116|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8130,8137|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8130,8137|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8130,8137|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|Hospital Course|8163,8173|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Hospital Course|8163,8173|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|Hospital Course|8163,8185|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|Hospital Course|8163,8185|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Biomedical or Dental Material|Hospital Course|8192,8198|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Hospital Course|8199,8207|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8199,8207|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8208,8215|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8208,8215|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8208,8215|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|8236,8242|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Hospital Course|8243,8251|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8243,8251|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8252,8259|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8252,8259|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8252,8259|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8290,8301|false|false|false|C0298130|montelukast|montelukast
Drug|Pharmacologic Substance|Hospital Course|8290,8301|false|false|false|C0298130|montelukast|montelukast
Drug|Biomedical or Dental Material|Hospital Course|8308,8314|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8328,8334|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|8360,8370|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|8360,8370|false|false|false|C0028978|omeprazole|omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8377,8384|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8377,8384|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8377,8384|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|8386,8393|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|8386,8401|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|Hospital Course|8394,8401|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8394,8401|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8394,8401|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8422,8429|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8422,8429|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8422,8429|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|8431,8438|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|8431,8446|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|Hospital Course|8439,8446|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8439,8446|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8439,8446|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8477,8487|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Hospital Course|8477,8487|false|false|false|C0213771|tiotropium|tiotropium
Drug|Organic Chemical|Hospital Course|8477,8495|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Hospital Course|8477,8495|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Hospital Course|8488,8495|false|false|false|C0006222|Bromides|bromide
Procedure|Laboratory Procedure|Hospital Course|8488,8495|false|false|false|C0202341|Bromides measurement|bromide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8503,8510|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|8503,8510|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|8503,8510|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|8514,8524|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|8514,8524|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Functional Concept|Hospital Course|8525,8531|false|false|false|C1550509|Participation Type - device|Device
Disorder|Congenital Abnormality|Hospital Course|8546,8549|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|8546,8549|false|false|false|C0006935|capsule (pharmacologic)|Cap
Finding|Gene or Genome|Hospital Course|8546,8549|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8546,8549|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Finding|Functional Concept|Hospital Course|8550,8560|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|8550,8560|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Drug|Biologically Active Substance|Hospital Course|8582,8589|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|8582,8589|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|8582,8589|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|8582,8589|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|8582,8589|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|Hospital Course|8582,8589|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|8582,8589|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Hospital Course|8582,8599|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Hospital Course|8582,8599|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Hospital Course|8590,8599|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Hospital Course|8590,8599|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Hospital Course|8590,8599|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Biomedical or Dental Material|Hospital Course|8616,8622|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8616,8632|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8633,8636|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8633,8636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|8633,8636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|8633,8636|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Hospital Course|8647,8653|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8647,8663|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Organic Chemical|Hospital Course|8688,8700|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|8688,8700|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|8688,8700|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|8688,8711|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|8705,8711|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8725,8731|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|8757,8764|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|8757,8764|false|false|false|C0004057|aspirin|aspirin
Drug|Biomedical or Dental Material|Hospital Course|8771,8777|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|8791,8797|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|8801,8805|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|8801,8811|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|8808,8811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|8808,8811|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biologically Active Substance|Hospital Course|8819,8825|false|false|false|C0030054|oxygen|Oxygen
Drug|Element, Ion, or Isotope|Hospital Course|8819,8825|false|false|false|C0030054|oxygen|Oxygen
Drug|Pharmacologic Substance|Hospital Course|8819,8825|false|false|false|C0030054|oxygen|Oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8819,8825|false|false|false|C0184633|Oxygen Therapy Care|Oxygen
Finding|Idea or Concept|Hospital Course|8826,8830|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8826,8830|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8826,8830|false|false|false|C1553498|home health encounter|Home
Finding|Finding|Hospital Course|8826,8837|false|false|false|C0421203|Home oxygen supply|Home Oxygen
Drug|Biologically Active Substance|Hospital Course|8831,8837|false|false|false|C0030054|oxygen|Oxygen
Drug|Element, Ion, or Isotope|Hospital Course|8831,8837|false|false|false|C0030054|oxygen|Oxygen
Drug|Pharmacologic Substance|Hospital Course|8831,8837|false|false|false|C0030054|oxygen|Oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8831,8837|false|false|false|C0184633|Oxygen Therapy Care|Oxygen
Finding|Idea or Concept|Hospital Course|8845,8855|false|false|false|C0549178|Continuous|Continuous
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8860,8865|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8860,8865|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8860,8865|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8860,8865|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8860,8865|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8860,8865|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8866,8873|false|false|false|C1550232|Body Parts - Cannula|cannula
Finding|Body Substance|Hospital Course|8866,8873|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Intellectual Product|Hospital Course|8866,8873|false|false|false|C1546577;C1550622|Specimen Type - Cannula|cannula
Finding|Functional Concept|Hospital Course|8887,8893|false|false|false|C1550509|Participation Type - device|device
Attribute|Clinical Attribute|Hospital Course|8912,8917|false|false|false|C0232117|Pulse Rate|Pulse
Finding|Physiologic Function|Hospital Course|8912,8917|false|false|false|C0391850|Physiologic pulse|Pulse
Phenomenon|Phenomenon or Process|Hospital Course|8912,8917|false|false|false|C1947910|Pulse phenomenon|Pulse
Procedure|Health Care Activity|Hospital Course|8912,8917|false|false|false|C0034107|Pulse taking|Pulse
Finding|Body Substance|Hospital Course|8943,8952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8943,8952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8943,8952|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8943,8952|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8943,8964|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8943,8964|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8953,8964|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|8953,8964|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|8966,8970|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8966,8970|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8966,8970|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|8976,8983|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|8976,8983|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|Hospital Course|8986,8994|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|9002,9011|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9002,9011|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9002,9011|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9002,9011|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9002,9021|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9012,9021|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|9012,9021|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9012,9021|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9012,9021|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|9042,9051|false|false|false|C0021400|Influenza|Influenza
Drug|Immunologic Factor|Principle Diagnosis|9042,9051|false|false|false|C0021403|Influenza virus vaccine|Influenza
Drug|Pharmacologic Substance|Principle Diagnosis|9042,9051|false|false|false|C0021403|Influenza virus vaccine|Influenza
Disorder|Disease or Syndrome|Principle Diagnosis|9052,9056|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Principle Diagnosis|9052,9056|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Principle Diagnosis|9052,9056|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Principle Diagnosis|9052,9069|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Principle Diagnosis|9057,9069|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Neoplastic Process|Principle Diagnosis|9072,9081|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Principle Diagnosis|9072,9081|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Principle Diagnosis|9072,9091|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|Principle Diagnosis|9072,9091|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|Principle Diagnosis|9082,9091|false|false|false|C0945731||Diagnosis
Finding|Classification|Principle Diagnosis|9082,9091|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Principle Diagnosis|9082,9091|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Principle Diagnosis|9082,9091|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Principle Diagnosis|9093,9099|false|false|false|C0004096|Asthma|ASTHMA
Disorder|Disease or Syndrome|Principle Diagnosis|9103,9115|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Disorder|Disease or Syndrome|Principle Diagnosis|9119,9133|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Finding|Finding|Principle Diagnosis|9119,9133|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Finding|Sign or Symptom|Principle Diagnosis|9137,9145|false|false|false|C0018681|Headache|HEADACHE
Disorder|Disease or Syndrome|Principle Diagnosis|9149,9163|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Finding|Finding|Principle Diagnosis|9167,9175|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Principle Diagnosis|9167,9186|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Principle Diagnosis|9176,9181|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Principle Diagnosis|9176,9181|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Principle Diagnosis|9176,9186|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Principle Diagnosis|9176,9186|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Principle Diagnosis|9182,9186|false|true|false|C2598155||PAIN
Finding|Functional Concept|Principle Diagnosis|9182,9186|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Principle Diagnosis|9182,9186|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Drug|Hazardous or Poisonous Substance|Principle Diagnosis|9190,9197|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Principle Diagnosis|9190,9197|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Principle Diagnosis|9190,9197|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Principle Diagnosis|9190,9197|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Principle Diagnosis|9190,9203|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Principle Diagnosis|9198,9203|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Principle Diagnosis|9198,9203|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Principle Diagnosis|9198,9203|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Finding|Principle Diagnosis|9207,9215|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Idea or Concept|Principle Diagnosis|9207,9215|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Finding|Principle Diagnosis|9207,9221|false|false|false|C0742257|chest abnormal|ABNORMAL CHEST
Finding|Finding|Principle Diagnosis|9207,9226|false|false|false|C0436503|Standard chest X-ray abnormal|ABNORMAL CHEST XRAY
Anatomy|Body Location or Region|Principle Diagnosis|9216,9221|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Principle Diagnosis|9216,9221|false|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|Principle Diagnosis|9216,9226|false|false|false|C0039985|Plain chest X-ray|CHEST XRAY
Phenomenon|Natural Phenomenon or Process|Principle Diagnosis|9222,9226|false|false|false|C0043309|Roentgen Rays|XRAY
Procedure|Diagnostic Procedure|Principle Diagnosis|9222,9226|false|false|false|C0043299|Diagnostic radiologic examination|XRAY
Disorder|Disease or Syndrome|Principle Diagnosis|9230,9234|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Principle Diagnosis|9230,9234|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Principle Diagnosis|9230,9234|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Mental Process|Discharge Condition|9260,9266|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9260,9273|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9260,9273|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9267,9273|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9267,9273|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|9275,9280|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|9285,9293|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|9295,9317|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9295,9317|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|9304,9317|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9304,9317|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9319,9324|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9319,9324|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9319,9324|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|9319,9324|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9319,9324|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9319,9324|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9329,9340|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9342,9350|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9342,9350|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9342,9350|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9351,9357|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9351,9357|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|9359,9369|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9359,9369|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9359,9369|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9359,9369|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|9372,9383|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|9372,9383|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Intellectual Product|Discharge Instructions|9458,9466|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9458,9466|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|9474,9478|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|9474,9478|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9474,9478|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9474,9481|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|Discharge Instructions|9514,9522|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Functional Concept|Discharge Instructions|9527,9535|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|9527,9535|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Functional Concept|Discharge Instructions|9559,9565|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Discharge Instructions|9559,9565|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Disorder|Disease or Syndrome|Discharge Instructions|9559,9570|false|false|false|C0009443|Common Cold|common cold
Disorder|Disease or Syndrome|Discharge Instructions|9566,9570|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|Discharge Instructions|9566,9570|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|Discharge Instructions|9566,9570|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Finding|Organism Function|Discharge Instructions|9566,9570|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|9566,9570|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9566,9570|false|false|false|C0010412|Cold Therapy|cold
Finding|Finding|Discharge Instructions|9574,9578|false|false|false|C5575035|Well (answer to question)|well
Finding|Idea or Concept|Discharge Instructions|9583,9592|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Attribute|Clinical Attribute|Discharge Instructions|9593,9604|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|Discharge Instructions|9593,9604|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|Discharge Instructions|9593,9604|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|Discharge Instructions|9593,9604|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Attribute|Clinical Attribute|Discharge Instructions|9593,9611|false|false|false|C2598168||respiratory status
Finding|Finding|Discharge Instructions|9593,9611|false|false|false|C1998827|Respiratory Status|respiratory status
Attribute|Clinical Attribute|Discharge Instructions|9605,9611|false|false|false|C5889824||status
Finding|Idea or Concept|Discharge Instructions|9605,9611|false|false|false|C1546481|What subject filter - Status|status
Disorder|Cell or Molecular Dysfunction|Discharge Instructions|9625,9633|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Discharge Instructions|9625,9633|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Discharge Instructions|9625,9633|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Discharge Instructions|9625,9637|false|false|false|C1446409|Positive|positive for
Disorder|Disease or Syndrome|Discharge Instructions|9643,9646|false|false|false|C0021400|Influenza|flu
Finding|Gene or Genome|Discharge Instructions|9643,9646|false|false|false|C3811318|ZMYND10 wt Allele|flu
Disorder|Disease or Syndrome|Discharge Instructions|9689,9693|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|9689,9693|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Discharge Instructions|9689,9693|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Discharge Instructions|9689,9706|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Finding|Finding|Discharge Instructions|9694,9706|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Finding|Discharge Instructions|9730,9734|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Discharge Instructions|9730,9734|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Discharge Instructions|9730,9734|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Organic Chemical|Discharge Instructions|9740,9748|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Discharge Instructions|9740,9748|false|false|false|C0038317|Steroids|steroids
Drug|Antibiotic|Discharge Instructions|9750,9762|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Discharge Instructions|9750,9762|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Discharge Instructions|9750,9762|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Discharge Instructions|9764,9771|false|false|false|C0876173|Tamiflu|tamiflu
Drug|Pharmacologic Substance|Discharge Instructions|9764,9771|false|false|false|C0876173|Tamiflu|tamiflu
Drug|Pharmacologic Substance|Discharge Instructions|9777,9787|false|false|false|C2064916|nebulizers (medication)|nebulizers
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9811,9820|false|false|false|C0184633|Oxygen Therapy Care|on oxygen
Drug|Biologically Active Substance|Discharge Instructions|9814,9820|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|9814,9820|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|9814,9820|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9814,9820|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Finding|Idea or Concept|Discharge Instructions|9842,9848|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Finding|Discharge Instructions|9869,9876|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|9872,9876|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|9872,9876|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|9872,9876|false|false|false|C1553498|home health encounter|home
Finding|Finding|Discharge Instructions|9886,9890|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|9886,9890|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|9886,9890|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|Discharge Instructions|9900,9909|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Discharge Instructions|9900,9909|false|false|false|C3714514|Infection|infection
Finding|Pathologic Function|Discharge Instructions|9928,9940|false|false|false|C0021368|Inflammation|inflammation
Attribute|Clinical Attribute|Discharge Instructions|9967,9978|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9967,9978|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|9967,9978|false|false|false|C4284232|Medications|medications
Drug|Hormone|Discharge Instructions|9993,10003|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Discharge Instructions|9993,10003|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Discharge Instructions|9993,10003|false|false|false|C0032952|prednisone|Prednisone
Finding|Idea or Concept|Discharge Instructions|10011,10014|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|10011,10014|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|10136,10140|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|Discharge Instructions|10136,10145|false|false|false|C1720393|Then stop|then stop
Drug|Antibiotic|Discharge Instructions|10148,10160|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Discharge Instructions|10148,10160|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Discharge Instructions|10148,10160|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Finding|Functional Concept|Discharge Instructions|10167,10175|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Discharge Instructions|10170,10175|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|10170,10175|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Idea or Concept|Discharge Instructions|10184,10187|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|10184,10187|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Discharge Instructions|10206,10213|false|false|false|C0876173|Tamiflu|Tamiflu
Drug|Pharmacologic Substance|Discharge Instructions|10206,10213|false|false|false|C0876173|Tamiflu|Tamiflu
Disorder|Disease or Syndrome|Discharge Instructions|10223,10228|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Discharge Instructions|10231,10234|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|10231,10234|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Discharge Instructions|10291,10295|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|10291,10295|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|10291,10295|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|10324,10335|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|10324,10335|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|10324,10335|false|false|false|C4284232|Medications|medications
Procedure|Health Care Activity|Discharge Instructions|10353,10361|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10362,10374|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|10362,10374|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

