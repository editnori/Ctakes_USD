CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Known|Modifier|false|false||Knownnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Adverse reaction to drug|Finding|true|false||Adverse Drug Reactionsnull|Adverse reaction to drug|Finding|true|false||Drug Reactionsnull|Pharmaceutical Preparations|Drug|false|false||Drug
null|Pharmacologic Substance|Drug|false|false||Drugnull|Drug problem|Finding|false|false||Drugnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Epistaxis|Finding|false|false||Epistaxisnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C0016658;C1272939;C0721966;C4520890;C1522019|nasalnull|Fracture|Disorder|false|false|C0028429|fracturesnull|Fractured|Finding|false|false||fracturesnull|Epistaxis|Finding|false|false||epistaxisnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Early|Time|false|false||earliernull|Afternoon (qualifier value)|Time|false|false||afternoonnull|Curb|Disorder|false|false||curbnull|Physical trauma|Disorder|false|false|C0015450;C4266571|trauma
null|Traumatic injury|Disorder|false|false|C0015450;C4266571|trauma
null|Trauma|Disorder|false|false|C0015450;C4266571|traumanull|Trauma assessment and care|Procedure|false|false|C0015450;C4266571|traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C3714660;C3263723;C1368081;C0548346|face
null|Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C3714660;C3263723;C1368081;C0548346|facenull|Face (spatial concept)|Modifier|false|false||facenull|Loss (adaptation)|Finding|true|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Consciousness related finding|Finding|false|false||consciousness
null|Conscious|Finding|false|false||consciousness
null|null|Finding|false|false||consciousnessnull|Persistent|Time|false|false||persistentnull|Physical trauma|Disorder|false|false|C0015450;C4266571|trauma
null|Traumatic injury|Disorder|false|false|C0015450;C4266571|trauma
null|Trauma|Disorder|false|false|C0015450;C4266571|traumanull|Trauma assessment and care|Procedure|false|false|C0015450;C4266571|traumanull|Trauma, nursing specialty|Title|false|false||traumanull|trauma qualifier|Modifier|false|false||traumanull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C1423759;C2828055;C1414531;C3160739;C3714660;C3263723;C1368081;C0548346|face
null|Face|Anatomy|false|false|C1423759;C2828055;C1414531;C3160739;C3714660;C3263723;C1368081;C0548346|facenull|Face (spatial concept)|Modifier|false|false||facenull|Further|Modifier|false|false||furthernull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C1423759;C2828055;C1414531;C0812434;C0684335;C0876917;C0362076;C3160739|head
null|Head|Anatomy|false|false|C1423759;C2828055;C1414531;C0812434;C0684335;C0876917;C0362076;C3160739|headnull|Head Device|Device|false|false||headnull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206;C0018670;C0152336|neck
null|Neck problem|Finding|false|false|C0027530;C3159206;C0018670;C0152336|necknull|dendritic spine neck|Anatomy|false|false|C3160739;C0812434;C0684335;C1423759;C2828055;C1414531|neck
null|Neck|Anatomy|false|false|C3160739;C0812434;C0684335;C1423759;C2828055;C1414531|necknull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0027530;C3159206;C0015450;C4266571;C0018670;C0152336|facenull|FANCE wt Allele|Finding|false|false|C0018670;C0152336;C0027530;C3159206;C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0018670;C0152336;C0027530;C3159206;C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0018670;C0152336;C0027530;C3159206;C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531|face
null|Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531|facenull|Face (spatial concept)|Modifier|false|false||facenull|Nasal bone structure|Anatomy|false|false|C4520890;C1522019;C1546560;C1550616|nasal bonenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0027422;C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0027422;C0028429|nasalnull|null|Anatomy|false|false|C1272939;C0721966;C4520890;C1522019|nasalnull|Specimen Type - Bone|Finding|false|false|C0027422;C1442209;C0262950|bone
null|null|Finding|false|false|C0027422;C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|Septal|Modifier|false|false||septalnull|Fracture|Disorder|false|false||fracturenull|Persistent|Time|false|false||persistentnull|Epistaxis|Finding|false|false||epistaxisnull|Bilateral|Modifier|false|false||bilateralnull|Small|LabModifier|false|false||smallnull|Abrasion Pharmacologic Substance|Drug|false|false||abrasionnull|Superficial abrasion|Disorder|false|false||abrasion
null|Abrasion|Disorder|false|false||abrasion
null|skin abrasion|Disorder|false|false||abrasionnull|Surgical abrasion|Procedure|false|false||abrasionnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Hemorrhage|Finding|false|false||Bleedingnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Lightheadedness|Finding|false|false||lightheadednull|Hypotensive|Finding|false|false||hypotensivenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Brief loss of consciousness|Disorder|false|false||brief loss of consciousnessnull|Behavior Rating Inventory of Executive Function|Finding|false|false||brief
null|BRIEF Health Literacy Screening Tool|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Unconscious State|Finding|false|false||loss of consciousnessnull|Loss (adaptation)|Finding|false|false||lossnull|Loss (quantitative)|LabModifier|false|false||lossnull|Consciousness related finding|Finding|false|false||consciousness
null|Conscious|Finding|false|false||consciousness
null|null|Finding|false|false||consciousnessnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Eye|Anatomy|false|false|C5848506|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Problems with head|Disorder|false|false|C0018670;C0152336|headnull|Procedure on head|Procedure|false|false|C0018670;C0152336|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0876917;C0362076|head
null|Head|Anatomy|false|false|C0876917;C0362076|headnull|Head Device|Device|false|false||headnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Event|Event|false|false||eventnull|Confusion|Disorder|false|false||confusionnull|Clouded consciousness|Finding|false|false||confusionnull|Further|Modifier|false|false||furthernull|Episode of|Time|false|false||episodesnull|Syncope|Finding|true|false||syncopenull|Syncope <Gastrophryninae>|Entity|true|false||syncopenull|Hemodynamics|Finding|false|false||hemodynamicnull|hemodynamics (procedure)|Procedure|false|false||hemodynamicnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Event|Event|false|false||eventnull|Epistaxis|Finding|false|false||epistaxisnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Further|Modifier|false|false||furthernull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Laboratory test finding|Lab|false|false||Labsnull|Leukocytes|Anatomy|false|false||WBCnull|Primed lymphocyte test|Procedure|false|false||pltnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false||BUNnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Urinalysis; qualitative or semiquantitative, except immunoassays|Procedure|false|false||urinalysis
null|Urinalysis|Procedure|false|false||urinalysisnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Plain chest X-ray|Procedure|false|false||CXRnull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Basal segment of lung|Anatomy|false|false|C1720922;C0740941;C1549548;C1705938;C1843354;C0024115;C0220787;C2712334;C0700198;C0332149;C0349707|lung basenull|Lung diseases|Disorder|false|false|C2987514;C0225704;C4037972;C0024109|lungnull|Lung Problem|Finding|false|false|C0225704;C2987514;C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0740941;C0024115|lung
null|Lung|Anatomy|false|false|C1549548;C1705938;C1843354;C0740941;C0024115|lungnull|nitrogenous base|Drug|false|false|C2987514|base
null|Base|Drug|false|false|C2987514|base
null|Dental Base|Drug|false|false|C2987514|base
null|base - RoleClass|Drug|false|false|C2987514|basenull|Base - General Qualifier|Finding|false|false|C2987514;C0225704;C4037972;C0024109|base
null|BPIFA4P gene|Finding|false|false|C2987514;C0225704;C4037972;C0024109|base
null|Base - RX Component Type|Finding|false|false|C2987514;C0225704;C4037972;C0024109|basenull|Anatomical base|Anatomy|false|false|C1549548;C1705938;C1843354;C0024115;C0740941;C0220787;C2712334;C0700198;C0349707;C0332149;C1720922;C1704464;C0178499;C1550601;C1880279|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Possible|Finding|false|false|C0225704;C2987514|possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Respiratory Aspiration|Disorder|false|false|C0225704;C2987514|aspirationnull|Aspiration into respiratory tract|Finding|false|false|C2987514;C0225704|aspiration
null|Endotracheal aspiration|Finding|false|false|C2987514;C0225704|aspiration
null|Pulmonary aspiration|Finding|false|false|C2987514;C0225704|aspirationnull|null|Procedure|false|false|C2987514;C0225704|aspirationnull|Pneumonia|Disorder|false|false||pneumonianull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Drug|false|false||Tdap
null|diphtheria, tetanus toxoids and acellular pertussis vaccine|Drug|false|false||Tdap
null|diphtheria, tetanus toxoids and acellular pertussis vaccine|Drug|false|false||Tdap
null|tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Drug|false|false||Tdapnull|amoxicillin / clavulanate|Drug|false|false||amoxicillin-clavulanatenull|amoxicillin|Drug|false|false||amoxicillin
null|amoxicillin|Drug|false|false||amoxicillinnull|clavulanate|Drug|false|false||clavulanate
null|clavulanate|Drug|false|false||clavulanatenull|Antibiotic Prophylaxis|Procedure|false|false||antibiotic prophylaxisnull|Antibiotics|Drug|false|false||antibioticnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|ondansetron|Drug|false|false||ondansetron
null|ondansetron|Drug|false|false||ondansetronnull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Hypertensive disease|Disorder|false|false||HTNnull|Hypercholesterolemia|Disorder|false|false||Hypercholesterolemianull|Hypercholesterolemia result|Finding|false|false||Hypercholesterolemianull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|unaware|Procedure|false|false||unawarenull|Family Medical History|Finding|false|false||family history ofnull|Family Medical History|Finding|false|false||family historynull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Blood Coagulation Disorders|Disorder|false|false||bleeding diathesisnull|Bleeding tendency|Finding|false|false||bleeding diathesisnull|Hemorrhage|Finding|false|false||bleedingnull|Disease susceptibility|Attribute|false|false||diathesisnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C0009938;C2136686;C1550016|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Contusions|Disorder|false|false|C0521367|bruisingnull|reported bruising (history)|Finding|false|false|C0521367|bruisingnull|Structure of both eyes|Anatomy|false|false|C0038999;C0684239;C0234233;C1547225;C0240577|both eyesnull|Eye|Anatomy|false|false|C0684239;C0234233;C0240577;C0038999;C5848506;C1547225|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Swollen nose|Finding|false|false|C0015392;C0229118|swollen nosenull|Swelling|Finding|false|false|C0229118;C0015392|swollennull|Mild Severity of Illness Code|Finding|false|false|C0229118;C0015392|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Emotional tenderness|Finding|false|false|C0015392;C0229118|tenderness
null|Sore to touch|Finding|false|false|C0015392;C0229118|tendernessnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|true|false||LADnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||RESPnull|Respiratory rate|Attribute|false|false||RESPnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKIN
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKINnull|Excoriation|Disorder|true|false||excoriationsnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Oropharyngeal|Anatomy|false|false|C1550016;C2136686;C0009938|oropharynxnull|Remote control command - Clear|Finding|false|false|C0521367|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Contusions|Disorder|false|false|C0521367|bruisingnull|reported bruising (history)|Finding|false|false|C0521367|bruisingnull|Structure of both eyes|Anatomy|false|false|C0684239;C0234233;C0240577;C0038999;C1547225|both eyesnull|Eye|Anatomy|false|false|C0684239;C0234233;C5848506;C0038999;C0240577;C1547225|eyesnull|null|Attribute|false|false|C0015392|eyesnull|Swollen nose|Finding|false|false|C0229118;C0015392|swollen nosenull|Swelling|Finding|false|false|C0015392;C0229118|swollennull|Mild Severity of Illness Code|Finding|false|false|C0229118;C0015392|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Emotional tenderness|Finding|false|false|C0229118;C0015392|tenderness
null|Sore to touch|Finding|false|false|C0229118;C0015392|tendernessnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|NECK
null|Neck problem|Finding|false|false|C0027530;C3159206|NECKnull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|NECK
null|Neck|Anatomy|false|false|C0812434;C0684335|NECKnull|Supple|Finding|false|false||Supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||RESPnull|Respiratory rate|Attribute|false|false||RESPnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|ABDnull|ABD (body structure)|Anatomy|false|false|C3811055|ABD
null|Abdomen|Anatomy|false|false|C3811055|ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Hereditary Multiple Exostoses|Disorder|false|false||EXTnull|EXT1 wt Allele|Finding|false|false||EXT
null|EXT1 gene|Finding|false|false||EXTnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|SKINnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|SKIN
null|Skin Specimen|Finding|false|false|C1123023;C4520765|SKINnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKIN
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|SKINnull|Excoriation|Disorder|true|false||excoriationsnull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Maxillary left second molar mesial prosthesis|Device|false|false||15PMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Maxillary left second molar mesial prosthesis|Device|false|false||15PMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Maxillary left second molar mesial prosthesis|Device|false|false||15PMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Cardiac markers|Procedure|false|false|C0018787|CARDIAC MARKERnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974;C1271630;C4554533|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Marker|Modifier|false|false||MARKERnull|null|Attribute|false|false|C0018787|TRENDnull|trend|Time|false|false||TRENDnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 5|Drug|false|false||MB-5null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|MB 2|Drug|false|false||MB-2null|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Plain chest X-ray|Procedure|false|false||CXRnull|Lateral|Modifier|false|false||lateralnull|View|Modifier|false|false||viewsnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|Lung|Anatomy|false|false||lungsnull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|false|false|C2987514;C0225732;C0225704;C4037972;C0024109;C0225730|consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Structure of base of left lung|Anatomy|false|false|C1552822;C0740941;C0024115;C0521530;C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279|left lung basenull|Left lung|Anatomy|false|false|C0024115;C1552822;C0740941;C1549548;C1705938;C1843354;C0521530|left lungnull|Table Cell Horizontal Align - left|Finding|false|false|C4037972;C0024109;C0225732;C0225730;C0225704|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Basal segment of lung|Anatomy|false|false|C0521530;C1549548;C1705938;C1843354;C0740941;C1552822;C1704464;C0178499;C1550601;C1880279;C0024115|lung basenull|Lung diseases|Disorder|false|false|C0225730;C0225732;C4037972;C0024109;C2987514;C0225704|lungnull|Lung Problem|Finding|false|false|C0225732;C4037972;C0024109;C0225704;C0225730;C2987514|lungnull|Chest>Lung|Anatomy|false|false|C1552822;C0740941;C0024115;C1549548;C1705938;C1843354;C0521530|lung
null|Lung|Anatomy|false|false|C1552822;C0740941;C0024115;C1549548;C1705938;C1843354;C0521530|lungnull|nitrogenous base|Drug|false|false|C2987514;C0225704;C0225732|base
null|Base|Drug|false|false|C2987514;C0225704;C0225732|base
null|Dental Base|Drug|false|false|C2987514;C0225704;C0225732|base
null|base - RoleClass|Drug|false|false|C2987514;C0225704;C0225732|basenull|Base - General Qualifier|Finding|false|false|C0225732;C2987514;C0225704;C4037972;C0024109;C0225730|base
null|BPIFA4P gene|Finding|false|false|C0225732;C2987514;C0225704;C4037972;C0024109;C0225730|base
null|Base - RX Component Type|Finding|false|false|C0225732;C2987514;C0225704;C4037972;C0024109;C0225730|basenull|Anatomical base|Anatomy|false|false|C0521530;C1704464;C0178499;C1550601;C1880279;C1549548;C1705938;C1843354;C0024115;C0740941|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Adjacent|Modifier|false|false||adjacent tonull|Adjacent|Modifier|false|false||adjacentnull|Lateral|Modifier|false|false||lateralnull|Structure of hemidiaphragm|Anatomy|false|false||hemidiaphragmnull|Mild Severity of Illness Code|Finding|false|false|C0005847|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Blood Vessel|Anatomy|false|false|C1547225|vascularnull|Vascular|Modifier|false|false||vascularnull|Hyperemia|Disorder|false|false||engorgementnull|Tick Engorgement|Finding|false|false||engorgementnull|Bilateral|Modifier|false|false||bilateralnull|Apical pulmonary opacity|Finding|false|false|C0032225|apical pleural thickeningnull|Apical|Modifier|false|false||apicalnull|Thickening of pleura|Disorder|false|false|C0032225|pleural thickeningnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0032226;C5139173;C0205400;C0264545|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Thickened|Finding|false|false|C0032225|thickeningnull|Aortic arch malformation|Disorder|false|false|C0003483;C0003489;C4037976;C0003741;C0230467;C0741204|aortic archnull|Aortic arch structure|Anatomy|false|false|C4759703;C4722404;C1538146|aortic arch
null|Chest>Aortic arch|Anatomy|false|false|C4759703;C4722404;C1538146|aortic archnull|Aorta|Anatomy|false|false|C4759703;C4722404;C1538146|aorticnull|Age-Related Clonal Hematopoiesis|Finding|false|false|C0003741;C0230467;C0741204;C0003489;C4037976;C0003483|arch
null|ZBTB8OS gene|Finding|false|false|C0003741;C0230467;C0741204;C0003489;C4037976;C0003483|archnull|Arch of foot|Anatomy|false|false|C4722404;C1538146;C4759703|arch
null|Structure of nucleus infundibularis hypothalami|Anatomy|false|false|C4722404;C1538146;C4759703|arch
null|ARCH|Anatomy|false|false|C4722404;C1538146;C4759703|archnull|Pathologic calcification, calcified structure|Finding|false|false||calcifications
null|Physiologic calcification|Finding|false|false||calcificationsnull|Calcified (qualifier value)|Modifier|false|false||calcificationsnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|ECHO protocol|Procedure|false|false||ECHO
null|Extension for Community Healthcare Outcomes|Procedure|false|false||ECHOnull|Echo <Calopterygidae>|Entity|false|false||ECHOnull|Left atrial structure|Anatomy|false|false|C1552822|left atriumnull|Table Cell Horizontal Align - left|Finding|false|false|C0018792;C0225860|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Atrium|Anatomy|false|false|C1552822|atriumnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Wall of left ventricle|Anatomy|false|false|C1552822|Left ventricular wallnull|Table Cell Horizontal Align - left|Finding|false|false|C0507618;C0504053|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Wall of ventricle|Anatomy|false|false|C1552822|ventricular wallnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Walls of a building|Device|false|false||wallnull|Dental caries|Disorder|false|false|C0333343|cavity
null|Cavitation|Disorder|false|false|C0333343|cavitynull|Body cavities|Anatomy|false|false|C1510420;C0011334|cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Left ventricular systolic dysfunction|Disorder|false|false|C0018827|left ventricular systolic dysfunctionnull|Table Cell Horizontal Align - left|Finding|false|false|C0018827|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false|C1552822;C0039155;C3887505;C1277187;C0749225;C0031847;C0277785;C3887504|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Systolic dysfunction|Finding|false|false|C0018827|systolic dysfunctionnull|Systole|Finding|false|false|C0018827|systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false|C0018827|dysfunctionnull|Dysfunction|Finding|false|false|C0018827|dysfunction
null|physiopathological|Finding|false|false|C0018827|dysfunction
null|Functional disorder|Finding|false|false|C0018827|dysfunctionnull|Focal|Modifier|false|false||focalnull|Apical|Modifier|false|false||apicalnull|Hypokinesia|Finding|false|false||hypokinesisnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Thrombus|Finding|true|false|C4266612;C0225897;C2355627;C0018827;C0007799|thrombinull|Chest>Heart.ventricle.left|Anatomy|false|false|C1552822;C0087086|left ventricle
null|Left ventricular structure|Anatomy|false|false|C1552822;C0087086|left ventriclenull|Table Cell Horizontal Align - left|Finding|false|false|C4266612;C0225897;C2355627;C0018827;C0007799|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Heart Ventricle|Anatomy|false|false|C0087086;C1552822|ventricle
null|Cerebral Ventricles|Anatomy|false|false|C0087086;C1552822|ventricle
null|Ventricle|Anatomy|false|false|C0087086;C1552822|ventriclenull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Heart Ventricle|Anatomy|false|false||ventricularnull|Ventricular|Modifier|false|false||ventricularnull|chamber [body part]|Anatomy|false|false||chambernull|Chamber (physical object)|Device|false|false||chambernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Aortic valve structure|Anatomy|false|false||aortic valve
null|Chest>Aortic valve|Anatomy|false|false||aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Mild Severity of Illness Code|Finding|false|false|C4533215;C0003501;C1186983|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Aortic valve structure|Anatomy|false|false|C1547225|aortic valve
null|Chest>Aortic valve|Anatomy|false|false|C1547225|aortic valvenull|Aorta|Anatomy|false|false||aorticnull|Anatomical valve|Anatomy|false|false|C1547225|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Valve Area|Finding|false|false|C1186983|valve areanull|Anatomical valve|Anatomy|false|false|C1510751;C4687749;C0555206|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Academic Research Enhancement Awards|Event|false|false|C1186983|areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Chiari malformation type II|Disorder|false|false|C1186983|cm2null|sq. cm|LabModifier|false|false||cm2null|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Aortic Valve Insufficiency|Disorder|false|false|C0003483|aortic regurgitationnull|Aorta|Anatomy|false|false|C0003504|aorticnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Mitral Valve|Anatomy|false|false||mitral valvenull|mitral|Modifier|false|false||mitralnull|Anatomical valve|Anatomy|false|false||valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Mitral Valve Insufficiency|Disorder|false|false||mitral regurgitationnull|mitral|Modifier|false|false||mitralnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Pulmonary artery structure|Anatomy|false|false|C0039155;C4522268;C2707265|pulmonary arterynull|Pulmonary (intended site)|Finding|false|false|C0024109;C0034052;C0226004;C0003842|pulmonarynull|Lung|Anatomy|false|false|C2707265;C4522268|pulmonarynull|null|Attribute|false|false|C0024109;C0226004;C0003842;C0034052|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Arterial system|Anatomy|false|false|C0039155;C2707265;C4522268|artery
null|Arteries|Anatomy|false|false|C0039155;C2707265;C4522268|arterynull|Systole|Finding|false|false|C0226004;C0003842;C0034052|systolicnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Physiological|Finding|false|false||physiologicnull|Pericardial effusion|Disorder|false|false|C0031050;C0442031|pericardial effusionnull|Pericardial effusion body substance|Finding|false|false|C0031050;C0442031|pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false|C0031039;C1253937;C2317432;C1546613;C0013687|pericardial
null|Pericardial sac structure|Anatomy|false|false|C0031039;C1253937;C2317432;C1546613;C0013687|pericardialnull|Effusion (substance)|Finding|false|false|C0031050;C0442031|effusion
null|null|Finding|false|false|C0031050;C0442031|effusion
null|effusion|Finding|false|false|C0031050;C0442031|effusionnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Left ventricular cavity size|Attribute|false|false|C0507083;C0503990;C0333343;C0018827|left ventricular cavity sizenull|Cavity of left ventricle|Anatomy|false|false|C1510420;C0011334;C0455830|left ventricular cavitynull|Table Cell Horizontal Align - left|Finding|false|false|C0018827|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Cavity of ventricle|Anatomy|false|false|C0455830;C1510420;C0011334|ventricular cavitynull|Heart Ventricle|Anatomy|false|false|C1552822;C1510420;C0011334;C0455830|ventricularnull|Ventricular|Modifier|false|false||ventricularnull|Dental caries|Disorder|false|false|C0503990;C0507083;C0018827;C0333343|cavity
null|Cavitation|Disorder|false|false|C0503990;C0507083;C0018827;C0333343|cavitynull|Body cavities|Anatomy|false|false|C0455830;C1510420;C0011334|cavitynull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|regional|Modifier|false|false||regional
null|Local|Modifier|false|false||regionalnull|Systolic dysfunction|Finding|false|false||systolic dysfunctionnull|Systole|Finding|false|false||systolicnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false|C0226032|CAD
null|Coronary heart disease|Disorder|false|false|C0226032|CAD
null|Coronary Artery Disease|Disorder|false|false|C0226032|CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1956346;C0010068;C0175816;C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Distribution [PK]|Finding|false|false||distribution
null|Distribution|Finding|false|false||distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|Mild aortic valve stenosis|Disorder|false|false|C0003483;C4533215;C0003501;C1186983|Mild aortic valve stenosisnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|AORTIC VALVE DISEASE 3|Disorder|false|false|C4533215;C0003501;C0003483;C1186983|aortic valve stenosis
null|Stenosis of aorta|Disorder|false|false|C4533215;C0003501;C0003483;C1186983|aortic valve stenosisnull|Aortic Valve Stenosis|Finding|false|false|C4533215;C0003501;C0003483;C1186983|aortic valve stenosisnull|Aortic valve structure|Anatomy|false|false|C0003507;C5700069;C5193127;C3276923;C1261287|aortic valve
null|Chest>Aortic valve|Anatomy|false|false|C0003507;C5700069;C5193127;C3276923;C1261287|aortic valvenull|Aorta|Anatomy|false|false|C3276923;C0003507;C5700069;C5193127|aorticnull|Anatomical valve|Anatomy|false|false|C1261287;C0003507;C5700069;C5193127;C3276923|valvenull|Valve (physical object)|Device|false|false||valve
null|Valve Device|Device|false|false||valve
null|medical valve|Device|false|false||valvenull|Stenosis|Finding|false|false|C1186983;C4533215;C0003501|stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Mild Severity of Illness Code|Finding|false|false|C0003483|Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Aorta|Anatomy|false|false|C1547225|aorticnull|Regurgitation|Finding|false|false||regurgitation
null|Regurgitates after swallowing|Finding|false|false||regurgitationnull|Regurgitation - mechanism|Phenomenon|false|false||regurgitationnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Hypertensive disease|Disorder|false|false||hypertensionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4554413;C1272939;C0721966;C0016658;C4520890;C1522019|nasalnull|Fracture|Disorder|false|false|C0028429|fracturesnull|Fractured|Finding|false|false|C0028429|fracturesnull|Epistaxis|Finding|false|false||epistaxisnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Epistaxis|Finding|false|false||Epistaxisnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C0016658;C1272939;C0721966;C4554413|nasalnull|Fracture|Disorder|false|false|C0028429|fracturesnull|Fractured|Finding|false|false|C0028429|fracturesnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|mechanical method|Finding|false|false||mechanicalnull|Mechanical Treatments|Procedure|false|false||mechanicalnull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Continuous|Finding|false|false||ongoingnull|Epistaxis|Finding|false|false||epistaxisnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Nasal bone structure|Anatomy|false|false|C0016658;C1546560;C1550616;C4554413|nasal bonenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966|nasalnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950;C0027422|bone
null|null|Finding|false|false|C1442209;C0262950;C0027422|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|Septal|Modifier|false|false||septalnull|Fracture|Disorder|false|false|C0027422|fracturesnull|Fractured|Finding|false|false|C0027422|fracturesnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4520890;C1522019;C1272939;C0721966|nasalnull|Spray Dosage Form|Drug|false|false||spraynull|Spray (administration method)|Finding|false|false||spraynull|Spray (action)|Event|false|false||spraynull|Spray Dosing Unit|LabModifier|false|false||spraynull|Hold - dosing instruction fragment|Finding|false|false||hold
null|hold - Data Operation|Finding|false|false||holdnull|Hold (action)|Event|false|false||holdnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Hemorrhage|Finding|false|false||bleedingnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Troponin|Drug|false|false||troponin
null|Troponin|Drug|false|false||troponinnull|Troponin measurement|Procedure|false|false||troponinnull|Protein Component|Drug|false|false||component
null|Protein Component|Drug|false|false||componentnull|Component, LOINC Axis 1|Finding|false|false||component
null|Specimen Child Role - Component|Finding|false|false||component
null|Component (part)|Finding|false|false||componentnull|Component object|Device|false|false||componentnull|Course|Time|false|false||coursenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0008031;C0741025;C2926613;C1549543;C0030193|chest
null|Anterior thoracic region|Anatomy|false|false|C0008031;C0741025;C2926613;C1549543;C0030193|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|cardiac symptom|Finding|false|false|C0018787|cardiac symptomsnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C0741933;C0683368;C1457887;C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Symptoms aspect|Finding|false|false|C0018787|symptoms
null|Symptoms|Finding|false|false|C0018787|symptomsnull|Cardiovascular system|Anatomy|false|false||Cardiologynull|cardiology (field)|Title|false|false||Cardiologynull|Cardiology service|Entity|false|false||Cardiologynull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Economic demand|Finding|false|false||demandnull|Demand (clinical)|Procedure|false|false||demandnull|Ischemia|Finding|false|false||ischemianull|Ischemia Procedure|Procedure|false|false||ischemianull|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Falls|Finding|false|false||fallnull|Autumn|Time|false|false||fallnull|Echocardiography|Procedure|false|false||echocardiogramnull|Aortic Valve Stenosis|Finding|false|false|C0003483|aortic stenosisnull|Aorta|Anatomy|false|false|C0003507|aorticnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Probable diagnosis|Finding|false|false|C0226032|likely
null|Probably|Finding|false|false|C0226032|likelynull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C0012634;C0332148;C0750492;C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Disease|Disorder|false|false|C0226032|diseasenull|Wall motion|Attribute|false|false||wall motionnull|Walls of a building|Device|false|false||wallnull|Motion|Phenomenon|false|false||motionnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|pravastatin|Drug|false|false||pravastatin
null|pravastatin|Drug|false|false||pravastatinnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Hypoxemia|Finding|false|false||Hypoxemia
null|Blood oxygen concentration below reference range (finding)|Finding|false|false||Hypoxemianull|Basilar|Modifier|false|false||basilarnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|Hypoxia|Finding|false|false||hypoxicnull|Oxygen Saturation|Attribute|false|false||oxygen saturationsnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Saturated|Phenomenon|false|false||saturationsnull|on room air|Finding|false|false||on room airnull|Room Air|Drug|false|false||room airnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Fever|Finding|false|false||feversnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Plain chest X-ray|Procedure|false|false||CXRnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Left lung|Anatomy|false|false|C0332149;C0740941;C0445223;C1552599;C0700198;C0851353;C1552822;C4319827;C0039869;C1720922;C0005768;C0229664;C0005767;C0024115|left lungnull|Table Cell Horizontal Align - left|Finding|false|false|C0225730;C4037972;C0024109|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lung diseases|Disorder|false|false|C4037972;C0024109;C0225730|lungnull|Lung Problem|Finding|false|false|C0225730;C4037972;C0024109|lungnull|Chest>Lung|Anatomy|false|false|C0332149;C1720922;C4319827;C0039869;C0024115;C0700198;C0740941;C1552822|lung
null|Lung|Anatomy|false|false|C0332149;C1720922;C4319827;C0039869;C0024115;C0700198;C0740941;C1552822|lungnull|Thought|Finding|false|false|C4037972;C0024109;C0225730|thought
null|null|Finding|false|false|C4037972;C0024109;C0225730|thoughtnull|Possibly Related to Intervention|Modifier|false|false||possibly relatednull|Possible|Finding|false|false|C0225730;C4037972;C0024109|possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false|C0225730|related
null|Related (finding)|Finding|false|false|C0225730|relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Respiratory Aspiration|Disorder|false|false|C4037972;C0024109;C0225730|aspiratednull|Pulmonary aspiration|Finding|false|false|C4037972;C0024109;C0225730|aspiratednull|Blood and lymphatic system disorders|Disorder|false|false|C0225730|bloodnull|In Blood|Finding|false|false|C0225730|blood
null|peripheral blood|Finding|false|false|C0225730|blood
null|Blood|Finding|false|false|C0225730|bloodnull|Monitor brand of insecticide|Drug|false|false||monitor
null|Monitor brand of insecticide|Drug|false|false||monitornull|Monitor Device|Device|false|false||monitor
null|Monitoring Device|Device|false|false||monitornull|Monitor, occupation|Subject|false|false||monitornull|Oxygen saturation measurement|Procedure|false|false||O2 saturationnull|Saturated|Phenomenon|false|false||saturationnull|Body temperature measurement|Procedure|false|false||temperaturenull|Body Temperature|Subject|false|false||temperaturenull|Temperature|LabModifier|false|false||temperaturenull|null|Attribute|false|false||trendnull|trend|Time|false|false||trendnull|Leukocytes|Anatomy|false|false||WBCnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Acute kidney injury|Disorder|false|false|C0227665;C0022646|Acute kidney injury
null|Kidney Failure, Acute|Disorder|false|false|C0227665;C0022646|Acute kidney injurynull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Injury of kidney|Disorder|false|false|C0227665;C0022646|kidney injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0160420;C0022660;C2609414;C0812426;C0496927;C0496892;C4554465;C0869841;C3263723;C3263722|kidney
null|Both kidneys|Anatomy|false|false|C0160420;C0022660;C2609414;C0812426;C0496927;C0496892;C4554465;C0869841;C3263723;C3263722|kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false|C0227665;C0022646|injury
null|Traumatic injury|Disorder|false|false|C0227665;C0022646|injurynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Last|Modifier|false|false||lastnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|unaware|Procedure|false|false||unawarenull|null|Finding|false|false|C0227665;C0022646|history of kidney diseasenull|Medical History|Finding|false|false|C0227665;C0022646|history ofnull|History of present illness (finding)|Finding|false|false|C0227665;C0022646|history
null|History of previous events|Finding|false|false|C0227665;C0022646|history
null|Historical aspects qualifier|Finding|false|false|C0227665;C0022646|history
null|Medical History|Finding|false|false|C0227665;C0022646|history
null|Concept History|Finding|false|false|C0227665;C0022646|historynull|History|Subject|false|false||historynull|Kidney Diseases|Disorder|false|false|C0227665;C0022646|kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|kidneynull|Kidney|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0262926;C0012634;C0022658;C0455686;C0812426;C0262926;C1705255;C0019665;C0262512;C2004062|kidney
null|Both kidneys|Anatomy|false|false|C0496927;C0496892;C4554465;C0869841;C0262926;C0012634;C0022658;C0455686;C0812426;C0262926;C1705255;C0019665;C0262512;C2004062|kidneynull|Disease|Disorder|false|false|C0227665;C0022646|diseasenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Peripheral Vascular Diseases|Disorder|false|false|C0005847|Peripheral vascular diseasenull|Peripheral|Modifier|false|false||Peripheralnull|Vascular Diseases|Disorder|false|false|C0005847|vascular diseasenull|Blood Vessel|Anatomy|false|false|C0085096;C0012634;C0042373|vascularnull|Vascular|Modifier|false|false||vascularnull|Disease|Disorder|false|false|C0005847|diseasenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|AAA brand of benzocaine-cetalkonium chloride combination|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAA
null|APP protein, human|Drug|false|false||AAAnull|Aortic Aneurysm, Abdominal|Disorder|false|false||AAA
null|Aortic Aneurysm|Disorder|false|false||AAAnull|AAAS wt Allele|Finding|false|false||AAA
null|APP gene|Finding|false|false||AAA
null|APP wt Allele|Finding|false|false||AAAnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|false|false||historynull|Coronary Artery Bypass Surgery|Procedure|true|false||CABGnull|Cardiac attachment|Finding|true|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Peripheral|Modifier|false|false||peripheralnull|null|Device|false|false||stentsnull|Cardiac attachment|Finding|false|false|C0018787|cardiacnull|Heart|Anatomy|false|false|C5237222;C0040808;C1314974|cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|GDC Regimen Terminology|Finding|false|false|C0018787|regimennull|Treatment Protocols|Procedure|false|false|C0018787|regimennull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|Echocardiography, Stress|Procedure|false|false|C0226032|stress echonull|Stress bismuth subsalicylate|Drug|false|false||stress
null|Stress bismuth subsalicylate|Drug|false|false||stressnull|Stress|Finding|false|false||stressnull|W stress|Attribute|false|false||stressnull|Extension for Community Healthcare Outcomes|Procedure|false|false|C0226032|echo
null|ECHO protocol|Procedure|false|false|C0226032|echonull|Echo <Calopterygidae>|Entity|false|false||echonull|Processing type - Evaluation|Finding|false|false|C0226032|evaluationnull|Evaluation procedure|Procedure|false|false|C0226032|evaluation
null|Evaluation|Procedure|false|false|C0226032|evaluationnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C0920208;C0012634;C1550157;C5575284;C0058928;C1261322;C0220825;C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|false|false||LADnull|Disease|Disorder|false|false|C0226032|diseasenull|Possible|Finding|false|false||possiblynull|Possible diagnosis|Modifier|false|false||possiblynull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Territory|Entity|false|false||territory
null|Geographic state|Entity|false|false||territorynull|At risk|Modifier|false|false||at risknull|Risk|Finding|false|false||risknull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Echocardiography|Procedure|false|false||echocardiogramnull|year|Time|false|false||yearsnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Epistaxis|Finding|false|false||epistaxisnull|Nasal Spray brand of phenylephrine|Drug|false|false|C0028429|nasal spraynull|Nasal spray (device)|Device|false|false||nasal spray
null|Nasal Sprays|Device|false|false||nasal spray
null|Nasal Spray|Device|false|false||nasal spraynull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C4521772;C4520890;C1522019;C1272939;C0721966;C2608294|nasalnull|Spray Dosage Form|Drug|false|false||spraynull|Spray (administration method)|Finding|false|false|C0028429|spraynull|Spray (action)|Event|false|false||spraynull|Spray Dosing Unit|LabModifier|false|false||spraynull|Repeat Object|Finding|false|false|C1261077;C1527391;C0817096|Repeat
null|Repeat|Finding|false|false|C1261077;C1527391;C0817096|Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Plain chest X-ray|Procedure|false|false|C1261077;C1527391;C0817096|chest x-raynull|Chest problem|Finding|false|false|C1261077;C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0043299;C1962945;C1306645;C0034571;C3244296;C0043309;C1705914;C0205341;C0039985;C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0043299;C1962945;C1306645;C0034571;C3244296;C0043309;C1705914;C0205341;C0039985;C0741025|chestnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false|C1527391;C0817096;C1261077|x-ray
null|roentgenographic|Finding|false|false|C1527391;C0817096;C1261077|x-raynull|Plain x-ray|Procedure|false|false|C1261077;C1527391;C0817096|x-ray
null|Diagnostic radiologic examination|Procedure|false|false|C1261077;C1527391;C0817096|x-ray
null|Radiographic imaging procedure|Procedure|false|false|C1261077;C1527391;C0817096|x-raynull|Roentgen Rays|Phenomenon|false|false|C1527391;C0817096;C1261077|x-raynull|week|Time|false|false||weeksnull|physiologic resolution|Finding|false|false|C1261077|resolution
null|Resolution|Finding|false|false|C1261077|resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Structure of left lower lobe of lung|Anatomy|false|false|C0043299;C1962945;C1306645;C1705914;C0205341;C0039985;C0034571;C3244296;C0741025;C0043309;C1514893;C2699488|LLLnull|Infiltrative Tumor Margin|Finding|false|false|C1184743|infiltrativenull|Process Pharmacologic Substance|Drug|false|false|C1184743|processnull|Process (qualifier value)|Finding|false|false|C1184743|processnull|bony process|Anatomy|false|false|C1951340;C4521054;C4527217;C1522240|processnull|Process|Phenomenon|false|false|C1184743|processnull|consider|Finding|false|false||Considernull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|ENT problem|Finding|false|false|C0150934;C0175196|ENT
null|NT5E gene|Finding|false|false|C0150934;C0175196|ENT
null|NT5E wt Allele|Finding|false|false|C0150934;C0175196|ENTnull|Structure of entorhinal cortex|Anatomy|false|false|C0262471;C3889152;C1417861|ENT
null|Ear, nose and throat|Anatomy|false|false|C0262471;C3889152;C1417861|ENTnull|Otolaryngology specialty|Title|false|false||ENTnull|Plastic Surgical Procedures|Procedure|false|false||Plastic Surgerynull|Plastic Surgery Specialty|Title|false|false||Plastic Surgerynull|Plastics|Drug|false|false||Plasticnull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Late|Time|false|false||laternull|Processing type - Evaluation|Finding|false|false|C0028429|evaluationnull|Evaluation procedure|Procedure|false|false|C0028429|evaluation
null|Evaluation|Procedure|false|false|C0028429|evaluationnull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|nasal
null|Nasal dosage form|Drug|false|false|C0028429|nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|nasal
null|Nasal (intended site)|Finding|false|false|C0028429|nasalnull|null|Anatomy|false|false|C0016658;C4554413;C1272939;C0721966;C4520890;C1522019;C1550157;C1261322;C0220825|nasalnull|Fracture|Disorder|false|false|C0028429|fracturesnull|Fractured|Finding|false|false|C0028429|fracturesnull|Repeat Object|Finding|false|false|C2263086|Repeat
null|Repeat|Finding|false|false|C2263086|Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C1561540;C0009555;C0472699;C0018935;C1705914;C0205341|CBCnull|1 Week|Time|false|false||one weeknull|Transaction counts and value totals - week|Finding|false|false|C2263086|weeknull|week|Time|false|false||weeknull|Medical Product Stability|Modifier|false|false||stability
null|Stable status|Modifier|false|false||stabilitynull|Hemopoietic stem cell transplant|Procedure|false|false|C2263086|HCT
null|Hematocrit Measurement|Procedure|false|false|C2263086|HCTnull|Platelets Product|Drug|false|false|C0005821|plateletsnull|Platelet count (procedure)|Procedure|false|false|C0005821|plateletsnull|Blood Platelets|Anatomy|false|false|C0443116;C0032181|plateletsnull|consider|Finding|false|false||Considernull|Conversions (qualifier value)|Finding|false|false||conversionnull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|succinate|Drug|false|false||succinate
null|Succinates|Drug|false|false||succinatenull|Comfort|Finding|false|false||easenull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|pravastatin|Drug|false|false||Pravastatin
null|pravastatin|Drug|false|false||Pravastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|clopidogrel|Drug|false|false||Clopidogrel
null|clopidogrel|Drug|false|false||Clopidogrelnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|null|Drug|false|false||NSAID
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|ibuprofen|Drug|false|false||ibuprofen
null|ibuprofen|Drug|false|false||ibuprofennull|Hemorrhage|Finding|false|false||bleedingnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|30 days|Time|false|false||30 Daysnull|day|Time|false|false||Daysnull|metoprolol tartrate|Drug|false|false||Metoprolol Tartrate
null|metoprolol tartrate|Drug|false|false||Metoprolol Tartratenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C5975557|mouth
null|Oral region|Anatomy|false|false|C1527415;C5975557|mouthnull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false|C0230028;C0226896|timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C2828567;C1527415|mouth
null|Oral region|Anatomy|false|false|C2828567;C1527415|mouthnull|Every evening|Modifier|false|false||every eveningnull|Evening|Time|false|false||eveningnull|PRSS30P gene|Finding|false|false|C0230028;C0226896|Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|oxymetazoline|Drug|false|false||Oxymetazoline
null|oxymetazoline|Drug|false|false||Oxymetazolinenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Counter brand of Terbufos|Drug|false|false||counter
null|Counter brand of Terbufos|Drug|false|false||counternull|Counter device|Device|false|false||counternull|Proprietary Name|Finding|false|false||brand namenull|MDF Attribute Type - Name|Finding|false|false||name
null|Person Name|Finding|false|false||name
null|Name|Finding|false|false||namenull|Name (property) (qualifier value)|Modifier|false|false||namenull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Fractured nasal bones|Disorder|false|false|C0028429|Nasal fracturenull|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal brand of oxymetazoline|Drug|false|false|C0028429|Nasal
null|Nasal dosage form|Drug|false|false|C0028429|Nasalnull|Nasal Route of Administration|Finding|false|false|C0028429|Nasal
null|Nasal (intended site)|Finding|false|false|C0028429|Nasalnull|null|Anatomy|false|false|C1272939;C0721966;C0016658;C4520890;C1522019;C0339848|Nasalnull|Fracture|Disorder|false|false|C0028429|fracturenull|Epistaxis|Finding|false|false||Epistaxisnull|null|Disorder|false|false||NSTEMInull|null|Finding|false|false||NSTEMInull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Hemorrhage|Finding|false|false||bleedsnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Plug (physical object)|Device|false|false||plugsnull|Hemorrhage|Finding|false|false||bleedingnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Troponin|Drug|false|false||troponins
null|Troponin|Drug|false|false||troponinsnull|Hematologic Tests|Procedure|false|false|C4318744|blood testnull|Blood test device|Device|false|false||blood testnull|Blood and lymphatic system disorders|Disorder|false|false|C4318744|bloodnull|peripheral blood|Finding|false|false|C4318744|blood
null|Blood|Finding|false|false|C4318744|blood
null|In Blood|Finding|false|false|C4318744|bloodnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C0022885;C0456984;C0018941;C0005768;C0229664;C0005767;C0039593;C0392366;C0851353|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heart
null|Heart|Anatomy|false|false|C0153957;C0153500;C0795691|heartnull|Ultrasonic|Finding|false|false|C4037974;C0018787|ultrasoundnull|Urological ultrasound|Procedure|false|false|C4037974;C0018787|ultrasound
null|Ultrasonography|Procedure|false|false|C4037974;C0018787|ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false|C4037974;C0018787|ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false|C4037974;C0018787|ultrasoundnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C1315081;C0041618;C0795691;C0220934;C0153957;C0153500;C0041621;C1456803|heart
null|Heart|Anatomy|false|false|C1315081;C0041618;C0795691;C0220934;C0153957;C0153500;C0041621;C1456803|heartnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Exercise stress test|Procedure|false|false|C4318744|stress test
null|Stress Test|Procedure|false|false|C4318744|stress testnull|Stress bismuth subsalicylate|Drug|false|false|C4318744|stress
null|Stress bismuth subsalicylate|Drug|false|false|C4318744|stressnull|Stress|Finding|false|false|C4318744|stressnull|W stress|Attribute|false|false|C4318744|stressnull|Tests (qualifier value)|Finding|false|false|C4318744|test
null|Testing|Finding|false|false|C4318744|testnull|Laboratory Procedures|Procedure|false|false|C4318744|testnull|Test - temporal region|Anatomy|false|false|C1718621;C0723460;C0022885;C0038435;C0039593;C0392366;C0456984;C0015260;C3494508|testnull|Test Result|Lab|false|false|C4318744|testnull|Test Dosing Unit|LabModifier|false|false||testnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Choose (action)|Event|false|false||choosingnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions