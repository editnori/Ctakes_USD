CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|sulfa|Drug|false|false||Sulfanull|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamide [EPC]|Drug|false|false||Sulfonamidenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Bactrim|Drug|false|false||Bactrim
null|Bactrim|Drug|false|false||Bactrimnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Percutaneous liver biopsy|Procedure|false|false||Percutaneous liver biopsynull|Percutaneous Route of Drug Administration|Finding|false|false||Percutaneousnull|Percutaneous|Modifier|false|false||Percutaneousnull|Consent Type - Liver Biopsy|Procedure|false|false||liver biopsy
null|Biopsy of liver (procedure)|Procedure|false|false||liver biopsynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Known|Modifier|false|false||knownnull|Lesion|Finding|false|false||lesionsnull|Lung|Anatomy|false|false||lungsnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Breath|Finding|false|false||breathnull|Initially|Time|false|false||initiallynull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Processing type - Evaluation|Finding|false|false||Evaluationnull|Evaluation procedure|Procedure|false|false||Evaluation
null|Evaluation|Procedure|false|false||Evaluationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|CT of abdomen|Procedure|false|false||abdominal CT scannull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Numerous|LabModifier|false|false||multiplenull|Lung and Liver|Anatomy|false|false||lung and livernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Definitely Related to Intervention|Modifier|false|false||definite
null|Definite|Modifier|false|false||definitenull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Recent|Time|false|false||recentnull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|Documentation|Finding|false|false||documentationnull|Act of Documentation|Procedure|false|false||documentationnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Usual|Modifier|false|false||usualnull|personal health|Finding|false|false||state of healthnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Health|Finding|false|false||healthnull|Evening|Time|false|false||eveningnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Acute-on-chronic|Time|false|false||acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|ACHE protein, human|Drug|false|false||ache
null|acetylcholinesterase|Drug|false|false||ache
null|acetylcholinesterase|Drug|false|false||ache
null|ACHE protein, human|Drug|false|false||achenull|ACHE Gene|Finding|false|false||ache
null|Pain|Finding|false|false||ache
null|Ache|Finding|false|false||achenull|Associated with|Modifier|false|false||associated withnull|Associated with|Modifier|false|false||associatednull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Direct - PostalAddressUse|Finding|false|false||direct
null|direct address|Finding|false|false||directnull|Direct type of relationship|Modifier|false|false||direct
null|Direct (qualifier)|Modifier|false|false||directnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|exercise induced|Finding|false|false||exertionalnull|Protein Component|Drug|true|false||component
null|Protein Component|Drug|true|false||componentnull|Specimen Child Role - Component|Finding|true|false||component
null|Component (part)|Finding|true|false||component
null|Component, LOINC Axis 1|Finding|true|false||componentnull|Component object|Device|true|false||componentnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Smear - instruction imperative|Event|false|false||spreadnull|Spreading (qualifier value)|Modifier|false|false||spreadnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|null|Time|false|false||precedingnull|month|Time|false|false||monthsnull|Recent|Time|false|false||recentlynull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Greater|LabModifier|false|false||greaternull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Edema of lower extremity|Finding|false|false||lower extremity edemanull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false||extremity edemanull|Limb structure|Anatomy|false|false||extremitynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Veins|Anatomy|false|false||venousnull|Venous|Modifier|false|false||venousnull|Ultrasonography|Procedure|false|false||ultrasoundsnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Changing|Finding|true|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Visit|Finding|false|false||visitnull|Associated with|Modifier|false|false||associatednull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Sweating|Finding|false|false||sweats
null|Sweat|Finding|false|false||sweatsnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|positional|Finding|false|false||positionalnull|Protein Component|Drug|false|false||component
null|Protein Component|Drug|false|false||componentnull|Specimen Child Role - Component|Finding|false|false||component
null|Component (part)|Finding|false|false||component
null|Component, LOINC Axis 1|Finding|false|false||componentnull|Component object|Device|false|false||componentnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Laboratory test finding|Lab|false|false||Labsnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Urinalysis; qualitative or semiquantitative, except immunoassays|Procedure|false|false||Urinalysis
null|Urinalysis|Procedure|false|false||Urinalysisnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Epithelial|Modifier|false|false||epithelialnull|Cells|Anatomy|false|false||cellsnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Central brand of multivitamin with minerals|Drug|false|false||central
null|Central brand of multivitamin with minerals|Drug|false|false||centralnull|Central Minus|Procedure|false|false||centralnull|Central|Modifier|false|false||centralnull|Pulmonary Embolism|Finding|false|false||pulmonary embolusnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|null|Finding|false|false||embolus
null|Embolus|Finding|false|false||embolusnull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Registry to Evaluate Early and Long-Term Pulmonary Arterial (PAH) Hypertension Disease Management (REVEAL)|Finding|false|false||revealnull|Revealed|Modifier|false|false||revealnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Hepatomegaly|Finding|false|false||enlarged livernull|Enlargement procedure|Procedure|false|false||enlargednull|Enlarged|Modifier|false|false||enlargednull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus Tachycardia|Disorder|false|false||sinus tachycardianull|continuous electrocardiogram sinus tachycardia|Finding|false|false||sinus tachycardia
null|Sinus Tachycardia by ECG Finding|Finding|false|false||sinus tachycardianull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Overall Publication Type|Finding|false|false||overallnull|Overall|Modifier|false|false||overallnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|null|Time|false|false||priornull|ceftriaxone|Drug|false|false||Ceftriaxone
null|ceftriaxone|Drug|false|false||Ceftriaxonenull|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycin
null|azithromycin|Drug|false|false||azithromycinnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Pneumonia|Disorder|false|false||pneumonianull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Pain-Free|Drug|false|false||pain freenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|ATP5F1A gene|Finding|false|false||OMRnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Enneking High Surgical Grade|Finding|false|false||high grade
null|Severe (severity modifier)|Finding|false|false||high gradenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Histopathologic Grade|Finding|false|false||grade
null|Grade|Finding|false|false||grade
null|School Grade|Finding|false|false||gradenull|Exploratory laparotomy|Procedure|false|false||exploratory laparotomynull|Laparotomy|Procedure|false|false||laparotomynull|Lysis|Finding|false|false||lysis
null|pathologic cytolysis|Finding|false|false||lysisnull|Tissue Adhesions|Finding|false|false||adhesionsnull|Small intestine excision|Procedure|false|false||small bowel resectionnull|Abdomen>Small bowel|Anatomy|false|false||small bowel
null|Intestines, Small|Anatomy|false|false||small bowelnull|Small|LabModifier|false|false||smallnull|Bowel resection|Procedure|false|false||bowel resectionnull|Intestines|Anatomy|false|false||bowelnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Anastomosis of small intestine to small intestine|Procedure|false|false||enteroenterostomy
null|Anastomosis of intestine|Procedure|false|false||enteroenterostomynull|Carcinoid Tumor|Disorder|false|false||carcinoidnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Vitamin B 12 Deficiency|Disorder|false|false||vitamin B12 deficiencynull|Decreased circulating vitamin B12 concentration|Finding|false|false||vitamin B12 deficiencynull|Vitamin B12 [EPC]|Drug|false|false||vitamin B12
null|cobalamins|Drug|false|false||vitamin B12
null|cobalamins|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12
null|vitamin B12|Drug|false|false||vitamin B12null|VITAMIN B12 MEASUREMENT|Procedure|false|false||vitamin B12null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|TNFAIP1 wt Allele|Finding|false|false||B12
null|NDUFB3 gene|Finding|false|false||B12
null|TNFAIP1 gene|Finding|false|false||B12null|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Neck|Anatomy|false|false||cervicalnull|Cervical|Modifier|false|false||cervicalnull|Degenerative polyarthritis|Disorder|false|false||DJDnull|Degenerative polyarthritis|Disorder|false|false||osteoarthritisnull|Lung excision|Procedure|false|false||lung resectionnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|removal technique|Procedure|false|false||resection
null|Excision|Procedure|false|false||resectionnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Right arm|Anatomy|false|false||R armnull|Anorectal Malformations|Disorder|false|false||armnull|AKR1A1 wt Allele|Finding|false|false||arm
null|ARMC9 gene|Finding|false|false||armnull|Protocol Treatment Arm|Procedure|false|false||arm
null|Axillary Reverse Mapping|Procedure|false|false||arm
null|Study Arm|Procedure|false|false||armnull|Upper arm|Anatomy|false|false||arm
null|null|Anatomy|false|false||arm
null|Upper Extremity|Anatomy|false|false||armnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|ATP5F1A gene|Finding|false|false||OMRnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Cessation of life|Finding|false|false||Died
null|Death (finding)|Finding|false|false||Died
null|Dead (finding)|Finding|false|false||Diednull|Malignant neoplasm of pancreas|Disorder|false|false||pancreatic cancer
null|Pancreatic carcinoma|Disorder|false|false||pancreatic cancernull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false||pancreaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Glycation End Products, Advanced|Drug|false|true||age
null|Glycation End Products, Advanced|Drug|false|true||agenull|null|Attribute|false|true||agenull|Age|Subject|false|false||agenull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Cessation of life|Finding|false|false||Died
null|Death (finding)|Finding|false|false||Died
null|Dead (finding)|Finding|false|false||Diednull|Disease|Disorder|false|false||diseasenull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||sinusnull|pathologic fistula|Disorder|false|false||sinusnull|Sinus - general anatomical term|Anatomy|false|false||sinus
null|Nasal sinus|Anatomy|false|false||sinusnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Full|Modifier|false|false||fullnull|Sentence|Finding|false|false||sentencesnull|HEENT|Anatomy|false|false||HEENTnull|PERRLA|Finding|false|false||PERRLAnull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Jugular venous engorgement|Finding|true|false||JVDnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Palp - CHV concept|Finding|false|false||palp
null|ALPP gene|Finding|false|false||palp
null|ALPP wt Allele|Finding|false|false||palpnull|Palpable|Modifier|false|false||palpablenull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Lung|Anatomy|false|false||LUNGSnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|aeration|Procedure|false|false||aerationnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||respnull|Respiratory rate|Attribute|false|false||respnull|Unlabored|Finding|false|false||unlaborednull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Malignant neoplasm of heart|Disorder|false|false||HEART
null|benign neoplasm of heart|Disorder|false|false||HEARTnull|HEART PROBLEM|Finding|false|false||HEARTnull|Chest>Heart|Anatomy|false|false||HEART
null|Heart|Anatomy|false|false||HEARTnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Heart Sounds|Finding|false|false||heart soundsnull|auscultation of heart sounds|Procedure|false|false||heart soundsnull|null|Attribute|false|false||heart soundsnull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Regular|Modifier|false|false||regularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|SYSTOLIC EJECTION MURMUR|Finding|false|false||SEMnull|Microscopes, Electron, Scanning|Device|false|false||SEMnull|Standard Error|LabModifier|false|false||SEMnull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Palp - CHV concept|Finding|false|false||palp
null|ALPP gene|Finding|false|false||palp
null|ALPP wt Allele|Finding|false|false||palpnull|More|LabModifier|false|false||morenull|Structure of right upper quadrant of abdomen|Anatomy|false|false||RUQnull|RUQ - Right upper quadrant|Modifier|false|false||RUQnull|Protective muscle spasm|Finding|false|false||guardingnull|Liver palpable|Finding|false|false||palpable livernull|Palpable|Modifier|false|false||palpablenull|Liver edge|Finding|false|false||liver edgenull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|1+ pitting edema|Finding|false|false||1+ pitting edemanull|Pitting edema|Finding|false|false||pitting edemanull|Pitting|Finding|false|false||pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Middle|Modifier|false|false||midnull|Shin|Anatomy|false|false||shinnull|null|Finding|false|false||pulses radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Awake (finding)|Finding|false|false||awakenull|Awakening (time frame)|Time|false|false||awakenull|Central Nervous System|Anatomy|false|false||CNsnull|Clinical Nurse Specialists|Subject|false|false||CNsnull|Certified Nurse Specialist|Title|false|false||CNsnull|Staphylococcus, coagulase negative (organism)|Entity|false|false||CNsnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Muscle Strength|Finding|false|false||muscle strengthnull|null|Attribute|false|false||muscle strengthnull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|At discharge|Time|false|false||At dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Obesity|Disorder|false|false||obesenull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Flat affect|Finding|false|false||flat affectnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Poor eye contact|Finding|false|false||poor eye contactnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|eye contact|Finding|false|false||eye contactnull|Carcinoma in situ of eye|Disorder|false|false||eye
null|Disorder of eye|Disorder|false|false||eyenull|Eye - Specimen Source Code|Finding|false|false||eye
null|Eye problem|Finding|false|false||eye
null|Eye Specimen|Finding|false|false||eyenull|Head>Eye|Anatomy|false|false||eye
null|Eye|Anatomy|false|false||eye
null|Orbital region|Anatomy|false|false||eyenull|Contact - HL7 Attribution|Finding|false|false||contact
null|Contact with|Finding|false|false||contact
null|Communication Contact|Finding|false|false||contactnull|contact person|Subject|false|false||contactnull|Physical contact|Phenomenon|false|false||contactnull|Personal Contact|Event|false|false||contactnull|HEENT|Anatomy|false|false||HEENTnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Scleral icterus|Finding|false|false||scleral icterusnull|Sclera|Anatomy|false|false||scleralnull|Icterus|Finding|false|false||icterusnull|Icterus <Icteridae>|Entity|false|false||icterusnull|null|LabModifier|false|false||icterusnull|Pink color|Modifier|false|false||pinknull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Poor dentition|Finding|false|false||poor dentitionnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Dentition|Anatomy|false|false||dentition
null|Tooth structure|Anatomy|false|false||dentitionnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Malignant neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Benign neoplasm of conjunctiva|Disorder|false|false||conjunctiva
null|Conjunctival Diseases|Disorder|false|false||conjunctivanull|Specimen Type - Conjunctiva|Finding|false|false||conjunctiva
null|null|Finding|false|false||conjunctivanull|examination of conjunctiva|Procedure|false|false||conjunctiva
null|Procedure on conjunctiva|Procedure|false|false||conjunctivanull|Structure of palpebral conjunctiva|Anatomy|false|false||conjunctiva
null|conjunctiva|Anatomy|false|false||conjunctivanull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Supple|Finding|false|false||supplenull|Leukocyte adhesion deficiency type 1|Disorder|true|false||LAD
null|Leukocyte adhesion deficiency|Disorder|true|false||LADnull|ITGB2 wt Allele|Finding|true|false||LAD
null|DLD gene|Finding|true|false||LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false||LADnull|Ladino Language|Entity|true|false||LADnull|Cardiac attachment|Finding|false|false||CARDIACnull|Heart|Anatomy|false|false||CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|Regular|Modifier|false|false||regularnull|Lung diseases|Disorder|false|false||LUNGnull|Lung Problem|Finding|false|false||LUNGnull|Chest>Lung|Anatomy|false|false||LUNG
null|Lung|Anatomy|false|false||LUNGnull|cetrimonium bromide|Drug|false|false||CTABnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Decreased breath sounds|Finding|false|false||decreased breath soundsnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Assessment of body build|Procedure|false|false||body habitusnull|Document Body|Finding|false|false||bodynull|Structure of body of caudate nucleus|Anatomy|false|false||body
null|Human body structure|Anatomy|false|false||body
null|Body structure|Anatomy|false|false||body
null|Adult human body|Anatomy|false|false||body
null|Whole body|Anatomy|false|false||bodynull|Human body|Subject|false|false||bodynull|Mobility finding|Finding|false|false||mobilitynull|Range of Motion, Articular|Attribute|false|false||mobilitynull|Mobility (attribute)|Modifier|false|false||mobilitynull|Use of accessory muscles|Finding|true|false||accessory muscle usenull|Accessory skeletal muscle|Disorder|true|false||accessory musclenull|Accessory|Device|true|false||accessorynull|Muscle (organ)|Anatomy|false|false||muscle
null|Muscle Tissue|Anatomy|false|false||musclenull|Use - dosing instruction imperative|Finding|true|false||use
null|utilization qualifier|Finding|true|false||use
null|Usage|Finding|true|false||usenull|Malignant neoplasm of abdomen|Disorder|false|false||ABDOMENnull|Abdomen problem|Finding|false|false||ABDOMENnull|Abdomen|Anatomy|false|false||ABDOMEN
null|Abdominal Cavity|Anatomy|false|false||ABDOMENnull|Obesity|Disorder|false|false||obesenull|Protective muscle spasm|Finding|false|false||guardingnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Firmness|Modifier|false|false||firmnessnull|Abdomen|Anatomy|false|false||abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|1+ pitting edema|Finding|false|false||1+ pitting edemanull|Pitting edema|Finding|false|false||pitting edemanull|Pitting|Finding|false|false||pittingnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Neurology speciality|Title|false|false||NEUROnull|Neurologic (qualifier value)|Modifier|false|false||NEUROnull|Asterixis|Finding|true|false||asterixisnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Movement|Finding|false|false||movementnull|Gravity (physical force)|Phenomenon|false|false||gravitynull|Gravity - Unit of Force|LabModifier|false|false||gravitynull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Set of muscles|Anatomy|false|false||muscles
null|Muscle (organ)|Anatomy|false|false||muscles
null|Muscle Tissue|Anatomy|false|false||musclesnull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Hand problem|Finding|false|false||handnull|Upper extremity>Hand|Anatomy|false|false||hand
null|Hand|Anatomy|false|false||handnull|null|Attribute|false|false||grip strengthnull|Grip strength|Subject|false|false||grip strengthnull|Hand Strength|LabModifier|false|false||grip strengthnull|Influenza|Disorder|false|false||gripnull|grasp|Finding|false|false||gripnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false||ALT
null|Atypical Lipoma|Disorder|false|false||ALTnull|null|Finding|false|false||ALT
null|Alternative Billing Concepts|Finding|false|false||ALT
null|GPT gene|Finding|false|false||ALTnull|Antibiotic Lock Therapy|Procedure|false|false||ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Creatine Kinase|Drug|false|false||CPK
null|Creatine Kinase|Drug|false|false||CPKnull|PIK3C2A gene|Finding|false|false||CPKnull|Creatine kinase measurement|Procedure|false|false||CPKnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MB
null|Creatine Kinase MB Isoenzyme|Drug|false|false||CK-MBnull|creatine kinase activity|Finding|false|false||CK-MBnull|Serum creatine phosphokinase MB isoenzyme measurement|Procedure|false|false||CK-MB
null|Creatine kinase MB measurement|Procedure|false|false||CK-MBnull|CD79A wt Allele|Finding|false|false||MB-1
null|CD79A gene|Finding|false|false||MB-1null|Blood albumin|Procedure|false|false||BLOOD Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Albumin|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumins|Drug|false|false||Albumin
null|Albumin|Drug|false|false||Albuminnull|Albumin metabolic function|Finding|false|false||Albumin
null|ALB gene|Finding|false|false||Albuminnull|Albumin measurement|Procedure|false|false||Albuminnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Yellow color|Modifier|false|false||YELLOWnull|Cloudy|Modifier|false|false||Cloudynull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||Ketonenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||MODnull|null|Lab|false|false||URINE RBC
null|Red blood cells urine positive|Lab|false|false||URINE RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Leukocytes|Anatomy|false|false||WBCnull|Yeast, Dried|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeastnull|Saccharomyces cerevisiae|Entity|false|false||Yeast
null|Yeasts|Entity|false|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|At discharge|Time|false|false||At dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Microbiology Diagnostic Service Section ID|Finding|false|false||Microbiology
null|Microbiological|Finding|false|false||Microbiology
null|Microbiology - Laboratory Class|Finding|false|false||Microbiologynull|Microbiology procedure|Procedure|false|false||Microbiologynull|Science of Microbiology|Title|false|false||Microbiologynull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Pathology processes|Finding|false|false||Pathology
null|Pathological aspects|Finding|false|false||Pathologynull|Pathology procedure|Procedure|false|false||Pathologynull|Pathology|Title|false|false||Pathologynull|Consent Type - Liver Biopsy|Procedure|false|false||Liver biopsy
null|Biopsy of liver (procedure)|Procedure|false|false||Liver biopsynull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|Core needle biopsy|Procedure|false|false||core needle biopsynull|Core Specimen|Finding|false|false||corenull|viral nucleocapsid location|Anatomy|false|false||corenull|Processor Core|Device|false|false||core
null|Core Device|Device|false|false||corenull|Core|Modifier|false|false||corenull|Consent Type - Needle Biopsy|Procedure|false|false||needle biopsy
null|Puncture biopsy|Procedure|false|false||needle biopsy
null|Needle biopsy (procedure)|Procedure|false|false||needle biopsynull|null|Finding|false|false||needlenull|Needle device|Device|false|false||needlenull|Needle Shape|Modifier|false|false||needlenull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Adenocarcinoma|Disorder|false|false||Adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||Adenocarcinomanull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|immunohistochemical stains|Drug|false|false||Immunohistochemical stainsnull|immunohistochemical stains procedure|Procedure|false|false||Immunohistochemical stainsnull|Stains|Drug|false|false||stainsnull|Dyes [MoA]|Finding|false|false||stainsnull|Staining method|Procedure|false|false||stainsnull|Tumor cells, uncertain whether benign or malignant|Anatomy|false|false||tumor cells
null|Tumor cells|Anatomy|false|false||tumor cellsnull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Cells|Anatomy|false|false||cellsnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|KRT20 wt Allele|Finding|false|false||CK20
null|KRT20 gene|Finding|false|false||CK20null|bicalutamide|Drug|false|false||CDX
null|cefadroxil|Drug|false|false||CDX
null|cefadroxil|Drug|false|false||CDX
null|bicalutamide|Drug|false|false||CDXnull|Cell Line-Derived Xenograft|Finding|false|false||CDXnull|Companion Diagnostic Test|Procedure|false|false||CDXnull|Negative for CK7 and TTF-1|Lab|false|false||negative for CK7 and TTF-1null|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|KRT7 wt Allele|Finding|false|false||CK7
null|KRT7 gene|Finding|false|false||CK7null|thyroid transcription factor 1|Drug|false|false||TTF-1
null|thyroid transcription factor 1|Drug|false|false||TTF-1
null|NKX2-1 protein, human|Drug|false|false||TTF-1
null|NKX2-1 protein, human|Drug|false|false||TTF-1
null|TTF1 protein, human|Drug|false|false||TTF-1
null|TTF1 protein, human|Drug|false|false||TTF-1null|NKX2-1 wt Allele|Finding|false|false||TTF-1
null|TTF1 wt Allele|Finding|false|false||TTF-1
null|NKX2-1 gene|Finding|false|false||TTF-1null|RHOH wt Allele|Finding|false|false||TTF
null|RHOH gene|Finding|false|false||TTFnull|Tumour treating fields therapy|Procedure|false|false||TTFnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Neoplasm Metastasis|Disorder|false|false||metastasis
null|Metastatic malignant neoplasm|Disorder|false|false||metastasisnull|Metastasis|Finding|false|false||metastasis
null|Metastatic Lesion|Finding|false|false||metastasisnull|Colorectal|Modifier|false|false||colorectalnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus Tachycardia|Disorder|false|false||Sinus tachycardianull|continuous electrocardiogram sinus tachycardia|Finding|false|false||Sinus tachycardia
null|Sinus Tachycardia by ECG Finding|Finding|false|false||Sinus tachycardianull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinusnull|pathologic fistula|Disorder|false|false||Sinusnull|Sinus - general anatomical term|Anatomy|false|false||Sinus
null|Nasal sinus|Anatomy|false|false||Sinusnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Voltage|LabModifier|false|false||voltagenull|Diffuse|Modifier|false|false||Diffusenull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|More|LabModifier|false|false||morenull|Prominent|Modifier|false|false||prominentnull|portable x-ray of chest|Procedure|false|false||Portable CXRnull|Portable|Modifier|false|false||Portablenull|Plain chest X-ray|Procedure|false|false||CXRnull|Secondary malignant neoplasm of lung|Disorder|false|false||pulmonary metastasesnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Possible|Finding|false|false||Possiblenull|Possible diagnosis|Modifier|false|false||Possible
null|Possibly Related to Intervention|Modifier|false|false||Possiblenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Congestion|Finding|false|false||congestionnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Lung Volumes|Finding|false|false||lung volumesnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Volume|LabModifier|false|false||volumesnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Central brand of multivitamin with minerals|Drug|true|false||central
null|Central brand of multivitamin with minerals|Drug|true|false||centralnull|Central Minus|Procedure|true|false||centralnull|Central|Modifier|false|false||centralnull|Segmental|Modifier|false|false||segmentalnull|Filling defect|Finding|true|false||filling defectnull|THYROID HORMONE PLASMA MEMBRANE TRANSPORT DEFECT|Disorder|true|false||defectnull|Defect|Finding|true|false||defectnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Procedure on artery|Procedure|false|false||arteriesnull|Arteries|Anatomy|false|false||arteries
null|Arterial system|Anatomy|false|false||arteriesnull|Processing type - Evaluation|Finding|false|false||Evaluationnull|Evaluation procedure|Procedure|false|false||Evaluation
null|Evaluation|Procedure|false|false||Evaluationnull|Limited a Little|Finding|false|false||slightly limitednull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Limited component (foundation metadata concept)|Finding|false|false||limited
null|Limited (extensiveness)|Finding|false|false||limitednull|Suboptimal|Modifier|false|false||suboptimalnull|Intravenous Bolus|Finding|false|false||IV bolusnull|Response Modality - Bolus|Finding|false|false||bolus
null|Bolus of ingested food|Finding|false|false||bolusnull|bolus infusion|Procedure|false|false||bolusnull|Bolus Dosing Unit|LabModifier|false|false||bolusnull|Bilateral|Modifier|false|false||bilateralnull|Multiple Pulmonary Nodules|Finding|false|false||pulmonary nodulesnull|Pulmonary (intended site)|Finding|true|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|true|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|null|Time|false|false||priornull|null|Attribute|false|false||CT studynull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Focal|Modifier|false|false||focalnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Hepatomegaly|Finding|false|false||Enlarged livernull|Enlargement procedure|Procedure|false|false||Enlargednull|Enlarged|Modifier|false|false||Enlargednull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Numerous|LabModifier|false|false||multiplenull|Lesion|Finding|false|false||lesionsnull|therapeutic suggestion|Finding|false|false||suggestion
null|suggestion|Finding|false|false||suggestionnull|Cost of Illness|Modifier|false|false||burden of diseasenull|Burden|Finding|false|false||burdennull|Disease|Disorder|false|false||diseasenull|Structure of right upper quadrant of abdomen|Anatomy|false|false||Right upper quadrantnull|RUQ - Right upper quadrant|Modifier|false|false||Right upper quadrantnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Quadrant|Modifier|false|false||quadrantnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Extensive|Modifier|false|false||Extensivenull|Diffuse|Modifier|false|false||diffusenull|Hepatic|Anatomy|false|false||hepaticnull|Metastatic malignant neoplasm|Disorder|false|false||metastatic disease
null|Metastatic Neoplasm|Disorder|false|false||metastatic disease
null|Neoplasm Metastasis|Disorder|false|false||metastatic diseasenull|Metastatic Lesion|Finding|false|false||metastatic diseasenull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Disease|Disorder|false|false||diseasenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Bile duct structure|Anatomy|false|false||biliary ductnull|Biliary|Finding|false|false||biliarynull|Duct (organ) structure|Anatomy|false|false||duct
null|canal [body parts]|Anatomy|false|false||ductnull|Duct Device|Device|false|false||ductnull|Obstruction|Finding|false|false||obstructionnull|portable x-ray of chest|Procedure|false|false||Portable CXRnull|Portable|Modifier|false|false||Portablenull|Plain chest X-ray|Procedure|false|false||CXRnull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Lung Volumes|Finding|false|false||lung volumesnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Volume|LabModifier|false|false||volumesnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Pulmonary vascular congestion|Disorder|false|false||pulmonary vascular congestionnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Congestion|Finding|false|false||congestionnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Small|LabModifier|false|false||smallnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Fissural|Modifier|false|false||fissuralnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|false|false||newnull|Focal|Modifier|false|false||focalnull|Abnormally opaque structure (morphologic abnormality)|Finding|true|false||opacities
null|Decreased translucency|Finding|true|false||opacitiesnull|Pneumonia|Disorder|false|false||pneumonianull|CAT scan of head|Procedure|false|false||head CTnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Process Pharmacologic Substance|Drug|true|false||processnull|Process (qualifier value)|Finding|true|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|true|false||processnull|Mass of body structure|Finding|true|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false||mass
null|null|Finding|true|false||mass
null|FBN1 wt Allele|Finding|true|false||mass
null|FBN1 gene|Finding|true|false||mass
null|Mass of body region|Finding|true|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|More|LabModifier|false|false||morenull|Sensitive|Finding|false|false||sensitivenull|stimulus sensitivity|Modifier|false|false||sensitivenull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Left hip region structure|Anatomy|false|false||Left hipnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Definite|Modifier|false|false||definite
null|Definitely Related to Intervention|Modifier|false|false||definitenull|Lytic lesion|Finding|true|false||lytic lesion
null|null|Finding|true|false||lytic lesionnull|Lysis|Finding|false|false||lyticnull|Lytic|Modifier|false|false||lyticnull|Lesion|Finding|true|false||lesion
null|null|Finding|true|false||lesionnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Bone Tissue, Human|Anatomy|false|false||osseous
null|Skeletal bone|Anatomy|false|false||osseousnull|Lesion|Finding|false|false||lesion
null|null|Finding|false|false||lesionnull|Portable|Modifier|false|false||Portablenull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Plain x-ray|Procedure|false|false||Radiographsnull|Abdominopelvic structure|Anatomy|false|false||abdomen and pelvisnull|Abdomen|Anatomy|false|false||abdomen andnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Malignant neoplasm of pelvis|Disorder|false|false||pelvisnull|Pelvis problem|Finding|false|false||pelvisnull|Pelvis+|Anatomy|false|false||pelvis
null|Pelvic cavity structure|Anatomy|false|false||pelvis
null|Pelvis|Anatomy|false|false||pelvisnull|Intestines|Anatomy|false|false||bowelnull|Gas - SpecimenType|Drug|false|false||gas
null|Gases|Drug|false|false||gas
null|Gas Dosage Form|Drug|false|false||gasnull|Gas - Specimen Source Codes|Finding|false|false||gas
null|gastrointestinal gas|Finding|false|false||gas
null|PAGR1 wt Allele|Finding|false|false||gas
null|GALNS wt Allele|Finding|false|false||gas
null|GALNS gene|Finding|false|false||gas
null|GAST wt Allele|Finding|false|false||gas
null|GAST gene|Finding|false|false||gas
null|germacrene-A synthase activity|Finding|false|false||gas
null|PAGR1 gene|Finding|false|false||gasnull|Patterns|Modifier|false|false||patternnull|Living Arrangement - Relative|Finding|false|false||relativenull|null|Attribute|false|false||relativenull|Relative (related person)|Subject|false|false||relativenull|Relative|Modifier|false|false||relativenull|Intestines|Anatomy|false|false||bowelnull|Gas - SpecimenType|Drug|false|false||gas
null|Gases|Drug|false|false||gas
null|Gas Dosage Form|Drug|false|false||gasnull|Gas - Specimen Source Codes|Finding|false|false||gas
null|gastrointestinal gas|Finding|false|false||gas
null|PAGR1 wt Allele|Finding|false|false||gas
null|GALNS wt Allele|Finding|false|false||gas
null|GALNS gene|Finding|false|false||gas
null|GAST wt Allele|Finding|false|false||gas
null|GAST gene|Finding|false|false||gas
null|germacrene-A synthase activity|Finding|false|false||gas
null|PAGR1 gene|Finding|false|false||gasnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Structure of mid abdomen (surface region)|Anatomy|false|false||mid abdomennull|Middle|Modifier|false|false||midnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Marked|Modifier|false|false||marked
null|Massive|Modifier|false|false||markednull|Enlargement (morphologic abnormality)|Disorder|false|false||enlargementnull|Hypertrophy|Finding|false|false||enlargementnull|Enlargement procedure|Procedure|false|false||enlargementnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||loopsnull|Special Handling Code - Upright|Finding|false|false||uprightnull|Entity Handling - upright|Phenomenon|false|false||uprightnull|Upright|Modifier|false|false||uprightnull|View|Modifier|false|false||viewnull|Suboptimal|Modifier|false|false||suboptimalnull|Limited (extensiveness)|Finding|false|false||limitsnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Intraperitoneal Route of Administration|Finding|false|false||intraperitoneal
null|Intraperitoneal (intended site)|Finding|false|false||intraperitonealnull|Intraperitoneal|Modifier|false|false||intraperitonealnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Free of (attribute)|Finding|false|false||freenull|Empty (qualifier)|Modifier|false|false||freenull|Intraperitoneal Route of Administration|Finding|false|false||intraperitoneal
null|Intraperitoneal (intended site)|Finding|false|false||intraperitonealnull|Intraperitoneal|Modifier|false|false||intraperitonealnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Left lateral decubitus position|Modifier|false|false||left lateral decubitusnull|Lateral to the left|Modifier|false|false||left lateralnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lateral|Modifier|false|false||lateralnull|Pressure injury|Disorder|false|false||decubitusnull|Decubitus direction|Modifier|false|false||decubitusnull|View|Modifier|false|false||viewnull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Metastatic malignant neoplasm|Disorder|false|false||metastatic cancer
null|Disseminated Malignant Neoplasm|Disorder|false|false||metastatic cancer
null|Neoplasm Metastasis|Disorder|false|false||metastatic cancernull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Lesion|Finding|false|false||lesionsnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Lung|Anatomy|false|false||lungsnull|Initially|Time|false|false||initiallynull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Intrapulmonary Route of Administration|Finding|false|false||intrapulmonarynull|Intrapulmonary|Modifier|false|false||intrapulmonarynull|Tumor Burden|Procedure|false|false||tumor burdennull|Neoplasms|Disorder|false|false||tumornull|Tumor Mass|Finding|false|false||tumor
null|null|Finding|false|false||tumornull|Burden|Finding|false|false||burdennull|Late|Time|false|false||laternull|Percutaneous Route of Drug Administration|Finding|false|false||percutaneousnull|Percutaneous|Modifier|false|false||percutaneousnull|Consent Type - Liver Biopsy|Procedure|false|false||liver biopsy
null|Biopsy of liver (procedure)|Procedure|false|false||liver biopsynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|oncology services|Procedure|false|false||oncology servicenull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Adenocarcinoma of colon metastatic|Disorder|false|false||Metastatic colon adenocarcinomanull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Adenocarcinoma of colon|Disorder|false|false||colon adenocarcinomanull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|null|Finding|false|false||embolus
null|Embolus|Finding|false|false||embolusnull|Structure of right upper quadrant of abdomen|Anatomy|false|false||right upper quadrantnull|RUQ - Right upper quadrant|Modifier|false|false||right upper quadrantnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Quadrant|Modifier|false|false||quadrantnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|unknown vaccine or immune globulin|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|Unknown - Vaccines administered|Drug|false|false||unknown
null|unknown vaccine or immune globulin|Drug|false|false||unknownnull|Unknown - mode of arrival code|Finding|false|false||unknown
null|Unknown - Special Program Code|Finding|false|false||unknown
null|Unknown - Production Class Code|Finding|false|false||unknown
null|Unknown - Patient Outcome|Finding|false|false||unknown
null|Unknown - Recreational Drug Use Code|Finding|false|false||unknown
null|Unknown - Escort Required|Finding|false|false||unknown
null|Unknown - Transport Arranged|Finding|false|false||unknown
null|Unknown - Living Arrangement|Finding|false|false||unknown
null|Unknown - Employment Status|Finding|false|false||unknown
null|Unknown - Relationship|Finding|false|false||unknown
null|Unknown - publishing section|Finding|false|false||unknown
null|Unknown Publicity Code|Finding|false|false||unknown
null|Unknown - Event reason|Finding|false|false||unknown
null|Unknown - Religion|Finding|false|false||unknown
null|Unknown - Organ Donor Code|Finding|false|false||unknown
null|unknown - NullFlavor|Finding|false|false||unknown
null|Unknown - Notify Clergy Code|Finding|false|false||unknown
null|Unknown - Administrative Gender|Finding|false|false||unknown
null|Unknown - Patient Condition Code|Finding|false|false||unknown
null|Unknown - Living Will Code|Finding|false|false||unknown
null|Marital Status - Unknown|Finding|false|false||unknown
null|Unknown - Patient Class|Finding|false|false||unknown
null|Unknown - Event Expected|Finding|false|false||unknown
null|Unknown - Expanded yes/no indicator|Finding|false|false||unknown
null|Unknown - Immunization Registry Status|Finding|false|false||unknown
null|Unknown - Container status|Finding|false|false||unknown
null|Unknown - CWE statuses|Finding|false|false||unknown
null|Unknown - Patient_s Relationship to Insured|Finding|false|false||unknown
null|Unknown - Job Status|Finding|false|false||unknown
null|Unknown - Precaution Code|Finding|false|false||unknown
null|Unknown - Contact Role|Finding|false|false||unknown
null|Unknown - Living Dependency|Finding|false|false||unknownnull|Ethnic group unknown|Subject|false|false||unknownnull|Unknown - Allergy Severity|Modifier|false|false||unknown
null|Unknown - HL7 update mode|Modifier|false|false||unknown
null|Unknown|Modifier|false|false||unknownnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Lung|Anatomy|false|false||lungsnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Patient Class - Outpatient|Finding|false|false||outpatient
null|Referral category - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Reluctance|Finding|false|false||reluctancenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Percutaneous liver biopsy|Procedure|false|false||Percutaneous liver biopsynull|Percutaneous Route of Drug Administration|Finding|false|false||Percutaneousnull|Percutaneous|Modifier|false|false||Percutaneousnull|Consent Type - Liver Biopsy|Procedure|false|false||liver biopsy
null|Biopsy of liver (procedure)|Procedure|false|false||liver biopsynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Adenocarcinoma of colon|Disorder|false|false||colonic adenocarcinomanull|Colon structure (body structure)|Anatomy|false|false||colonicnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Following|Time|false|false||Following
null|Status post|Time|false|false||Followingnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|Provider|Finding|false|false||providersnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|oncology services|Procedure|false|false||oncology servicenull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Potential|Modifier|false|false||potentialnull|Clinical Trials|Procedure|false|false||trialnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Very Poor|Finding|false|false||very poornull|Very|Modifier|false|false||verynull|Patient Condition Code - Poor|Finding|false|false||poor
null|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Functional Relationship|Finding|false|false||functional
null|Function (attribute)|Finding|false|false||functional
null|Functional|Finding|false|false||functionalnull|Nutritional status|Finding|false|false||nutritional statusnull|null|Attribute|false|false||nutritionalnull|Nutritional|Modifier|false|false||nutritionalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Goals of Care|Procedure|false|false||goals of carenull|What subject filter - Goals|Finding|false|false||goals
null|objective (goal)|Finding|false|false||goals
null|treatment goals|Finding|false|false||goalsnull|null|Attribute|false|false||goalsnull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|Goals of Care|Procedure|false|false||goals of carenull|What subject filter - Goals|Finding|false|false||goals
null|objective (goal)|Finding|false|false||goals
null|treatment goals|Finding|false|false||goalsnull|null|Attribute|false|false||goalsnull|care of - AddressPartType|Finding|false|false||care ofnull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfort
null|Comfort brand of hydroxyethyl cellulose|Drug|false|false||comfortnull|Comfort|Finding|false|false||comfortnull|Symptom Management|Procedure|false|false||symptom management
null|Palliative Care|Procedure|false|false||symptom managementnull|Symptoms|Finding|false|false||symptomnull|null|Attribute|false|false||symptomnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Home Hospice|Procedure|false|false||home hospicenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Structure of left thigh|Anatomy|false|false||Left thighnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|thigh weakness|Finding|false|false||thigh weaknessnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Focal|Modifier|false|false||focalnull|Structure of left thigh|Anatomy|false|false||left thighnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|thigh weakness|Finding|false|false||thigh weaknessnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Relationship by association|Finding|false|false||association
null|Mental association|Finding|false|false||association
null|NCI Thesaurus Association|Finding|false|false||association
null|Association Class|Finding|false|false||associationnull|Chemical Association|Phenomenon|false|false||associationnull|Relationships|Modifier|false|false||associationnull|Diffuse|Modifier|false|false||diffusenull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Chronicity|Time|false|false||chronicitynull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Rectal Dosage Form|Drug|false|false||rectalnull|Rectal Route of Administration|Finding|false|false||rectal
null|Rectal (intended site)|Finding|false|false||rectalnull|TUBE,RECTAL,24FR,PLASTIC B#6510|Device|false|false||rectalnull|rectal|Modifier|false|false||rectalnull|Numbness of saddle area|Finding|true|false||saddle anesthesianull|Anesthesia substance|Drug|true|false||anesthesianull|null|Finding|true|false||anesthesia
null|Absence of sensation|Finding|true|false||anesthesianull|Anesthesia procedures|Procedure|true|false||anesthesia
null|Dental anesthesia|Procedure|true|false||anesthesianull|null|Attribute|true|false||anesthesianull|incontinent of urine on urethra exam|Finding|false|false||incontinent of urine
null|Urinary Incontinence|Finding|false|false||incontinent of urinenull|Incontinent|Finding|false|false||incontinentnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Feces|Finding|false|false||fecesnull|Underlying|Finding|false|false||underlyingnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Concern|Finding|false|false||concernnull|Metastatic malignant neoplasm to bone|Disorder|false|false||bony metastasesnull|Bony|Finding|false|false||bonynull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Cone-Rod Dystrophy 2|Disorder|false|false||cordnull|Cord - Body Parts|Anatomy|false|false||cordnull|Cord Device|Device|false|false||cordnull|Involvement with|Finding|false|false||involvementnull|Alternative|Modifier|false|false||alternativenull|Consideration|Finding|false|false||considerationnull|Epidural Route of Administration|Finding|false|false||epiduralnull|null|Procedure|false|false||epiduralnull|Body Parts - Epidural|Anatomy|false|false||epiduralnull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Living Arrangement - Transient|Finding|false|false||transient
null|Encounter due to vagabond status|Finding|false|false||transientnull|Transient Population Group|Subject|false|false||transientnull|Transitory|Time|false|false||transientnull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|Empiric|Modifier|false|false||empiricnull|Antibiotics|Drug|false|false||antibioticnull|coverage - HL7PublishingDomain|Finding|false|false||coverage
null|null|Finding|false|false||coverage
null|coverage - financial contract|Finding|false|false||coveragenull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|cefepime|Drug|false|false||cefepim
null|cefepime|Drug|false|false||cefepimnull|Frequently|Time|false|false||frequentnull|Numerous|LabModifier|false|false||multiplenull|Lumbosacral|Modifier|false|false||lumbosacralnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|lorazepam|Drug|false|false||lorazepam
null|lorazepam|Drug|false|false||lorazepamnull|Premedication|Procedure|false|false||premedicationnull|Claustrophobia|Disorder|false|false||claustrophobianull|Neurologic Examination|Procedure|false|false||Neuro examnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Abdominal Pain|Finding|false|false||Abdominal painnull|Abdomen|Anatomy|false|false||Abdominalnull|Abdominal (qualifier value)|Modifier|false|false||Abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Intermittent abdominal pain|Finding|false|false||intermittent abdominal painnull|Intermittent|Time|false|false||intermittentnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|peritoneal|Anatomy|false|false||peritoneal
null|Peritoneum|Anatomy|false|false||peritonealnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Obstruction|Finding|false|false||obstructionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Abdominal Cavity|Anatomy|false|false||intraabdominalnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Episode of|Time|false|false||episodesnull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Hematemesis|Finding|false|false||hematemesisnull|Numerous|LabModifier|false|false||multiplenull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Obstruction|Finding|true|false||obstructionnull|CT of abdomen|Procedure|false|false||CT abdomennull|null|Attribute|false|false||CT abdomennull|Malignant neoplasm of abdomen|Disorder|false|false||abdomennull|Abdomen problem|Finding|false|false||abdomennull|Abdomen|Anatomy|false|false||abdomen
null|Abdominal Cavity|Anatomy|false|false||abdomennull|Alternative|Modifier|false|false||alternativenull|Source|Finding|false|false||sourcesnull|Abdominal Cavity|Anatomy|false|false||intraabdominalnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Numerous|LabModifier|false|false||multiplenull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Hematemesis|Finding|false|false||Hematemesisnull|Single episode|Time|false|false||single episodenull|Marital Status - Single|Finding|false|false||single
null|Unmarried|Finding|false|false||singlenull|Singular|LabModifier|false|false||singlenull|Episode of|Time|false|false||episode ofnull|Episode of|Time|false|false||episodenull|Small|LabModifier|false|false||smallnull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Approximate|Modifier|false|false||approximatelynull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|pantoprazole|Drug|false|false||pantoprazole
null|pantoprazole|Drug|false|false||pantoprazolenull|Gastrointestinal attachment|Finding|false|false||gastrointestinalnull|gastrointestinal|Modifier|false|false||gastrointestinalnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Following|Time|false|false||subsequentnull|Discontinuation (procedure)|Finding|false|false||discontinuation
null|Discontinued|Finding|false|false||discontinuationnull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|Recurrent Malignant Neoplasm|Disorder|true|false||recurrencenull|Recurrence (disease attribute)|Finding|true|false||recurrencenull|Recurrence|Phenomenon|true|false||recurrencenull|Equivocal|Modifier|false|false||questionablenull|First episode|Time|false|false||first episodenull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Episode of|Time|false|false||episodenull|True|Modifier|false|false||truenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Popsicle|Drug|false|false||popsiclenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Esophagogastroduodenoscopy|Procedure|false|false||Esophagogastroduodenoscopynull|Absent|Finding|false|false||absence ofnull|Absence (morphologic abnormality)|Disorder|false|false||absencenull|Absent|Finding|false|false||absencenull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Hematemesis|Finding|false|false||hematemesisnull|null|Time|false|false||priornull|Esophagogastroduodenoscopy|Procedure|true|false||EGDsnull|Esophagogastroduodenoscopes|Device|true|false||EGDsnull|Availability of|Finding|false|false||availablenull|ATP5F1A gene|Finding|false|false||OMRnull|Mental state|Finding|false|false||mental statusnull|null|Attribute|false|false||mental status
null|null|Attribute|false|false||mental statusnull|Psyche structure|Finding|false|false||mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Infrequent|Time|false|false||occasionalnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|LITAF gene|Finding|false|false||simplenull|Simple|Modifier|false|false||simplenull|Uncertainty|Finding|false|false||uncertainnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Communicable Diseases|Disorder|false|false||Infectiousnull|infectious - Entity Risk|Modifier|false|false||Infectiousnull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Culture (Anthropological)|Finding|false|false||culturesnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Following|Time|false|false||subsequentnull|CAT scan of head|Procedure|false|false||head CTnull|Problems with head|Disorder|false|false||headnull|Procedure on head|Procedure|false|false||headnull|Structure of head of caudate nucleus|Anatomy|false|false||head
null|Head|Anatomy|false|false||headnull|Head Device|Device|false|false||headnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Intracranial Route of Administration|Finding|false|false||intracranialnull|Intracranial|Anatomy|false|false||intracranialnull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Nuclear magnetic resonance imaging brain|Procedure|false|false||Brain MRInull|Brain Diseases|Disorder|false|false||Brainnull|Head>Brain|Anatomy|false|false||Brain
null|Brain|Anatomy|false|false||Brainnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Definitive|Time|false|false||definitivenull|Exclusion Criteria|Finding|false|false||exclusionnull|Exclusion|Event|false|false||exclusionnull|Metastatic malignant neoplasm|Disorder|false|false||metastases
null|Neoplasm Metastasis|Disorder|false|false||metastasesnull|Metastatic Lesion|Finding|false|false||metastasesnull|Claustrophobia|Disorder|false|false||claustrophobianull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Aversion|Drug|false|false||aversion
null|Aversion|Drug|false|false||aversionnull|Aversion (finding)|Finding|false|false||aversionnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|A1BG gene|Finding|false|false||ABGnull|Analysis of arterial blood gases and pH|Procedure|false|false||ABGnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hypercapnia|Finding|false|false||CO2 retentionnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|Retention of content|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Urinary Retention|Finding|false|false||retention
null|cellular entity retention|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiates|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiates
null|Opiate Alkaloids|Drug|false|false||opiatesnull|Opiate Measurement|Procedure|false|false||opiatesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Drowsiness|Finding|false|false||sleepynull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Mathematical Factor|Finding|false|false||factor
null|Factor|Finding|false|false||factor
null|Feelings about Genomic Testing Results|Finding|false|false||factornull|Hepatic Encephalopathy|Disorder|false|false||Hepatic encephalopathynull|Hepatic|Anatomy|false|false||Hepaticnull|Encephalopathies|Disorder|false|false||encephalopathynull|Amount type - Differential|Finding|false|false||differentialnull|Differential (qualifier value)|Modifier|false|false||differential
null|Different|Modifier|false|false||differential
null|Differential - view|Modifier|false|false||differentialnull|metastatic qualifier|Finding|false|false||metastatic
null|Metastatic to|Finding|false|false||metastaticnull|Lesion|Finding|false|false||lesionsnull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Asterixis|Finding|false|false||asterixisnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|ABLEPHARON-MACROSTOMIA SYNDROME|Disorder|false|false||AMSnull|TWIST2 wt Allele|Finding|false|false||AMSnull|Accelerator Mass Spectrometry|Procedure|false|false||AMSnull|Severe depression|Disorder|false|false||severe depressionnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Mental state|Finding|false|false||Mental statusnull|null|Attribute|false|false||Mental status
null|null|Attribute|false|false||Mental statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|On discharge|Time|false|false||on dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|Sudden onset (contextual qualifier) (qualifier value)|Finding|false|false||acute onsetnull|Sudden onset (attribute)|Time|false|false||acute onset
null|acute|Time|false|false||acute onsetnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Onset of (contextual qualifier)|Modifier|false|false||onsetnull|Age of Onset|LabModifier|false|false||onsetnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Immune thrombocytopenic purpura|Disorder|false|false||franknull|Hypoxia, CTCAE|Finding|true|false||hypoxia
null|Hypoxia|Finding|true|false||hypoxianull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Pulmonary Embolism|Finding|false|false||pulmonary embolusnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|null|Finding|true|false||embolus
null|Embolus|Finding|true|false||embolusnull|clotrimazole|Drug|false|false||clot
null|clotrimazole|Drug|false|false||clotnull|Blood Clot|Finding|false|false||clotnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Focal|Modifier|false|false||focalnull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Cardiac enzymes|Drug|false|false||cardiac enzymes
null|Cardiac enzymes|Drug|false|false||cardiac enzymesnull|Cardiac enzymes/isoenzymes measurement|Procedure|false|false||cardiac enzymesnull|null|Attribute|false|false||cardiac enzymesnull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes, peripheral vasodilators|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|Enzymes, antithrombotic|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes, hematological|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymes
null|Enzymes for ALIMENTARY TRACT AND METABOLISM|Drug|false|false||enzymesnull|enzymology|Finding|false|false||enzymesnull|Acute Coronary Syndrome|Disorder|false|false||acute coronary syndromenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Heart|Anatomy|false|false||coronarynull|Coronary|Modifier|false|false||coronarynull|Syndrome|Disorder|false|false||syndromenull|IPSS-R Risk Category Low|Finding|false|false||Low
null|IPSS Risk Category Low|Finding|false|false||Low
null|low confidentiality|Finding|false|false||Lownull|Low - MessageWaitingPriority|Modifier|false|false||Low
null|low|Modifier|false|false||Low
null|low exposure|Modifier|false|false||Lownull|null|LabModifier|false|false||Lownull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Consistent with|Finding|false|false||consistentnull|null|Time|false|false||priornull|Limited component (foundation metadata concept)|Finding|false|false||limited
null|Limited (extensiveness)|Finding|false|false||limitednull|Suspicion|Finding|false|false||suspicionnull|Pericardial effusion|Disorder|false|false||pericardial effusionnull|Pericardial effusion body substance|Finding|false|false||pericardial effusionnull|Pericardial (qualifier value)|Anatomy|false|false||pericardial
null|Pericardial sac structure|Anatomy|false|false||pericardialnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Dyspnea|Finding|false|false||Shortness of breathnull|null|Attribute|false|false||Shortness of breathnull|Breath|Finding|false|false||breathnull|Course|Time|false|false||coursenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Exception - Property or Attribute|Finding|false|false||exception
null|exception - ResponseLevel|Finding|false|false||exceptionnull|nebulizers (medication)|Drug|false|false||nebulizersnull|Nebulizers|Device|false|false||nebulizersnull|Expectorants|Drug|false|false||expectorantsnull|Poisoning by, adverse effect of and underdosing of expectorants|Disorder|false|false||expectorants
null|Poisoning by expectorant|Disorder|false|false||expectorants
null|Expectorants causing adverse effects in therapeutic use|Disorder|false|false||expectorantsnull|Leukocytosis|Disorder|false|false||Leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||Leukocytosisnull|White Blood Cell Count procedure|Procedure|false|false||White blood cell countnull|null|Lab|false|false||White blood cell countnull|Leukocytes|Anatomy|false|false||White blood cellnull|White (population group)|Subject|false|false||White
null|Caucasian|Subject|false|false||White
null|Caucasians|Subject|false|false||Whitenull|White color|Modifier|false|false||Whitenull|Blood Cell Count|Procedure|false|false||blood cell count
null|Complete Blood Count|Procedure|false|false||blood cell countnull|Blood Cells|Anatomy|false|false||blood cellnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Cell Count|Procedure|false|false||cell countnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Peak level|Modifier|false|false||peakednull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Recent|Time|false|false||recentnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Work-up|Procedure|false|false||work upnull|Work|Event|false|false||worknull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|Blood culture|Procedure|false|false||blood culturesnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|Apyrexial|Finding|false|false||afebrilenull|Exception - Property or Attribute|Finding|false|false||exception
null|exception - ResponseLevel|Finding|false|false||exceptionnull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|Encounter due to vagabond status|Finding|false|false||transient
null|Living Arrangement - Transient|Finding|false|false||transientnull|Transient Population Group|Subject|false|false||transientnull|Transitory|Time|false|false||transientnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Liver Function Tests|Procedure|false|false||Liver function testnull|Liver function|Finding|false|false||Liver functionnull|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|liver extract|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Liver
null|Liver brand of Vitamin B 12|Drug|false|false||Livernull|Benign neoplasm of liver|Disorder|false|false||Liver
null|Liver diseases|Disorder|false|false||Livernull|Liver problem|Finding|false|false||Livernull|Procedures on liver|Procedure|false|false||Livernull|Abdomen>Liver|Anatomy|false|false||Liver
null|null|Anatomy|false|false||Liver
null|Liver|Anatomy|false|false||Livernull|Function Test|Procedure|false|false||function testnull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Tests (qualifier value)|Finding|false|false||test
null|Testing|Finding|false|false||testnull|Laboratory Procedures|Procedure|false|false||testnull|Test - temporal region|Anatomy|false|false||testnull|Test Result|Lab|false|false||testnull|Test Dosing Unit|LabModifier|false|false||testnull|Congenital Abnormality|Disorder|false|false||abnormalitiesnull|teratologic|Finding|false|false||abnormalitiesnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|Aspartate Transaminase|Drug|false|false||AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||AST
null|SLC17A5 protein, human|Drug|false|false||ASTnull|Atypical Spitz Nevus|Disorder|false|false||ASTnull|SLC17A5 wt Allele|Finding|false|false||AST
null|SLC17A5 gene|Finding|false|false||AST
null|GOT1 gene|Finding|false|false||ASTnull|Asterion|Anatomy|false|false||ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alkaline Phosphatase|Drug|false|false||alkaline phosphatase
null|Alkaline Phosphatase|Drug|false|false||alkaline phosphatasenull|Alkaline phosphatase metabolic function|Finding|false|false||alkaline phosphatasenull|Alkaline phosphatase measurement|Procedure|false|false||alkaline phosphatasenull|Phosphoric Monoester Hydrolases|Drug|false|false||phosphatase
null|Phosphoric Monoester Hydrolases|Drug|false|false||phosphatasenull|phosphoric monoester hydrolase activity|Finding|false|false||phosphatasenull|Phosphatase (disposition)|Modifier|false|false||phosphatasenull|Bilirubin|Drug|false|false||total bilirubin
null|Bilirubin|Drug|false|false||total bilirubinnull|Total bilirubin metabolic function|Finding|false|false||total bilirubinnull|Bilirubin, total measurement|Procedure|false|false||total bilirubinnull|Total bilirubin level|Lab|false|false||total bilirubinnull|Total|Modifier|false|false||totalnull|bilirubin preparation|Drug|false|false||bilirubin
null|bilirubin preparation|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubin
null|Bilirubin|Drug|false|false||bilirubinnull|Bilirubin, total measurement|Procedure|false|false||bilirubin
null|blood bilirubin level test|Procedure|false|false||bilirubinnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hepatic|Anatomy|false|false||hepaticnull|Infiltration Route of Administration|Finding|false|false||infiltration
null|Infiltration|Finding|false|false||infiltration
null|Spread by direct extension|Finding|false|false||infiltrationnull|Infiltration (procedure)|Procedure|false|false||infiltrationnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Structure of right upper quadrant of abdomen|Anatomy|false|false||Right upper quadrantnull|RUQ - Right upper quadrant|Modifier|false|false||Right upper quadrantnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Upper Surface|Modifier|false|false||upper
null|Upper|Modifier|false|false||uppernull|Quadrant|Modifier|false|false||quadrantnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Cholecystitis|Disorder|false|false||cholecystitisnull|Obstructed|Finding|false|false||obstructivenull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Abdominal Cavity|Anatomy|false|false||intraabdominalnull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Elevated lactate level|Finding|false|false||Elevated lactatenull|Elevated|Modifier|false|false||Elevated
null|High|Modifier|false|false||Elevatednull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Copious|Finding|false|false||copiousnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Reflecting|Finding|false|false||reflectingnull|Hepatic|Anatomy|false|false||hepaticnull|Clearance procedure|Procedure|false|false||clearancenull|Clearance of substance|Attribute|false|false||clearancenull|Clearance [PK]|Phenomenon|false|false||clearancenull|Clearance|Modifier|false|false||clearancenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Malignant (qualifier value)|Modifier|false|false||malignantnull|Infiltration Route of Administration|Finding|false|false||infiltration
null|Infiltration|Finding|false|false||infiltration
null|Spread by direct extension|Finding|false|false||infiltrationnull|Infiltration (procedure)|Procedure|false|false||infiltrationnull|Sinus Tachycardia|Disorder|false|false||Sinus tachycardianull|continuous electrocardiogram sinus tachycardia|Finding|false|false||Sinus tachycardia
null|Sinus Tachycardia by ECG Finding|Finding|false|false||Sinus tachycardianull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinusnull|pathologic fistula|Disorder|false|false||Sinusnull|Sinus - general anatomical term|Anatomy|false|false||Sinus
null|Nasal sinus|Anatomy|false|false||Sinusnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|persistently|Finding|false|false||persistentlynull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Responsive|Finding|false|false||responsivenull|Copious|Finding|false|false||copiousnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Tachycardia by ECG Finding|Finding|false|false||Tachycardia
null|Tachycardia|Finding|false|false||Tachycardianull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Concurrent|Time|false|false||concurrentnull|Leukocytosis|Disorder|false|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|false|false||leukocytosisnull|Elevated lactate level|Finding|false|false||elevated lactatenull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|lactate|Drug|false|false||lactate
null|lactate|Drug|false|false||lactate
null|Lactates|Drug|false|false||lactatenull|Lactic acid measurement|Procedure|false|false||lactatenull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Source (property) (qualifier value)|Finding|false|false||source
null|Term Source|Finding|false|false||source
null|Source|Finding|false|false||sourcenull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Suspicion|Finding|false|false||suspicionnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|Pulmonary Embolism|Finding|false|false||pulmonary embolusnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|null|Finding|false|false||embolus
null|Embolus|Finding|false|false||embolusnull|Basis|Drug|false|false||basisnull|Basis - conceptual entity|Finding|false|false||basisnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Hypoxia|Finding|false|false||hypoxicnull|Hematocrit level|Finding|false|false||Hematocritnull|Hematocrit Measurement|Procedure|false|false||Hematocritnull|hematocrit attribute|Attribute|false|false||Hematocritnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|false|false||bleedingnull|Exception - Property or Attribute|Finding|false|false||exception
null|exception - ResponseLevel|Finding|false|false||exceptionnull|Living Arrangement - Transient|Finding|false|false||transient
null|Encounter due to vagabond status|Finding|false|false||transientnull|Transient Population Group|Subject|false|false||transientnull|Transitory|Time|false|false||transientnull|Hematemesis|Finding|false|false||hematemesisnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Depressed mood|Disorder|false|false||depressednull|Flat affect|Finding|false|false||flat affectnull|Residential flat|Device|false|false||flatnull|Flat shape|Modifier|false|false||flatnull|Affect (mental function)|Finding|false|false||affectnull|assessment of affect|Procedure|false|false||affectnull|Anhedonia|Disorder|false|false||anhedonianull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Underlying|Finding|false|false||underlyingnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Motivation|Finding|false|false||motivationnull|Diagnosis Classification - Diagnosis|Finding|false|false||diagnosis
null|diagnosis aspects|Finding|false|false||diagnosisnull|Diagnosis|Procedure|false|false||diagnosisnull|null|Attribute|false|false||diagnosisnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Known|Modifier|false|false||knownnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Suicidal|Disorder|true|false||suicidalnull|ideation|Finding|false|false||ideationnull|Frequently|Time|false|false||frequentlynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|sertraline|Drug|false|false||sertraline
null|sertraline|Drug|false|false||sertralinenull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Consent Type - Liver Biopsy|Procedure|false|false||liver biopsy
null|Biopsy of liver (procedure)|Procedure|false|false||liver biopsynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Explanation|Finding|false|false||explanationnull|Social Work (discipline)|Subject|false|false||social worknull|Social|Finding|false|false||socialnull|Work|Event|false|false||worknull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Hematocrit level|Finding|false|false||Hematocritnull|Hematocrit Measurement|Procedure|false|false||Hematocritnull|hematocrit attribute|Attribute|false|false||Hematocritnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Recent|Time|false|false||recentnull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Anemia of chronic disease|Disorder|false|false||anemia of chronic diseasenull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Chronic disease|Disorder|false|false||chronic diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Disease|Disorder|false|false||diseasenull|Basis|Drug|false|false||basisnull|Basis - conceptual entity|Finding|false|false||basisnull|Laboratory test finding|Lab|false|false||labsnull|Taking vital signs|Procedure|false|false||Vital signsnull|null|Attribute|false|false||Vital signs
null|Vital signs|Attribute|false|false||Vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||Vitalnull|Vital (qualifier value)|Modifier|false|false||Vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Exception - Property or Attribute|Finding|false|false||exception
null|exception - ResponseLevel|Finding|false|false||exceptionnull|Persistent|Time|false|false||persistentnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|false|false||bleedingnull|Bed Status - Isolated|Finding|false|false||isolated
null|Isolated|Finding|false|false||isolatednull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Emesis [PE]|Finding|false|false||emesis
null|Vomiting|Finding|false|false||emesis
null|Vomitus|Finding|false|false||emesisnull|Emesis <Emesidini>|Entity|false|false||emesis
null|Emesis <subgenus>|Entity|false|false||emesisnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Blood Coagulation Disorders|Disorder|false|false||Coagulopathynull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Reflecting|Finding|false|false||reflectnull|Synthesis|Event|false|false||syntheticnull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Hepatic|Anatomy|false|false||hepaticnull|Infiltration Route of Administration|Finding|false|false||infiltration
null|Infiltration|Finding|false|false||infiltration
null|Spread by direct extension|Finding|false|false||infiltrationnull|Infiltration (procedure)|Procedure|false|false||infiltrationnull|Primary malignant neoplasm|Disorder|false|false||malignancy
null|Malignant Neoplasms|Disorder|false|false||malignancynull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Oral intake|Finding|false|false||oral intakenull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Intake|Finding|false|false||intakenull|Measurement of fluid intake|Procedure|false|false||intake
null|Intake (treatment)|Procedure|false|false||intakenull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|false|false||bleedingnull|Exception - Property or Attribute|Finding|false|false||exception
null|exception - ResponseLevel|Finding|false|false||exceptionnull|Living Arrangement - Transient|Finding|false|false||transient
null|Encounter due to vagabond status|Finding|false|false||transientnull|Transient Population Group|Subject|false|false||transientnull|Transitory|Time|false|false||transientnull|Hematemesis|Finding|false|false||hematemesisnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Marketing basis - Transitional|Finding|false|false||Transitionalnull|Transitional cell morphology|Modifier|false|false||Transitionalnull|Patient Discharge|Procedure|false|false||Patient dischargenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Home Hospice|Procedure|false|false||home hospicenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Inaccurate|Modifier|false|false||inaccuratenull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||SOBnull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||DAILYnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Sedation|Finding|false|false||sedation
null|Sedated state|Finding|false|false||sedationnull|Sedation procedure|Procedure|false|false||sedationnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|bupropion|Drug|false|false||BuPROPion
null|bupropion|Drug|false|false||BuPROPionnull|Daily|Time|false|false||DAILYnull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|tramadol|Drug|false|false||TraMADOL
null|tramadol|Drug|false|false||TraMADOLnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADOLnull|Ultram|Drug|false|false||Ultram
null|Ultram|Drug|false|false||Ultramnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|sennosides, USP|Drug|false|false||sennosides
null|sennosides, USP|Drug|false|false||sennosidesnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||omeprazole
null|omeprazole|Drug|false|false||omeprazolenull|capsule (pharmacologic)|Drug|false|false||capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||capsule
null|Structure of organ capsule|Anatomy|false|false||capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||Dailynull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|Hospital bed|Device|false|false||Hospital Bednull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Hospital bed|Device|false|false||Hospital Bednull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|BORNHOLM EYE DISEASE|Disorder|false|false||Bednull|Bachelor of Education|Finding|false|false||Bednull|Beds|Device|false|false||Bednull|Patient Location - Bed|Modifier|false|false||Bednull|Therapeutic brand of coal tar|Drug|false|false||Therapeutic
null|Therapeutic brand of coal tar|Drug|false|false||Therapeuticnull|Therapeutic - Location Service Code|Finding|false|false||Therapeutic
null|Therapeutic|Finding|false|false||Therapeuticnull|Therapeutic procedure|Procedure|false|false||Therapeuticnull|Mattresses|Device|false|false||Mattressnull|Hospice Care|Procedure|false|false||Hospicenull|Hospice (environment)|Device|false|false||Hospicenull|Hospice (environment)|Entity|false|false||Hospicenull|What subject filter - Order|Finding|false|false||Order
null|Medical Order|Finding|false|false||Order
null|Order (taxonomic)|Finding|false|false||Order
null|Order (record artifact)|Finding|false|false||Order
null|Order (document)|Finding|false|false||Ordernull|Order [PK]|Phenomenon|false|false||Ordernull|Order (action)|Event|false|false||Ordernull|Order (arrangement)|Modifier|false|false||Order
null|Permutation|Modifier|false|false||Ordernull|Hospice Care|Procedure|false|false||Hospicenull|Hospice (environment)|Device|false|false||Hospicenull|Hospice (environment)|Entity|false|false||Hospicenull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||traZODONE
null|trazodone|Drug|false|false||traZODONEnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||constipationnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||Primarynull|Primary|Modifier|false|false||Primarynull|Adenocarcinoma of colon metastatic|Disorder|false|false||Metastatic colon adenocarcinomanull|metastatic qualifier|Finding|false|false||Metastatic
null|Metastatic to|Finding|false|false||Metastaticnull|Adenocarcinoma of colon|Disorder|false|false||colon adenocarcinomanull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Confusion|Disorder|false|false||Confusednull|Precaution Code - Confused|Finding|false|false||Confused
null|Clouded consciousness|Finding|false|false||Confusednull|Sometimes|Time|false|false||sometimesnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Bed-ridden|Finding|false|false||Bedboundnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Underlying|Finding|false|false||underlyingnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Pneumonia|Disorder|true|false||pneumonianull|Blood Clot|Finding|true|false||blood clot
null|Thrombus|Finding|true|false||blood clotnull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|In Blood|Finding|true|false||blood
null|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||bloodnull|clotrimazole|Drug|true|false||clot
null|clotrimazole|Drug|true|false||clotnull|Blood Clot|Finding|true|false||clotnull|Blood Vessel|Anatomy|false|false||blood vesselsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Blood Vessel|Anatomy|false|false||vesselsnull|Lung|Anatomy|false|false||lungsnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Structure of left thigh|Anatomy|false|false||left thighnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|imaging studies|Procedure|false|false||imaging studiesnull|Imaging problem|Finding|false|false||imagingnull|Diagnostic Imaging|Procedure|false|false||imaging
null|Imaging Techniques|Procedure|false|false||imagingnull|Imaging Technology|Title|false|false||imagingnull|Scientific Study|Procedure|false|false||studiesnull|Further|Modifier|false|false||furthernull|Act Class - investigation|Finding|false|false||investigationnull|Evaluation procedure|Procedure|false|false||investigation
null|Evaluation|Procedure|false|false||investigationnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Liver brand of Vitamin B 12|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|liver extract|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||liver
null|Liver brand of Vitamin B 12|Drug|false|false||livernull|Benign neoplasm of liver|Disorder|false|false||liver
null|Liver diseases|Disorder|false|false||livernull|Liver problem|Finding|false|false||livernull|Procedures on liver|Procedure|false|false||livernull|Abdomen>Liver|Anatomy|false|false||liver
null|null|Anatomy|false|false||liver
null|Liver|Anatomy|false|false||livernull|Lung|Anatomy|false|false||lungsnull|Carcinoma in situ of colon|Disorder|false|false||colon
null|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|Large Intestine|Anatomy|false|false||large bowelnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|Intestines|Anatomy|false|false||bowelnull|oncology services|Procedure|false|false||oncology servicenull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|More|LabModifier|false|false||morenull|Language Ability Proficiency - Good|Finding|false|false||good
null|Language Proficiency - Good|Finding|false|false||goodnull|Specimen Quality - Good|Modifier|false|false||good
null|Good|Modifier|false|false||goodnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Discussion (communication)|Finding|false|false||discussionnull|Discussion (procedure)|Procedure|false|false||discussionnull|Health Care|Procedure|false|false||health carenull|Health|Finding|false|false||healthnull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|Advance Directive - Proxy|Finding|false|false||proxynull|Proxy|Subject|false|false||proxynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Entity Name Part Type - family|Finding|false|false||family
null|Last Name|Finding|false|false||family
null|Living Arrangement - Family|Finding|false|false||family
null|Family (taxonomic)|Finding|false|false||family
null|Family Collection|Finding|false|false||familynull|Family|Subject|false|false||familynull|Love|Finding|false|false||lovednull|Purchased Services, Clinical and Biomedical, Home Healthcare, Hospice|Event|false|false||hospice servicesnull|Hospice Care|Procedure|false|false||hospicenull|Hospice (environment)|Device|false|false||hospicenull|Hospice (environment)|Entity|false|false||hospicenull|Clinical Service|Procedure|false|false||servicesnull|Services|Event|false|false||servicesnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions