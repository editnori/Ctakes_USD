 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|28,32
No|33,35
:|35,36
_|39,40
_|40,41
_|41,42
<EOL>|42,43
<EOL>|44,45
Admission|45,54
Date|55,59
:|59,60
_|62,63
_|63,64
_|64,65
Discharge|79,88
Date|89,93
:|93,94
_|97,98
_|98,99
_|99,100
<EOL>|100,101
<EOL>|102,103
Date|103,107
of|108,110
Birth|111,116
:|116,117
_|119,120
_|120,121
_|121,122
Sex|135,138
:|138,139
F|142,143
<EOL>|143,144
<EOL>|145,146
Service|146,153
:|153,154
NEUROLOGY|155,164
<EOL>|164,165
<EOL>|166,167
No|179,181
Known|182,187
Allergies|188,197
/|198,199
Adverse|200,207
Drug|208,212
Reactions|213,222
<EOL>|222,223
<EOL>|224,225
Attending|225,234
:|234,235
_|236,237
_|237,238
_|238,239
.|239,240
<EOL>|240,241
<EOL>|242,243
slurred|260,267
speech|268,274
<EOL>|274,275
<EOL>|276,277
Major|277,282
Surgical|283,291
or|292,294
Invasive|295,303
Procedure|304,313
:|313,314
<EOL>|314,315
None|315,319
<EOL>|319,320
<EOL>|321,322
_|350,351
_|351,352
_|352,353
year|354,358
old|359,362
right|363,368
-|368,369
handed|369,375
woman|376,381
with|382,386
hx|387,389
of|390,392
Atrial|393,399
fibrillation|400,412
on|413,415
<EOL>|416,417
Eliquis|417,424
(|425,426
only|426,430
once|431,435
daily|436,441
)|441,442
,|442,443
hypertension|444,456
,|456,457
hyperlipidemia|458,472
,|472,473
CHF|474,477
<EOL>|477,478
presents|478,486
as|487,489
transfer|490,498
from|499,503
OSH|504,507
after|508,513
she|514,517
had|518,521
acute|522,527
onset|528,533
<EOL>|534,535
dysarthria|535,545
and|546,549
CTA|550,553
showed|554,560
possible|561,569
partial|570,577
thrombus|578,586
or|587,589
stenosis|590,598
<EOL>|599,600
in|600,602
superior|603,611
division|612,620
of|621,623
L|624,625
MCA.|626,630
Transferred|631,642
here|643,647
for|648,651
closer|652,658
<EOL>|659,660
monitoring|660,670
and|671,674
possible|675,683
thrombectomy|684,696
if|697,699
her|700,703
exam|704,708
acutely|709,716
<EOL>|717,718
worsens|718,725
.|725,726
<EOL>|726,727
<EOL>|727,728
History|728,735
obtained|736,744
from|745,749
patient|750,757
and|758,761
daughter|762,770
at|771,773
bedside|774,781
.|781,782
Patient|783,790
<EOL>|791,792
is|792,794
an|795,797
excellent|798,807
historian|808,817
.|817,818
<EOL>|819,820
<EOL>|820,821
On|821,823
_|824,825
_|825,826
_|826,827
,|827,828
she|829,832
had|833,836
dinner|837,843
with|844,848
friends|849,856
and|857,860
then|861,865
returned|866,874
to|875,877
her|878,881
<EOL>|882,883
apartment|883,892
and|893,896
was|897,900
fooling|901,908
around|909,915
on|916,918
her|919,922
computer|923,931
.|931,932
Last|933,937
known|938,943
<EOL>|944,945
well|945,949
<EOL>|949,950
was|950,953
around|954,960
8|961,962
:|962,963
00|963,965
_|966,967
_|967,968
_|968,969
.|969,970
Then|971,975
,|975,976
she|977,980
had|981,984
an|985,987
odd|988,991
sensation|992,1001
and|1002,1005
started|1006,1013
<EOL>|1014,1015
throwing|1015,1023
her|1024,1027
arms|1028,1032
around|1033,1039
.|1039,1040
She|1041,1044
went|1045,1049
to|1050,1052
living|1053,1059
room|1060,1064
to|1065,1067
sit|1068,1071
down|1072,1076
<EOL>|1077,1078
and|1078,1081
<EOL>|1081,1082
tried|1082,1087
to|1088,1090
read|1091,1095
but|1096,1099
could|1100,1105
not|1106,1109
see|1110,1113
the|1114,1117
words|1118,1123
very|1124,1128
clearly|1129,1136
.|1136,1137
Then|1138,1142
,|1142,1143
<EOL>|1144,1145
two|1145,1148
family|1149,1155
members|1156,1163
were|1164,1168
knocking|1169,1177
at|1178,1180
the|1181,1184
door|1185,1189
and|1190,1193
she|1194,1197
had|1198,1201
a|1202,1203
tough|1204,1209
<EOL>|1210,1211
time|1211,1215
<EOL>|1215,1216
standing|1216,1224
up|1225,1227
to|1228,1230
open|1231,1235
door|1236,1240
.|1240,1241
She|1242,1245
was|1246,1249
able|1250,1254
to|1255,1257
eventually|1258,1268
stand|1269,1274
up|1275,1277
<EOL>|1278,1279
with|1279,1283
great|1284,1289
difficulty|1290,1300
and|1301,1304
walked|1305,1311
with|1312,1316
her|1317,1320
walker|1321,1327
.|1327,1328
She|1329,1332
usually|1333,1340
<EOL>|1341,1342
walks|1342,1347
with|1348,1352
a|1353,1354
walker|1355,1361
because|1362,1369
of|1370,1372
knee|1373,1377
replacement|1378,1389
.|1389,1390
Finally|1391,1398
,|1398,1399
got|1400,1403
up|1404,1406
<EOL>|1407,1408
out|1408,1411
of|1412,1414
chair|1415,1420
with|1421,1425
walker|1426,1432
and|1433,1436
walked|1437,1443
to|1444,1446
the|1447,1450
door|1451,1455
to|1456,1458
unlock|1459,1465
.|1465,1466
She|1467,1470
<EOL>|1471,1472
noticed|1472,1479
problems|1480,1488
talking|1489,1496
to|1497,1499
family|1500,1506
members|1507,1514
.|1514,1515
She|1516,1519
had|1520,1523
difficulty|1524,1534
<EOL>|1535,1536
forming|1536,1543
words|1544,1549
and|1550,1553
pronouncing|1554,1565
words|1566,1571
.|1571,1572
Denies|1573,1579
word|1580,1584
finding|1585,1592
<EOL>|1593,1594
difficulty|1594,1604
.|1604,1605
She|1606,1609
could|1610,1615
tell|1616,1620
it|1621,1623
was|1624,1627
slurred|1628,1635
like|1636,1640
a|1641,1642
person|1643,1649
who|1650,1653
had|1654,1657
<EOL>|1658,1659
too|1659,1662
much|1663,1667
to|1668,1670
drink|1671,1676
.|1676,1677
EMTs|1678,1682
asked|1683,1688
if|1689,1691
she|1692,1695
was|1696,1699
intoxicated|1700,1711
but|1712,1715
she|1716,1719
was|1720,1723
<EOL>|1724,1725
not|1725,1728
.|1728,1729
She|1730,1733
was|1734,1737
very|1738,1742
aware|1743,1748
of|1749,1751
her|1752,1755
dysarthria|1756,1766
and|1767,1770
told|1771,1775
her|1776,1779
daughters|1780,1789
<EOL>|1790,1791
that|1791,1795
she|1796,1799
thinks|1800,1806
she|1807,1810
's|1810,1812
having|1813,1819
a|1820,1821
stroke|1822,1828
.|1828,1829
Then|1830,1834
,|1834,1835
she|1836,1839
said|1840,1844
she|1845,1848
had|1849,1852
<EOL>|1853,1854
trouble|1854,1861
sitting|1862,1869
down|1870,1874
but|1875,1878
has|1879,1882
no|1883,1885
idea|1886,1890
why|1891,1894
she|1895,1898
thought|1899,1906
that|1907,1911
.|1911,1912
When|1913,1917
<EOL>|1918,1919
she|1919,1922
was|1923,1926
standing|1927,1935
,|1935,1936
she|1937,1940
was|1941,1944
able|1945,1949
to|1950,1952
walk|1953,1957
with|1958,1962
walker|1963,1969
but|1970,1973
she|1974,1977
felt|1978,1982
<EOL>|1983,1984
unsteady|1984,1992
and|1993,1996
almost|1997,2003
fell|2004,2008
.|2008,2009
No|2010,2012
visual|2013,2019
changes|2020,2027
.|2027,2028
No|2029,2031
numbness|2032,2040
or|2041,2043
<EOL>|2044,2045
tingling|2045,2053
.|2053,2054
Denies|2055,2061
focal|2062,2067
weakness|2068,2076
;|2076,2077
she|2078,2081
just|2082,2086
had|2087,2090
trouble|2091,2098
standing|2099,2107
<EOL>|2108,2109
up|2109,2111
.|2111,2112
She|2113,2116
was|2117,2120
able|2121,2125
to|2126,2128
unlock|2129,2135
her|2136,2139
door|2140,2144
without|2145,2152
issue|2153,2158
but|2159,2162
she|2163,2166
felt|2167,2171
<EOL>|2172,2173
shaky|2173,2178
.|2178,2179
<EOL>|2180,2181
<EOL>|2181,2182
She|2182,2185
was|2186,2189
brought|2190,2197
by|2198,2200
EMS|2201,2204
to|2205,2207
_|2208,2209
_|2209,2210
_|2210,2211
where|2212,2217
NIHSS|2218,2223
was|2224,2227
1|2228,2229
for|2230,2233
<EOL>|2234,2235
slurred|2235,2242
speech|2243,2249
.|2249,2250
There|2251,2256
,|2256,2257
she|2258,2261
felt|2262,2266
the|2267,2270
same|2271,2275
but|2276,2279
her|2280,2283
symptoms|2284,2292
<EOL>|2293,2294
started|2294,2301
to|2302,2304
improve|2305,2312
when|2313,2317
she|2318,2321
started|2322,2329
to|2330,2332
be|2333,2335
transferred|2336,2347
.|2347,2348
<EOL>|2349,2350
Paramedics|2350,2360
said|2361,2365
her|2366,2369
speech|2370,2376
was|2377,2380
improving|2381,2390
rapidly|2391,2398
en|2399,2401
route|2402,2407
.|2407,2408
<EOL>|2410,2411
<EOL>|2411,2412
Last|2412,2416
month|2417,2422
,|2422,2423
started|2424,2431
needing|2432,2439
naps|2440,2444
.|2444,2445
Her|2446,2449
hearing|2450,2457
is|2458,2460
poor|2461,2465
at|2466,2468
<EOL>|2469,2470
baseline|2470,2478
and|2479,2482
she|2483,2486
normally|2487,2495
uses|2496,2500
hearing|2501,2508
aids|2509,2513
.|2513,2514
<EOL>|2515,2516
<EOL>|2516,2517
For|2517,2520
the|2521,2524
past|2525,2529
_|2530,2531
_|2531,2532
_|2532,2533
months|2534,2540
,|2540,2541
she|2542,2545
has|2546,2549
had|2550,2553
_|2554,2555
_|2555,2556
_|2556,2557
nocturia|2558,2566
nightly|2567,2574
.|2574,2575
No|2576,2578
<EOL>|2579,2580
dysuria|2580,2587
.|2587,2588
<EOL>|2589,2590
<EOL>|2590,2591
She|2591,2594
has|2595,2598
noticed|2599,2606
more|2607,2611
frequent|2612,2620
headaches|2621,2630
lately|2631,2637
in|2638,2640
the|2641,2644
past|2645,2649
_|2650,2651
_|2651,2652
_|2652,2653
<EOL>|2654,2655
months|2655,2661
.|2661,2662
Last|2663,2667
headache|2668,2676
was|2677,2680
yesterday|2681,2690
.|2690,2691
She|2692,2695
takes|2696,2701
tramadol|2702,2710
and|2711,2714
<EOL>|2715,2716
acetaminophen|2716,2729
up|2730,2732
to|2733,2735
a|2736,2737
couple|2738,2744
times|2745,2750
a|2751,2752
night|2753,2758
.|2758,2759
She|2760,2763
reports|2764,2771
<EOL>|2772,2773
headaches|2773,2782
at|2783,2785
night|2786,2791
which|2792,2797
wake|2798,2802
her|2803,2806
up|2807,2809
.|2809,2810
She|2811,2814
denies|2815,2821
that|2822,2826
the|2827,2830
<EOL>|2831,2832
headache|2832,2840
is|2841,2843
<EOL>|2843,2844
positional|2844,2854
;|2854,2855
it|2856,2858
is|2859,2861
the|2862,2865
same|2866,2870
sitting|2871,2878
up|2879,2881
or|2882,2884
lying|2885,2890
down|2891,2895
.|2895,2896
She|2897,2900
has|2901,2904
had|2905,2908
<EOL>|2909,2910
some|2910,2914
gradual|2915,2922
weight|2923,2929
loss|2930,2934
over|2935,2939
the|2940,2943
past|2944,2948
~|2949,2950
12|2950,2952
months|2953,2959
;|2959,2960
_|2961,2962
_|2962,2963
_|2963,2964
year|2965,2969
ago|2970,2973
<EOL>|2974,2975
she|2975,2978
was|2979,2982
almost|2983,2989
140|2990,2993
lbs|2994,2997
,|2997,2998
and|2999,3002
now|3003,3006
she|3007,3010
is|3011,3013
_|3014,3015
_|3015,3016
_|3016,3017
lbs|3018,3021
.|3021,3022
Her|3023,3026
appetite|3027,3035
is|3036,3038
<EOL>|3039,3040
still|3040,3045
good|3046,3050
and|3051,3054
she|3055,3058
enjoys|3059,3065
eating|3066,3072
but|3073,3076
she|3077,3080
is|3081,3083
less|3084,3088
hungry|3089,3095
that|3096,3100
she|3101,3104
<EOL>|3105,3106
used|3106,3110
to|3111,3113
be|3114,3116
.|3116,3117
<EOL>|3119,3120
<EOL>|3120,3121
Daughter|3121,3129
says|3130,3134
that|3135,3139
she|3140,3143
has|3144,3147
had|3148,3151
marked|3152,3158
decline|3159,3166
in|3167,3169
memory|3170,3176
in|3177,3179
past|3180,3184
<EOL>|3185,3186
_|3186,3187
_|3187,3188
_|3188,3189
weeks|3190,3195
.|3195,3196
Over|3197,3201
past|3202,3206
few|3207,3210
years|3211,3216
,|3216,3217
she|3218,3221
has|3222,3225
been|3226,3230
forgetting|3231,3241
plans|3242,3247
,|3247,3248
<EOL>|3249,3250
times|3250,3255
for|3256,3259
pickpup|3260,3267
,|3267,3268
and|3269,3272
dinner|3273,3279
plans|3280,3285
,|3285,3286
which|3287,3292
has|3293,3296
become|3297,3303
normal|3304,3310
.|3310,3311
<EOL>|3312,3313
Over|3313,3317
the|3318,3321
past|3322,3326
_|3327,3328
_|3328,3329
_|3329,3330
weeks|3331,3336
,|3336,3337
family|3338,3344
has|3345,3348
noticed|3349,3356
dramatic|3357,3365
worsening|3366,3375
.|3375,3376
<EOL>|3377,3378
She|3378,3381
does|3382,3386
n't|3386,3389
remember|3390,3398
which|3399,3404
grandkids|3405,3414
were|3415,3419
coming|3420,3426
to|3427,3429
visit|3430,3435
when|3436,3440
<EOL>|3441,3442
she|3442,3445
bought|3446,3452
the|3453,3456
plane|3457,3462
tickets|3463,3470
herself|3471,3478
.|3478,3479
<EOL>|3479,3480
<EOL>|3480,3481
She|3481,3484
endorses|3485,3493
2|3494,3495
pillow|3496,3502
orthopnea|3503,3512
.|3512,3513
<EOL>|3514,3515
<EOL>|3516,3517
Divertoculosis|3539,3553
<EOL>|3553,3554
Atrial|3554,3560
fibrillation|3561,3573
on|3574,3576
Eliquis|3577,3584
<EOL>|3584,3585
CHF|3585,3588
<EOL>|3588,3589
Hypercholesterolemia|3589,3609
<EOL>|3609,3610
Hypertension|3610,3622
<EOL>|3622,3623
<EOL>|3624,3625
:|3639,3640
<EOL>|3640,3641
_|3641,3642
_|3642,3643
_|3643,3644
<EOL>|3644,3645
:|3659,3660
<EOL>|3660,3661
Father|3661,3667
-|3668,3669
severe|3670,3676
alcoholic|3677,3686
,|3686,3687
schizophrenia|3688,3701
<EOL>|3701,3702
Mother|3702,3708
-|3709,3710
CHF|3711,3714
<EOL>|3714,3715
Brother|3715,3722
-|3723,3724
stroke|3725,3731
,|3731,3732
carotid|3733,3740
stenosis|3741,3749
<EOL>|3749,3750
<EOL>|3751,3752
ADMISSION|3767,3776
EXAM|3777,3781
:|3781,3782
<EOL>|3782,3783
Vitals|3783,3789
:|3789,3790
T|3791,3792
:|3792,3793
97.9|3793,3797
HR|3800,3802
:|3802,3803
79|3804,3806
BP|3809,3811
:|3811,3812
164|3813,3816
/|3816,3817
121|3817,3820
RR|3823,3825
:|3825,3826
19|3827,3829
SaO2|3832,3836
:|3836,3837
94|3838,3840
%|3840,3841
on|3842,3844
RA|3845,3847
<EOL>|3847,3848
<EOL>|3848,3849
General|3849,3856
:|3856,3857
Awake|3858,3863
,|3863,3864
cooperative|3865,3876
elderly|3877,3884
woman|3885,3890
,|3890,3891
NAD|3892,3895
.|3895,3896
<EOL>|3896,3897
HEENT|3897,3902
:|3902,3903
NC|3904,3906
/|3906,3907
AT|3907,3909
,|3909,3910
no|3911,3913
scleral|3914,3921
icterus|3922,3929
noted|3930,3935
,|3935,3936
MMM|3937,3940
,|3940,3941
no|3942,3944
lesions|3945,3952
noted|3953,3958
in|3959,3961
<EOL>|3961,3962
oropharynx|3962,3972
.|3972,3973
<EOL>|3973,3974
Neck|3974,3978
:|3978,3979
Supple|3980,3986
.|3986,3987
No|3988,3990
nuchal|3991,3997
rigidity|3998,4006
.|4006,4007
<EOL>|4007,4008
Pulmonary|4008,4017
:|4017,4018
Normal|4019,4025
work|4026,4030
of|4031,4033
breathing|4034,4043
.|4043,4044
<EOL>|4044,4045
Cardiac|4045,4052
:|4052,4053
RRR|4054,4057
,|4057,4058
warm|4059,4063
,|4063,4064
well|4065,4069
-|4069,4070
perfused|4070,4078
.|4078,4079
<EOL>|4079,4080
Abdomen|4080,4087
:|4087,4088
Soft|4089,4093
,|4093,4094
non-distended|4095,4108
.|4108,4109
<EOL>|4109,4110
Extremities|4110,4121
:|4121,4122
No|4123,4125
_|4126,4127
_|4127,4128
_|4128,4129
edema|4130,4135
.|4135,4136
<EOL>|4136,4137
Skin|4137,4141
:|4141,4142
ecchymoses|4143,4153
in|4154,4156
L|4157,4158
shin|4159,4163
,|4163,4164
more|4165,4169
extensive|4170,4179
on|4180,4182
R|4183,4184
shin|4185,4189
.|4189,4190
<EOL>|4191,4192
<EOL>|4193,4194
Neurologic|4194,4204
:|4204,4205
<EOL>|4205,4206
-|4206,4207
Mental|4207,4213
Status|4214,4220
:|4220,4221
Alert|4222,4227
,|4227,4228
oriented|4229,4237
_|4238,4239
_|4239,4240
_|4240,4241
.|4241,4242
<EOL>|4242,4243
Able|4243,4247
to|4248,4250
relate|4251,4257
history|4258,4265
without|4266,4273
difficulty.|4274,4285
Attentive|4286,4295
,|4295,4296
able|4297,4301
to|4302,4304
<EOL>|4304,4305
name|4305,4309
_|4310,4311
_|4311,4312
_|4312,4313
backward|4314,4322
without|4323,4330
difficulty.|4331,4342
Language|4343,4351
is|4352,4354
fluent|4355,4361
with|4362,4366
<EOL>|4366,4367
intact|4367,4373
repetition|4374,4384
and|4385,4388
comprehension|4389,4402
.|4402,4403
Normal|4404,4410
prosody|4411,4418
.|4418,4419
There|4420,4425
were|4426,4430
<EOL>|4430,4431
no|4431,4433
paraphasic|4434,4444
errors|4445,4451
.|4451,4452
Able|4453,4457
to|4458,4460
name|4461,4465
both|4466,4470
high|4471,4475
and|4476,4479
low|4480,4483
frequency|4484,4493
<EOL>|4493,4494
objects|4494,4501
.|4501,4502
Able|4504,4508
to|4509,4511
read|4512,4516
without|4517,4524
difficulty|4525,4535
.|4535,4536
No|4537,4539
dysarthria|4540,4550
.|4550,4551
Able|4552,4556
<EOL>|4557,4558
to|4558,4560
<EOL>|4560,4561
follow|4561,4567
both|4568,4572
midline|4573,4580
and|4581,4584
appendicular|4585,4597
commands|4598,4606
.|4606,4607
There|4608,4613
was|4614,4617
no|4618,4620
<EOL>|4620,4621
evidence|4621,4629
of|4630,4632
apraxia|4633,4640
or|4641,4643
neglect|4644,4651
.|4651,4652
<EOL>|4652,4653
<EOL>|4653,4654
-|4654,4655
Cranial|4655,4662
Nerves|4663,4669
:|4669,4670
<EOL>|4670,4671
II|4671,4673
,|4673,4674
III|4675,4678
,|4678,4679
IV|4680,4682
,|4682,4683
VI|4684,4686
:|4686,4687
PERRL|4689,4694
3|4695,4696
to|4697,4699
2mm|4700,4703
and|4704,4707
brisk|4708,4713
.|4713,4714
EOMI|4715,4719
without|4720,4727
<EOL>|4727,4728
nystagmus|4728,4737
.|4737,4738
Normal|4739,4745
saccades|4746,4754
.|4754,4755
VFF|4756,4759
to|4760,4762
confrontation|4763,4776
.|4776,4777
<EOL>|4778,4779
V|4779,4780
:|4780,4781
Facial|4782,4788
sensation|4789,4798
intact|4799,4805
to|4806,4808
light|4809,4814
touch|4815,4820
and|4821,4824
pinprick|4825,4833
.|4833,4834
<EOL>|4834,4835
VII|4835,4838
:|4838,4839
No|4840,4842
facial|4843,4849
droop|4850,4855
,|4855,4856
facial|4857,4863
musculature|4864,4875
symmetric|4876,4885
.|4885,4886
<EOL>|4886,4887
VIII|4887,4891
:|4891,4892
Hearing|4893,4900
intact|4901,4907
to|4908,4910
finger|4911,4917
snapping|4918,4926
b|4927,4928
/|4928,4929
l|4929,4930
.|4930,4931
Did|4932,4935
not|4936,4939
bring|4940,4945
her|4946,4949
<EOL>|4949,4950
hearing|4950,4957
aids|4958,4962
.|4962,4963
<EOL>|4964,4965
IX|4965,4967
,|4967,4968
X|4969,4970
:|4970,4971
Palate|4972,4978
elevates|4979,4987
symmetrically|4988,5001
.|5001,5002
<EOL>|5002,5003
XI|5003,5005
:|5005,5006
_|5007,5008
_|5008,5009
_|5009,5010
strength|5011,5019
in|5020,5022
trapezii|5023,5031
bilaterally|5032,5043
.|5043,5044
<EOL>|5044,5045
XII|5045,5048
:|5048,5049
Tongue|5050,5056
protrudes|5057,5066
in|5067,5069
midline|5070,5077
with|5078,5082
good|5083,5087
excursions|5088,5098
.|5098,5099
Strength|5100,5108
<EOL>|5108,5109
full|5109,5113
with|5114,5118
tongue|5119,5125
-|5125,5126
in|5126,5128
-|5128,5129
cheek|5129,5134
testing|5135,5142
.|5142,5143
<EOL>|5143,5144
<EOL>|5144,5145
-|5145,5146
Motor|5146,5151
:|5151,5152
Normal|5153,5159
bulk|5160,5164
and|5165,5168
tone|5169,5173
throughout|5174,5184
.|5184,5185
No|5186,5188
pronator|5189,5197
drift|5198,5203
.|5203,5204
No|5205,5207
<EOL>|5207,5208
adventitious|5208,5220
movements|5221,5230
,|5230,5231
such|5232,5236
as|5237,5239
tremor|5240,5246
or|5247,5249
asterixis|5250,5259
noted|5260,5265
.|5265,5266
<EOL>|5266,5267
[|5269,5270
_|5270,5271
_|5271,5272
_|5272,5273
]|5273,5274
<EOL>|5274,5275
L|5275,5276
5|5280,5281
5|5285,5286
5|5290,5291
5|5295,5296
5|5300,5301
5|5305,5306
5|5309,5310
5|5314,5315
5|5319,5320
5|5323,5324
5|5328,5329
5|5333,5334
<EOL>|5334,5335
R|5335,5336
5|5340,5341
5|5345,5346
5|5350,5351
5|5355,5356
5|5360,5361
5|5365,5366
5|5369,5370
5|5374,5375
5|5379,5380
5|5383,5384
5|5388,5389
5|5393,5394
<EOL>|5394,5395
<EOL>|5395,5396
-|5396,5397
Sensory|5397,5404
:|5404,5405
No|5406,5408
deficits|5409,5417
to|5418,5420
light|5421,5426
touch|5427,5432
,|5432,5433
pinprick|5434,5442
,|5442,5443
temperature|5444,5455
<EOL>|5455,5456
throughout|5456,5466
.|5466,5467
Decreased|5468,5477
vibratory|5478,5487
sense|5488,5493
in|5494,5496
b|5497,5498
/|5498,5499
l|5499,5500
feet|5501,5505
up|5506,5508
to|5509,5511
ankles|5512,5518
.|5518,5519
<EOL>|5519,5520
Joint|5520,5525
position|5526,5534
sense|5535,5540
intact|5541,5547
in|5548,5550
b|5551,5552
/|5552,5553
l|5553,5554
great|5555,5560
toes|5561,5565
.|5565,5566
No|5567,5569
extinction|5570,5580
to|5581,5583
<EOL>|5583,5584
DSS|5584,5587
.|5587,5588
Romberg|5589,5596
absent|5597,5603
.|5603,5604
<EOL>|5604,5605
<EOL>|5605,5606
-|5606,5607
Reflexes|5607,5615
:|5615,5616
<EOL>|5616,5617
[|5619,5620
Bic|5620,5623
]|5623,5624
[|5625,5626
Tri|5626,5629
]|5629,5630
[|5631,5632
_|5632,5633
_|5633,5634
_|5634,5635
]|5635,5636
[|5637,5638
Pat|5638,5641
]|5641,5642
[|5643,5644
Ach|5644,5647
]|5647,5648
<EOL>|5648,5649
L|5649,5650
2|5653,5654
+|5654,5655
2|5659,5660
2|5666,5667
2|5673,5674
+|5674,5675
0|5679,5680
<EOL>|5680,5681
R|5681,5682
2|5685,5686
+|5686,5687
2|5691,5692
2|5698,5699
2|5705,5706
+|5706,5707
0|5711,5712
<EOL>|5713,5714
Plantar|5714,5721
response|5722,5730
was|5731,5734
flexor|5735,5741
bilaterally|5742,5753
.|5753,5754
<EOL>|5754,5755
<EOL>|5755,5756
-|5756,5757
Coordination|5757,5769
:|5769,5770
No|5771,5773
intention|5774,5783
tremor|5784,5790
.|5790,5791
No|5793,5795
dysmetria|5796,5805
on|5806,5808
FNF|5809,5812
<EOL>|5812,5813
bilaterally|5813,5824
.|5824,5825
HKS|5826,5829
with|5830,5834
L|5835,5836
heel|5837,5841
without|5842,5849
dysmetria|5850,5859
.|5859,5860
Unable|5861,5867
to|5868,5870
bend|5871,5875
R|5876,5877
<EOL>|5877,5878
knee|5878,5882
due|5883,5886
to|5887,5889
knee|5890,5894
surgery|5895,5902
.|5902,5903
<EOL>|5904,5905
<EOL>|5905,5906
-|5906,5907
Gait|5907,5911
:|5911,5912
unable|5913,5919
to|5920,5922
assess|5923,5929
as|5930,5932
patient|5933,5940
needs|5941,5946
a|5947,5948
walker|5949,5955
at|5956,5958
baseline|5959,5967
<EOL>|5967,5968
<EOL>|5968,5969
DISCHARGE|5969,5978
EXAM|5979,5983
:|5983,5984
<EOL>|5984,5985
24|5985,5987
HR|5988,5990
Data|5991,5995
(|5996,5997
last|5997,6001
updated|6002,6009
_|6010,6011
_|6011,6012
_|6012,6013
@|6014,6015
419|6016,6019
)|6019,6020
<EOL>|6020,6021
Temp|6021,6025
:|6025,6026
97.4|6027,6031
(|6032,6033
Tm|6033,6035
98.6|6036,6040
)|6040,6041
,|6041,6042
BP|6043,6045
:|6045,6046
146|6047,6050
/|6050,6051
76|6051,6053
(|6054,6055
116|6055,6058
-|6058,6059
155|6059,6062
/|6062,6063
65|6063,6065
-|6065,6066
94|6066,6068
)|6068,6069
,|6069,6070
HR|6071,6073
:|6073,6074
53|6075,6077
<EOL>|6078,6079
(|6079,6080
53|6080,6082
-|6082,6083
86|6083,6085
)|6085,6086
,|6086,6087
<EOL>|6087,6088
RR|6088,6090
:|6090,6091
17|6092,6094
(|6095,6096
_|6096,6097
_|6097,6098
_|6098,6099
)|6099,6100
,|6100,6101
O2|6102,6104
sat|6105,6108
:|6108,6109
96|6110,6112
%|6112,6113
(|6114,6115
92|6115,6117
-|6117,6118
97|6118,6120
)|6120,6121
,|6121,6122
O2|6123,6125
delivery|6126,6134
:|6134,6135
Ra|6136,6138
<EOL>|6138,6139
<EOL>|6139,6140
General|6140,6147
:|6147,6148
Awake|6149,6154
,|6154,6155
cooperative|6156,6167
elderly|6168,6175
woman|6176,6181
,|6181,6182
NAD|6183,6186
.|6186,6187
<EOL>|6187,6188
HEENT|6188,6193
:|6193,6194
NC|6195,6197
/|6197,6198
AT|6198,6200
,|6200,6201
no|6202,6204
scleral|6205,6212
icterus|6213,6220
noted|6221,6226
,|6226,6227
MMM|6228,6231
,|6231,6232
no|6233,6235
lesions|6236,6243
noted|6244,6249
in|6250,6252
<EOL>|6252,6253
oropharynx|6253,6263
.|6263,6264
<EOL>|6264,6265
Neck|6265,6269
:|6269,6270
Supple|6271,6277
.|6277,6278
No|6279,6281
nuchal|6282,6288
rigidity|6289,6297
.|6297,6298
<EOL>|6298,6299
Pulmonary|6299,6308
:|6308,6309
Normal|6310,6316
work|6317,6321
of|6322,6324
breathing|6325,6334
.|6334,6335
<EOL>|6335,6336
Cardiac|6336,6343
:|6343,6344
NR|6345,6347
,|6347,6348
RR|6349,6351
,|6351,6352
warm|6353,6357
,|6357,6358
well|6359,6363
-|6363,6364
perfused|6364,6372
.|6372,6373
<EOL>|6373,6374
Abdomen|6374,6381
:|6381,6382
Soft|6383,6387
,|6387,6388
non-distended|6389,6402
.|6402,6403
<EOL>|6403,6404
Extremities|6404,6415
:|6415,6416
No|6417,6419
_|6420,6421
_|6421,6422
_|6422,6423
edema|6424,6429
.|6429,6430
<EOL>|6430,6431
Skin|6431,6435
:|6435,6436
ecchymoses|6437,6447
in|6448,6450
L|6451,6452
shin|6453,6457
,|6457,6458
more|6459,6463
extensive|6464,6473
on|6474,6476
R|6477,6478
shin|6479,6483
.|6483,6484
<EOL>|6485,6486
<EOL>|6487,6488
Neurologic|6488,6498
:|6498,6499
<EOL>|6499,6500
-|6500,6501
Mental|6501,6507
Status|6508,6514
:|6514,6515
Alert|6516,6521
,|6521,6522
oriented|6523,6531
to|6532,6534
person|6535,6541
and|6542,6545
situation|6546,6555
.|6555,6556
Able|6557,6561
to|6562,6564
<EOL>|6564,6565
relate|6565,6571
history|6572,6579
without|6580,6587
difficulty.|6588,6599
Attentive|6600,6609
to|6610,6612
examiner|6613,6621
.|6621,6622
<EOL>|6622,6623
Language|6623,6631
is|6632,6634
fluent|6635,6641
with|6642,6646
intact|6647,6653
comprehension|6654,6667
.|6667,6668
Normal|6669,6675
prosody|6676,6683
.|6683,6684
<EOL>|6684,6685
There|6685,6690
were|6691,6695
no|6696,6698
paraphasic|6699,6709
errors|6710,6716
.|6716,6717
No|6718,6720
dysarthria|6721,6731
.|6731,6732
Able|6733,6737
to|6738,6740
follow|6741,6747
<EOL>|6747,6748
both|6748,6752
midline|6753,6760
and|6761,6764
appendicular|6765,6777
commands|6778,6786
.|6786,6787
There|6788,6793
was|6794,6797
no|6798,6800
evidence|6801,6809
of|6810,6812
<EOL>|6812,6813
apraxia|6813,6820
or|6821,6823
neglect|6824,6831
.|6831,6832
<EOL>|6832,6833
<EOL>|6833,6834
-|6834,6835
Cranial|6835,6842
Nerves|6843,6849
:|6849,6850
<EOL>|6850,6851
II|6851,6853
,|6853,6854
III|6855,6858
,|6858,6859
IV|6860,6862
,|6862,6863
VI|6864,6866
:|6866,6867
PERRL|6869,6874
3|6875,6876
to|6877,6879
2mm|6880,6883
and|6884,6887
brisk|6888,6893
.|6893,6894
EOMI|6895,6899
without|6900,6907
<EOL>|6907,6908
nystagmus|6908,6917
.|6917,6918
Normal|6919,6925
saccades|6926,6934
.|6934,6935
<EOL>|6935,6936
V|6936,6937
:|6937,6938
Facial|6939,6945
sensation|6946,6955
intact|6956,6962
to|6963,6965
light|6966,6971
touch|6972,6977
.|6977,6978
<EOL>|6978,6979
VII|6979,6982
:|6982,6983
No|6984,6986
facial|6987,6993
droop|6994,6999
,|6999,7000
facial|7001,7007
musculature|7008,7019
symmetric|7020,7029
.|7029,7030
<EOL>|7030,7031
VIII|7031,7035
:|7035,7036
Hearing|7037,7044
intact|7045,7051
to|7052,7054
conversation|7055,7067
.|7067,7068
<EOL>|7068,7069
IX|7069,7071
,|7071,7072
X|7073,7074
:|7074,7075
Palate|7076,7082
elevates|7083,7091
symmetrically|7092,7105
.|7105,7106
<EOL>|7106,7107
XI|7107,7109
:|7109,7110
_|7111,7112
_|7112,7113
_|7113,7114
strength|7115,7123
in|7124,7126
trapezii|7127,7135
bilaterally|7136,7147
.|7147,7148
<EOL>|7148,7149
XII|7149,7152
:|7152,7153
Tongue|7154,7160
protrudes|7161,7170
in|7171,7173
midline|7174,7181
with|7182,7186
good|7187,7191
excursions|7192,7202
.|7202,7203
<EOL>|7203,7204
<EOL>|7204,7205
-|7205,7206
Motor|7206,7211
:|7211,7212
Normal|7213,7219
bulk|7220,7224
and|7225,7228
tone|7229,7233
throughout|7234,7244
.|7244,7245
No|7246,7248
pronator|7249,7257
drift|7258,7263
.|7263,7264
No|7265,7267
<EOL>|7267,7268
adventitious|7268,7280
movements|7281,7290
,|7290,7291
such|7292,7296
as|7297,7299
tremor|7300,7306
or|7307,7309
asterixis|7310,7319
noted|7320,7325
.|7325,7326
<EOL>|7326,7327
[|7329,7330
Delt|7330,7334
]|7334,7335
[|7335,7336
Bic|7336,7339
]|7339,7340
[|7340,7341
Tri|7341,7344
]|7344,7345
[|7345,7346
ECR|7346,7349
]|7349,7350
[|7350,7351
FEx|7351,7354
]|7354,7355
[|7355,7356
IO|7356,7358
]|7358,7359
[|7359,7360
IP|7360,7362
]|7362,7363
[|7363,7364
Quad|7364,7368
]|7368,7369
[|7369,7370
Ham|7370,7373
]|7373,7374
[|7374,7375
TA|7375,7377
]|7377,7378
[|7378,7379
Gas|7379,7382
]|7382,7383
<EOL>|7383,7384
L|7384,7385
5|7389,7390
5|7394,7395
5|7399,7400
5|7404,7405
5|7409,7410
5|7414,7415
5|7418,7419
5|7423,7424
5|7428,7429
5|7432,7433
5|7437,7438
<EOL>|7442,7443
R|7443,7444
5|7448,7449
5|7453,7454
5|7458,7459
5|7463,7464
5|7468,7469
5|7473,7474
5|7477,7478
*|7482,7483
*|7487,7488
5|7491,7492
5|7496,7497
<EOL>|7501,7502
*|7502,7503
Knee|7503,7507
can|7508,7511
not|7511,7514
bend|7515,7519
after|7520,7525
prior|7526,7531
surgery|7532,7539
<EOL>|7539,7540
<EOL>|7540,7541
-|7541,7542
Sensory|7542,7549
:|7549,7550
No|7551,7553
deficits|7554,7562
to|7563,7565
light|7566,7571
touch|7572,7577
throughout|7578,7588
.|7588,7589
<EOL>|7589,7590
<EOL>|7590,7591
-|7591,7592
Coordination|7592,7604
:|7604,7605
No|7606,7608
intention|7609,7618
tremor|7619,7625
.|7625,7626
No|7628,7630
dysmetria|7631,7640
on|7641,7643
FNF|7644,7647
<EOL>|7647,7648
bilaterally|7648,7659
.|7659,7660
<EOL>|7661,7662
<EOL>|7662,7663
-|7663,7664
Gait|7664,7668
:|7668,7669
needs|7670,7675
a|7676,7677
walker|7678,7684
at|7685,7687
baseline|7688,7696
<EOL>|7696,7697
<EOL>|7698,7699
Pertinent|7699,7708
Results|7709,7716
:|7716,7717
<EOL>|7717,7718
_|7718,7719
_|7719,7720
_|7720,7721
01|7722,7724
:|7724,7725
50AM|7725,7729
BLOOD|7730,7735
WBC|7736,7739
-|7739,7740
7.2|7740,7743
RBC|7744,7747
-|7747,7748
4|7748,7749
.|7749,7750
75|7750,7752
Hgb|7753,7756
-|7756,7757
14.6|7757,7761
Hct|7762,7765
-|7765,7766
45|7766,7768
.|7768,7769
5|7769,7770
*|7770,7771
<EOL>|7772,7773
MCV|7773,7776
-|7776,7777
96|7777,7779
MCH|7780,7783
-|7783,7784
30.7|7784,7788
MCHC|7789,7793
-|7793,7794
32.1|7794,7798
RDW|7799,7802
-|7802,7803
13.2|7803,7807
RDWSD|7808,7813
-|7813,7814
46|7814,7816
.|7816,7817
5|7817,7818
*|7818,7819
Plt|7820,7823
_|7824,7825
_|7825,7826
_|7826,7827
<EOL>|7827,7828
_|7828,7829
_|7829,7830
_|7830,7831
01|7832,7834
:|7834,7835
50AM|7835,7839
BLOOD|7840,7845
Neuts|7846,7851
-|7851,7852
53.1|7852,7856
_|7857,7858
_|7858,7859
_|7859,7860
Monos|7861,7866
-|7866,7867
8.2|7867,7870
Eos|7871,7874
-|7874,7875
1.5|7875,7878
<EOL>|7879,7880
Baso|7880,7884
-|7884,7885
0.3|7885,7888
Im|7889,7891
_|7892,7893
_|7893,7894
_|7894,7895
AbsNeut|7896,7903
-|7903,7904
3|7904,7905
.|7905,7906
81|7906,7908
AbsLymp|7909,7916
-|7916,7917
2|7917,7918
.|7918,7919
63|7919,7921
AbsMono|7922,7929
-|7929,7930
0|7930,7931
.|7931,7932
59|7932,7934
<EOL>|7935,7936
AbsEos|7936,7942
-|7942,7943
0|7943,7944
.|7944,7945
11|7945,7947
AbsBaso|7948,7955
-|7955,7956
0|7956,7957
.|7957,7958
02|7958,7960
<EOL>|7960,7961
_|7961,7962
_|7962,7963
_|7963,7964
01|7965,7967
:|7967,7968
50AM|7968,7972
BLOOD|7973,7978
_|7979,7980
_|7980,7981
_|7981,7982
PTT|7983,7986
-|7986,7987
29.7|7987,7991
_|7992,7993
_|7993,7994
_|7994,7995
<EOL>|7995,7996
_|7996,7997
_|7997,7998
_|7998,7999
01|8000,8002
:|8002,8003
50AM|8003,8007
BLOOD|8008,8013
Glucose|8014,8021
-|8021,8022
97|8022,8024
UreaN|8025,8030
-|8030,8031
18|8031,8033
Creat|8034,8039
-|8039,8040
0.7|8040,8043
Na|8044,8046
-|8046,8047
139|8047,8050
<EOL>|8051,8052
K|8052,8053
-|8053,8054
4.3|8054,8057
Cl|8058,8060
-|8060,8061
102|8061,8064
HCO3|8065,8069
-|8069,8070
26|8070,8072
AnGap|8073,8078
-|8078,8079
11|8079,8081
<EOL>|8081,8082
_|8082,8083
_|8083,8084
_|8084,8085
07|8086,8088
:|8088,8089
35AM|8089,8093
BLOOD|8094,8099
CK|8100,8102
-|8102,8103
MB|8103,8105
-|8105,8106
4|8106,8107
cTropnT|8108,8115
-|8115,8116
<|8116,8117
0|8117,8118
.|8118,8119
01|8119,8121
<EOL>|8121,8122
_|8122,8123
_|8123,8124
_|8124,8125
07|8126,8128
:|8128,8129
35AM|8129,8133
BLOOD|8134,8139
Calcium|8140,8147
-|8147,8148
9.3|8148,8151
Phos|8152,8156
-|8156,8157
3.6|8157,8160
Mg|8161,8163
-|8163,8164
1.8|8164,8167
Cholest|8168,8175
-|8175,8176
207|8176,8179
*|8179,8180
<EOL>|8180,8181
_|8181,8182
_|8182,8183
_|8183,8184
07|8185,8187
:|8187,8188
35AM|8188,8192
BLOOD|8193,8198
Triglyc|8199,8206
-|8206,8207
62|8207,8209
HDL|8210,8213
-|8213,8214
69|8214,8216
CHOL|8217,8221
/|8221,8222
HD|8222,8224
-|8224,8225
3.0|8225,8228
LDLcalc|8229,8236
-|8236,8237
126|8237,8240
<EOL>|8240,8241
_|8241,8242
_|8242,8243
_|8243,8244
10|8245,8247
:|8247,8248
57AM|8248,8252
BLOOD|8253,8258
%|8259,8260
HbA1c|8260,8265
-|8265,8266
5.5|8266,8269
eAG|8270,8273
-|8273,8274
111|8274,8277
<EOL>|8277,8278
_|8278,8279
_|8279,8280
_|8280,8281
05|8282,8284
:|8284,8285
22AM|8285,8289
BLOOD|8290,8295
VitB12|8296,8302
-|8302,8303
249|8303,8306
<EOL>|8306,8307
_|8307,8308
_|8308,8309
_|8309,8310
05|8311,8313
:|8313,8314
22AM|8314,8318
BLOOD|8319,8324
TSH|8325,8328
-|8328,8329
5|8329,8330
.|8330,8331
8|8331,8332
*|8332,8333
<EOL>|8333,8334
_|8334,8335
_|8335,8336
_|8336,8337
05|8338,8340
:|8340,8341
22AM|8341,8345
BLOOD|8346,8351
Trep|8352,8356
Ab|8357,8359
-|8359,8360
NEG|8360,8363
<EOL>|8363,8364
_|8364,8365
_|8365,8366
_|8366,8367
03|8368,8370
:|8370,8371
12AM|8371,8375
URINE|8376,8381
Color|8382,8387
-|8387,8388
Straw|8388,8393
Appear|8394,8400
-|8400,8401
Clear|8401,8406
Sp|8407,8409
_|8410,8411
_|8411,8412
_|8412,8413
<EOL>|8413,8414
_|8414,8415
_|8415,8416
_|8416,8417
03|8418,8420
:|8420,8421
12AM|8421,8425
URINE|8426,8431
Blood|8432,8437
-|8437,8438
NEG|8438,8441
Nitrite|8442,8449
-|8449,8450
NEG|8450,8453
Protein|8454,8461
-|8461,8462
NEG|8462,8465
<EOL>|8466,8467
Glucose|8467,8474
-|8474,8475
NEG|8475,8478
Ketone|8479,8485
-|8485,8486
NEG|8486,8489
Bilirub|8490,8497
-|8497,8498
NEG|8498,8501
Urobiln|8502,8509
-|8509,8510
NEG|8510,8513
pH|8514,8516
-|8516,8517
6.5|8517,8520
Leuks|8521,8526
-|8526,8527
NEG|8527,8530
<EOL>|8530,8531
<EOL>|8531,8532
_|8532,8533
_|8533,8534
_|8534,8535
OSH|8536,8539
CTA|8540,8543
head|8544,8548
/|8548,8549
neck|8549,8553
_|8554,8555
_|8555,8556
_|8556,8557
opinion|8558,8565
(|8566,8567
_|8567,8568
_|8568,8569
_|8569,8570
)|8570,8571
<EOL>|8571,8572
1.|8585,8587
Segmental|8589,8598
left|8599,8603
vertebral|8604,8613
artery|8614,8620
occlusion|8621,8630
of|8631,8633
indeterminate|8634,8647
<EOL>|8648,8649
chronicity|8649,8659
.|8659,8660
No|8662,8664
evidence|8665,8673
of|8674,8676
ischemia|8677,8685
.|8685,8686
<EOL>|8686,8687
2.|8687,8689
Somewhat|8691,8699
small|8700,8705
caliber|8706,8713
attenuated|8714,8724
left|8725,8729
M2|8730,8732
inferior|8733,8741
branch|8742,8748
,|8748,8749
<EOL>|8750,8751
without|8751,8758
evidence|8759,8767
of|8768,8770
focal|8771,8776
occlusion|8777,8786
.|8786,8787
<EOL>|8787,8788
3.|8788,8790
No|8792,8794
acute|8795,8800
intracranial|8801,8813
abnormality|8814,8825
on|8826,8828
noncontrast|8829,8840
CT|8841,8843
head|8844,8848
.|8848,8849
<EOL>|8849,8850
<EOL>|8850,8851
_|8851,8852
_|8852,8853
_|8853,8854
MRI|8855,8858
head|8859,8863
w|8864,8865
/|8865,8866
o|8866,8867
contrast|8868,8876
<EOL>|8876,8877
1|8889,8890
.|8890,8891
No|8892,8894
acute|8895,8900
intracranial|8901,8913
abnormality|8914,8925
.|8925,8926
Specifically|8928,8940
,|8940,8941
no|8942,8944
large|8945,8950
<EOL>|8951,8952
territory|8952,8961
infarction|8962,8972
or|8973,8975
hemorrhage|8976,8986
.|8986,8987
<EOL>|8987,8988
2.|8988,8990
Scattered|8991,9000
foci|9001,9005
of|9006,9008
T2|9009,9011
/|9011,9012
high|9012,9016
-|9016,9017
signal|9017,9023
intensity|9024,9033
in|9034,9036
the|9037,9040
subcortical|9041,9052
<EOL>|9053,9054
and|9054,9057
periventricular|9058,9073
white|9074,9079
matter|9080,9086
are|9087,9090
nonspecific|9091,9102
and|9103,9106
may|9107,9110
reflect|9111,9118
<EOL>|9119,9120
changes|9120,9127
due|9128,9131
to|9132,9134
chronic|9135,9142
small|9143,9148
vessel|9149,9155
disease|9156,9163
.|9163,9164
<EOL>|9164,9165
<EOL>|9165,9166
_|9166,9167
_|9167,9168
_|9168,9169
TTE|9170,9173
<EOL>|9173,9174
IMPRESSION|9174,9184
:|9184,9185
No|9186,9188
structural|9189,9199
source|9200,9206
of|9207,9209
thromboembolism|9210,9225
identified|9226,9236
<EOL>|9237,9238
(|9238,9239
underlying|9239,9249
rhythm|9250,9256
predisposes|9257,9268
to|9269,9271
thrombus|9272,9280
formation|9281,9290
)|9290,9291
.|9291,9292
Preserved|9293,9302
<EOL>|9303,9304
left|9304,9308
ventricular|9309,9320
systolic|9321,9329
function|9330,9338
in|9339,9341
the|9342,9345
setting|9346,9353
of|9354,9356
<EOL>|9357,9358
beat|9358,9362
-|9362,9363
to|9363,9365
-|9365,9366
beat|9366,9370
variability|9371,9382
due|9383,9386
to|9387,9389
arrhythmia|9390,9400
.|9400,9401
Mild|9402,9406
to|9407,9409
moderate|9410,9418
<EOL>|9419,9420
mitral|9420,9426
and|9427,9430
tricuspid|9431,9440
regurgitation|9441,9454
.|9454,9455
Normal|9456,9462
pulmonary|9463,9472
pressure|9473,9481
.|9481,9482
<EOL>|9483,9484
Very|9484,9488
small|9489,9494
pericardial|9495,9506
effusion|9507,9515
<EOL>|9515,9516
<EOL>|9517,9518
Ms.|9541,9544
_|9545,9546
_|9546,9547
_|9547,9548
is|9549,9551
a|9552,9553
_|9554,9555
_|9555,9556
_|9556,9557
year|9558,9562
old|9563,9566
female|9567,9573
with|9574,9578
AFib|9579,9583
on|9584,9586
Eliquis|9587,9594
,|9594,9595
CHF|9596,9599
,|9599,9600
<EOL>|9601,9602
HLD|9602,9605
,|9605,9606
HTN|9607,9610
who|9611,9614
presented|9615,9624
w|9625,9626
/|9626,9627
sudden|9628,9634
onset|9635,9640
dysarthria|9641,9651
,|9651,9652
abnormal|9653,9661
arm|9662,9665
<EOL>|9666,9667
movements|9667,9676
,|9676,9677
and|9678,9681
poor|9682,9686
balance|9687,9694
(|9695,9696
walker|9696,9702
at|9703,9705
baseline|9706,9714
)|9714,9715
.|9715,9716
NIHSS|9717,9722
1|9723,9724
for|9725,9728
<EOL>|9729,9730
slurred|9730,9737
speech|9738,9744
at|9745,9747
OSH|9748,9751
.|9751,9752
There|9753,9758
,|9758,9759
a|9760,9761
CTA|9762,9765
head|9766,9770
and|9771,9774
neck|9775,9779
was|9780,9783
completed|9784,9793
,|9793,9794
<EOL>|9795,9796
and|9796,9799
there|9800,9805
was|9806,9809
concern|9810,9817
for|9818,9821
left|9822,9826
M2|9827,9829
branch|9830,9836
attenuation|9837,9848
concerning|9849,9859
<EOL>|9860,9861
for|9861,9864
stenosis|9865,9873
or|9874,9876
occlusion|9877,9886
,|9886,9887
and|9888,9891
she|9892,9895
was|9896,9899
subsequently|9900,9912
transferred|9913,9924
<EOL>|9925,9926
for|9926,9929
consideration|9930,9943
of|9944,9946
thrombectomy|9947,9959
but|9960,9963
NIHSS|9964,9969
0|9970,9971
on|9972,9974
arrival|9975,9982
so|9983,9985
she|9986,9989
<EOL>|9990,9991
was|9991,9994
not|9995,9998
deemed|9999,10005
a|10006,10007
candidate|10008,10017
.|10017,10018
She|10019,10022
was|10023,10026
admitted|10027,10035
to|10036,10038
the|10039,10042
Neurology|10043,10052
<EOL>|10053,10054
stroke|10054,10060
service|10061,10068
for|10069,10072
further|10073,10080
evaluation|10081,10091
of|10092,10094
possible|10095,10103
TIA|10104,10107
vs|10108,10110
stroke|10111,10117
.|10117,10118
<EOL>|10119,10120
No|10120,10122
further|10123,10130
symptoms|10131,10139
noted|10140,10145
during|10146,10152
admission|10153,10162
.|10162,10163
MRI|10164,10167
head|10168,10172
w|10173,10174
/|10174,10175
o|10175,10176
<EOL>|10177,10178
contrast|10178,10186
were|10187,10191
without|10192,10199
evidence|10200,10208
of|10209,10211
stroke|10212,10218
.|10218,10219
Reports|10220,10227
recent|10228,10234
<EOL>|10235,10236
echocardiogram|10236,10250
per|10251,10254
outpatient|10255,10265
PCP|10266,10269
/|10269,10270
cardiologist|10270,10282
,|10282,10283
reported|10284,10292
as|10293,10295
no|10296,10298
<EOL>|10299,10300
acute|10300,10305
findings|10306,10314
and|10315,10318
so|10319,10321
this|10322,10326
was|10327,10330
not|10331,10334
repeated|10335,10343
.|10343,10344
She|10345,10348
mentioned|10349,10358
<EOL>|10359,10360
concern|10360,10367
about|10368,10373
worsening|10374,10383
memory|10384,10390
,|10390,10391
but|10392,10395
able|10396,10400
to|10401,10403
perform|10404,10411
ADLs|10412,10416
w|10417,10418
/|10418,10419
<EOL>|10420,10421
meals|10421,10426
/|10426,10427
cleaning|10427,10435
provided|10436,10444
by|10445,10447
ALF|10448,10451
(|10452,10453
moved|10453,10458
10|10459,10461
months|10462,10468
ago|10469,10472
)|10472,10473
;|10473,10474
it|10475,10477
appears|10478,10485
<EOL>|10486,10487
there|10487,10492
has|10493,10496
been|10497,10501
no|10502,10504
acute|10505,10510
change|10511,10517
.|10517,10518
She|10519,10522
was|10523,10526
taking|10527,10533
apixiban|10534,10542
2.5|10543,10546
mg|10546,10548
<EOL>|10549,10550
once|10550,10554
daily|10555,10560
(|10561,10562
unclear|10562,10569
why|10570,10573
as|10574,10576
this|10577,10581
is|10582,10584
a|10585,10586
BID|10587,10590
medication|10591,10601
)|10601,10602
,|10602,10603
and|10604,10607
so|10608,10610
her|10611,10614
<EOL>|10615,10616
dose|10616,10620
was|10621,10624
increased|10625,10634
to|10635,10637
2.5|10638,10641
mg|10641,10643
BID|10644,10647
(|10648,10649
she|10649,10652
was|10653,10656
not|10657,10660
a|10661,10662
candidate|10663,10672
for|10673,10676
5mg|10677,10680
<EOL>|10681,10682
BID|10682,10685
due|10686,10689
to|10690,10692
her|10693,10696
age|10697,10700
and|10701,10704
weight|10705,10711
)|10711,10712
.|10712,10713
She|10714,10717
was|10718,10721
started|10722,10729
on|10730,10732
atorvastatin|10733,10745
<EOL>|10746,10747
for|10747,10750
her|10751,10754
hyperlipidemia|10755,10769
(|10770,10771
LDL|10771,10774
126|10775,10778
)|10778,10779
.|10779,10780
EP|10781,10783
cardiology|10784,10794
was|10795,10798
consulted|10799,10808
<EOL>|10809,10810
for|10810,10813
frequent|10814,10822
sinus|10823,10828
pauses|10829,10835
noted|10836,10841
on|10842,10844
telemetry|10845,10854
that|10855,10859
persisted|10860,10869
<EOL>|10870,10871
despite|10871,10878
holding|10879,10886
home|10887,10891
atenolol|10892,10900
,|10900,10901
recommending|10902,10914
discontinuing|10915,10928
home|10929,10933
<EOL>|10934,10935
digoxin|10935,10942
and|10943,10946
close|10947,10952
cardiology|10953,10963
_|10964,10965
_|10965,10966
_|10966,10967
.|10967,10968
Discharged|10969,10979
to|10980,10982
home|10983,10987
w|10988,10989
/|10989,10990
<EOL>|10991,10992
_|10992,10993
_|10993,10994
_|10994,10995
&|10996,10997
_|10998,10999
_|10999,11000
_|11000,11001
and|11002,11005
close|11006,11011
PCP|11012,11015
_|11016,11017
_|11017,11018
_|11018,11019
.|11019,11020
<EOL>|11020,11021
<EOL>|11021,11022
#|11022,11023
Transient|11023,11032
slurred|11033,11040
speech|11041,11047
and|11048,11051
instability|11052,11063
,|11063,11064
c|11065,11066
/|11066,11067
f|11067,11068
TIA|11069,11072
<EOL>|11072,11073
-|11073,11074
_|11075,11076
_|11076,11077
_|11077,11078
consult|11079,11086
-|11087,11088
cleared|11089,11096
for|11097,11100
home|11101,11105
with|11106,11110
home|11111,11115
services|11116,11124
<EOL>|11124,11125
-|11125,11126
Started|11127,11134
on|11135,11137
atorvastatin|11138,11150
for|11151,11154
HLD|11155,11158
and|11159,11162
increased|11163,11172
home|11173,11177
apixaban|11178,11186
to|11187,11189
<EOL>|11190,11191
therapeutic|11191,11202
level|11203,11208
<EOL>|11208,11209
-|11209,11210
_|11211,11212
_|11212,11213
_|11213,11214
with|11215,11219
stroke|11220,11226
neurology|11227,11236
after|11237,11242
discharge|11243,11252
<EOL>|11252,11253
<EOL>|11253,11254
Her|11254,11257
stroke|11258,11264
risk|11265,11269
factors|11270,11277
include|11278,11285
the|11286,11289
following|11290,11299
:|11299,11300
<EOL>|11300,11301
1|11301,11302
)|11302,11303
DM|11304,11306
:|11306,11307
A1c|11308,11311
5.5|11312,11315
%|11315,11316
<EOL>|11316,11317
2|11317,11318
)|11318,11319
Likely|11320,11326
chronic|11327,11334
segmental|11335,11344
left|11345,11349
vertebral|11350,11359
artery|11360,11366
occlusion|11367,11376
and|11377,11380
<EOL>|11381,11382
somewhat|11382,11390
small|11391,11396
caliber|11397,11404
attenuated|11405,11415
left|11416,11420
M2|11421,11423
inferior|11424,11432
branch|11433,11439
<EOL>|11439,11440
3|11440,11441
)|11441,11442
Hyperlipidemia|11443,11457
:|11457,11458
LDL|11459,11462
126|11463,11466
<EOL>|11466,11467
4|11467,11468
)|11468,11469
Obesity|11470,11477
<EOL>|11477,11478
5|11478,11479
)|11479,11480
No|11481,11483
concern|11484,11491
noted|11492,11497
for|11498,11501
sleep|11502,11507
apnea|11508,11513
-|11514,11515
she|11516,11519
does|11520,11524
not|11525,11528
carry|11529,11534
the|11535,11538
<EOL>|11539,11540
An|11550,11552
echocardiogram|11553,11567
did|11568,11571
not|11572,11575
show|11576,11580
a|11581,11582
PFO|11583,11586
on|11587,11589
bubble|11590,11596
study|11597,11602
.|11602,11603
<EOL>|11603,11604
<EOL>|11604,11605
AHA|11605,11608
/|11608,11609
ASA|11609,11612
Core|11613,11617
Measures|11618,11626
for|11627,11630
Ischemic|11631,11639
Stroke|11640,11646
and|11647,11650
Transient|11651,11660
Ischemic|11661,11669
<EOL>|11670,11671
Attack|11671,11677
<EOL>|11677,11678
1.|11678,11680
Dysphagia|11681,11690
screening|11691,11700
before|11701,11707
any|11708,11711
PO|11712,11714
intake|11715,11721
?|11721,11722
(|11723,11724
X|11724,11725
)|11725,11726
Yes|11727,11730
,|11730,11731
confirmed|11732,11741
<EOL>|11742,11743
done|11743,11747
-|11748,11749
(|11750,11751
)|11751,11752
Not|11753,11756
confirmed|11757,11766
(|11767,11768
)|11768,11769
No|11770,11772
<EOL>|11772,11773
2.|11773,11775
DVT|11776,11779
Prophylaxis|11780,11791
administered|11792,11804
?|11804,11805
(|11806,11807
X|11807,11808
)|11808,11809
Yes|11810,11813
-|11814,11815
(|11816,11817
)|11817,11818
No|11819,11821
<EOL>|11821,11822
3.|11822,11824
Antithrombotic|11825,11839
therapy|11840,11847
administered|11848,11860
by|11861,11863
end|11864,11867
of|11868,11870
hospital|11871,11879
day|11880,11883
2|11884,11885
?|11885,11886
<EOL>|11887,11888
(|11888,11889
X|11889,11890
)|11890,11891
Yes|11892,11895
-|11896,11897
(|11898,11899
)|11899,11900
No|11901,11903
<EOL>|11903,11904
4.|11904,11906
LDL|11907,11910
documented|11911,11921
?|11921,11922
(|11923,11924
X|11924,11925
)|11925,11926
Yes|11927,11930
(|11931,11932
LDL|11932,11935
=|11936,11937
126|11938,11941
)|11941,11942
-|11943,11944
(|11945,11946
)|11946,11947
No|11948,11950
<EOL>|11950,11951
5.|11951,11953
Intensive|11954,11963
statin|11964,11970
therapy|11971,11978
administered|11979,11991
?|11991,11992
(|11993,11994
simvastatin|11994,12005
80mg|12006,12010
,|12010,12011
<EOL>|12012,12013
simvastatin|12013,12024
80mg|12025,12029
/|12029,12030
ezetemibe|12030,12039
10mg|12040,12044
,|12044,12045
atorvastatin|12046,12058
40mg|12059,12063
or|12064,12066
80|12067,12069
mg|12070,12072
,|12072,12073
<EOL>|12074,12075
rosuvastatin|12075,12087
20mg|12088,12092
or|12093,12095
40mg|12096,12100
,|12100,12101
for|12102,12105
LDL|12106,12109
>|12110,12111
100|12112,12115
)|12115,12116
(|12117,12118
X|12118,12119
)|12119,12120
Yes|12121,12124
-|12125,12126
(|12127,12128
)|12128,12129
No|12130,12132
[|12133,12134
if|12134,12136
<EOL>|12137,12138
LDL|12138,12141
if|12142,12144
LDL|12145,12148
>|12149,12150
70|12150,12152
,|12152,12153
reason|12154,12160
not|12161,12164
given|12165,12170
:|12170,12171
<EOL>|12171,12172
[|12172,12173
]|12174,12175
Statin|12176,12182
medication|12183,12193
allergy|12194,12201
<EOL>|12201,12202
[|12202,12203
]|12204,12205
Other|12206,12211
reasons|12212,12219
documented|12220,12230
by|12231,12233
physician|12234,12243
/|12243,12244
advanced|12244,12252
practice|12253,12261
<EOL>|12262,12263
nurse|12263,12268
/|12268,12269
physician|12269,12278
_|12279,12280
_|12280,12281
_|12281,12282
(|12283,12284
physician|12284,12293
/|12293,12294
APN|12294,12297
/|12297,12298
PA|12298,12300
)|12300,12301
or|12302,12304
pharmacist|12305,12315
<EOL>|12315,12316
[|12316,12317
]|12318,12319
LDL|12320,12323
-|12323,12324
c|12324,12325
less|12326,12330
than|12331,12335
70|12336,12338
mg|12339,12341
/|12341,12342
dL|12342,12344
]|12344,12345
<EOL>|12345,12346
6.|12346,12348
Smoking|12349,12356
cessation|12357,12366
counseling|12367,12377
given|12378,12383
?|12383,12384
(|12385,12386
)|12386,12387
Yes|12388,12391
-|12392,12393
(|12394,12395
X|12395,12396
)|12396,12397
No|12398,12400
[|12401,12402
reason|12402,12408
<EOL>|12409,12410
(|12410,12411
X|12411,12412
)|12412,12413
non-smoker|12414,12424
-|12425,12426
(|12427,12428
)|12428,12429
unable|12430,12436
to|12437,12439
participate|12440,12451
]|12451,12452
<EOL>|12452,12453
7.|12453,12455
Stroke|12456,12462
education|12463,12472
(|12473,12474
personal|12474,12482
modifiable|12483,12493
risk|12494,12498
factors|12499,12506
,|12506,12507
how|12508,12511
to|12512,12514
<EOL>|12515,12516
activate|12516,12524
EMS|12525,12528
for|12529,12532
stroke|12533,12539
,|12539,12540
stroke|12541,12547
warning|12548,12555
signs|12556,12561
and|12562,12565
symptoms|12566,12574
,|12574,12575
<EOL>|12576,12577
prescribed|12577,12587
medications|12588,12599
,|12599,12600
need|12601,12605
for|12606,12609
followup|12610,12618
)|12618,12619
given|12620,12625
(|12626,12627
verbally|12627,12635
or|12636,12638
<EOL>|12639,12640
written|12640,12647
)|12647,12648
?|12648,12649
(|12650,12651
X|12651,12652
)|12652,12653
Yes|12654,12657
-|12658,12659
(|12660,12661
)|12661,12662
No|12663,12665
<EOL>|12665,12666
8.|12666,12668
Assessment|12669,12679
for|12680,12683
rehabilitation|12684,12698
or|12699,12701
rehab|12702,12707
services|12708,12716
considered|12717,12727
?|12727,12728
<EOL>|12729,12730
(|12730,12731
X|12731,12732
)|12732,12733
Yes|12734,12737
-|12738,12739
(|12740,12741
)|12741,12742
No|12743,12745
<EOL>|12745,12746
9.|12746,12748
Discharged|12749,12759
on|12760,12762
statin|12763,12769
therapy|12770,12777
?|12777,12778
(|12779,12780
X|12780,12781
)|12781,12782
Yes|12783,12786
-|12787,12788
(|12789,12790
)|12790,12791
No|12792,12794
[|12795,12796
if|12796,12798
LDL|12799,12802
>|12803,12804
70|12804,12806
,|12806,12807
<EOL>|12808,12809
reason|12809,12815
not|12816,12819
given|12820,12825
:|12825,12826
<EOL>|12826,12827
[|12827,12828
]|12829,12830
Statin|12831,12837
medication|12838,12848
allergy|12849,12856
<EOL>|12856,12857
[|12857,12858
]|12859,12860
Other|12861,12866
reasons|12867,12874
documented|12875,12885
by|12886,12888
physician|12889,12898
/|12898,12899
advanced|12899,12907
practice|12908,12916
<EOL>|12917,12918
nurse|12918,12923
/|12923,12924
physician|12924,12933
_|12934,12935
_|12935,12936
_|12936,12937
(|12938,12939
physician|12939,12948
/|12948,12949
APN|12949,12952
/|12952,12953
PA|12953,12955
)|12955,12956
or|12957,12959
pharmacist|12960,12970
<EOL>|12970,12971
[|12971,12972
]|12973,12974
LDL|12975,12978
-|12978,12979
c|12979,12980
less|12981,12985
than|12986,12990
70|12991,12993
mg|12994,12996
/|12996,12997
dL|12997,12999
<EOL>|12999,13000
10.|13000,13003
Discharged|13004,13014
on|13015,13017
antithrombotic|13018,13032
therapy|13033,13040
?|13040,13041
(|13042,13043
X|13043,13044
)|13044,13045
Yes|13046,13049
[|13050,13051
Type|13051,13055
:|13055,13056
(|13057,13058
)|13058,13059
<EOL>|13060,13061
Antiplatelet|13061,13073
-|13074,13075
(|13076,13077
X|13077,13078
)|13078,13079
Anticoagulation|13080,13095
]|13095,13096
-|13097,13098
(|13099,13100
)|13100,13101
No|13102,13104
<EOL>|13104,13105
11|13105,13107
.|13107,13108
Discharged|13109,13119
on|13120,13122
oral|13123,13127
anticoagulation|13128,13143
for|13144,13147
patients|13148,13156
with|13157,13161
atrial|13162,13168
<EOL>|13169,13170
fibrillation|13170,13182
/|13182,13183
flutter|13183,13190
?|13190,13191
(|13192,13193
X|13193,13194
)|13194,13195
Yes|13196,13199
-|13200,13201
(|13202,13203
)|13203,13204
No|13205,13207
-|13208,13209
(|13210,13211
)|13211,13212
N|13213,13214
/|13214,13215
A|13215,13216
<EOL>|13216,13217
<EOL>|13217,13218
#|13218,13219
Cognitive|13219,13228
complaints|13229,13239
<EOL>|13239,13240
-|13240,13241
B12|13242,13245
249|13246,13249
-|13250,13251
one|13252,13255
time|13256,13260
IM|13261,13263
supplementation|13264,13279
,|13279,13280
then|13281,13285
start|13286,13291
oral|13292,13296
B12|13297,13300
<EOL>|13301,13302
supplementation|13302,13317
<EOL>|13317,13318
-|13318,13319
Treponemal|13320,13330
antibodies|13331,13341
negative|13342,13350
<EOL>|13350,13351
-|13351,13352
consider|13353,13361
cognitive|13362,13371
neurology|13372,13381
referral|13382,13390
as|13391,13393
outpatient|13394,13404
for|13405,13408
memory|13409,13415
<EOL>|13416,13417
difficulties|13417,13429
not|13430,13433
appreciated|13434,13445
on|13446,13448
our|13449,13452
examination|13453,13464
<EOL>|13464,13465
<EOL>|13465,13466
#|13466,13467
Afib|13467,13471
<EOL>|13471,13472
#|13472,13473
frequent|13473,13481
sinus|13482,13487
pauses|13488,13494
<EOL>|13494,13495
-|13495,13496
stopped|13497,13504
digoxin|13505,13512
,|13512,13513
will|13514,13518
_|13519,13520
_|13520,13521
_|13521,13522
closely|13523,13530
w|13531,13532
/|13532,13533
otpt|13534,13538
cardiologist|13539,13551
<EOL>|13552,13553
(|13553,13554
also|13554,13558
PCP|13559,13562
)|13562,13563
<EOL>|13563,13564
-|13564,13565
increased|13566,13575
to|13576,13578
appropriate|13579,13590
therapeutic|13591,13602
dosing|13603,13609
at|13610,13612
Eliquis|13613,13620
2.5|13621,13624
mg|13625,13627
<EOL>|13628,13629
BID|13629,13632
(|13633,13634
reduced|13634,13641
dose|13642,13646
given|13647,13652
age|13653,13656
and|13657,13660
weight|13661,13667
<|13668,13669
60|13669,13671
kg|13672,13674
)|13674,13675
<EOL>|13675,13676
<EOL>|13676,13677
#|13677,13678
HLD|13678,13681
<EOL>|13681,13682
-|13682,13683
started|13684,13691
atorvastatin|13692,13704
<EOL>|13704,13705
<EOL>|13705,13706
#|13706,13707
HTN|13707,13710
<EOL>|13710,13711
-|13711,13712
continue|13713,13721
home|13722,13726
antihypertensives|13727,13744
<EOL>|13744,13745
<EOL>|13745,13746
#|13746,13747
elevated|13747,13755
troponin|13756,13764
(|13765,13766
RESOLVED|13766,13774
)|13774,13775
<EOL>|13775,13776
-|13776,13777
Troponin|13778,13786
elevated|13787,13795
at|13796,13798
OSH|13799,13802
,|13802,13803
negative|13804,13812
on|13813,13815
admission|13816,13825
<EOL>|13825,13826
<EOL>|13826,13827
#|13827,13828
elevated|13828,13836
TSH|13837,13840
<EOL>|13840,13841
-|13841,13842
should|13843,13849
recheck|13850,13857
as|13858,13860
otpt|13861,13865
w|13866,13867
/|13867,13868
PCP|13869,13872
_|13873,13874
_|13874,13875
_|13875,13876
<EOL>|13876,13877
<EOL>|13878,13879
Medications|13879,13890
on|13891,13893
Admission|13894,13903
:|13903,13904
<EOL>|13904,13905
The|13905,13908
Preadmission|13909,13921
Medication|13922,13932
list|13933,13937
is|13938,13940
accurate|13941,13949
and|13950,13953
complete|13954,13962
.|13962,13963
<EOL>|13963,13964
1.|13964,13966
Atenolol|13967,13975
50|13976,13978
mg|13979,13981
PO|13982,13984
DAILY|13985,13990
<EOL>|13991,13992
2.|13992,13994
Apixaban|13995,14003
2.5|14004,14007
mg|14008,14010
PO|14011,14013
DAILY|14014,14019
<EOL>|14020,14021
3.|14021,14023
Losartan|14024,14032
Potassium|14033,14042
50|14043,14045
mg|14046,14048
PO|14049,14051
DAILY|14052,14057
<EOL>|14058,14059
4.|14059,14061
Digoxin|14062,14069
0.125|14070,14075
mg|14076,14078
PO|14079,14081
DAILY|14082,14087
<EOL>|14088,14089
5.|14089,14091
LevoFLOXacin|14092,14104
500|14105,14108
mg|14109,14111
PO|14112,14114
Q24H|14115,14119
<EOL>|14120,14121
<EOL>|14121,14122
<EOL>|14123,14124
Discharge|14124,14133
Medications|14134,14145
:|14145,14146
<EOL>|14146,14147
1.|14147,14149
Atorvastatin|14151,14163
40|14164,14166
mg|14167,14169
PO|14170,14172
QPM|14173,14176
<EOL>|14177,14178
RX|14178,14180
*|14181,14182
atorvastatin|14182,14194
40|14195,14197
mg|14198,14200
1|14201,14202
tablet|14203,14209
(|14209,14210
s|14210,14211
)|14211,14212
by|14213,14215
mouth|14216,14221
once|14222,14226
daily|14227,14232
at|14233,14235
<EOL>|14236,14237
bedtime|14237,14244
Disp|14245,14249
#|14250,14251
*|14251,14252
30|14252,14254
Tablet|14255,14261
Refills|14262,14269
:|14269,14270
*|14270,14271
5|14271,14272
<EOL>|14273,14274
2.|14274,14276
Cyanocobalamin|14278,14292
500|14293,14296
mcg|14297,14300
PO|14301,14303
DAILY|14304,14309
<EOL>|14310,14311
RX|14311,14313
*|14314,14315
cyanocobalamin|14315,14329
(|14330,14331
vitamin|14331,14338
B|14339,14340
-|14340,14341
12|14341,14343
)|14343,14344
500|14345,14348
mcg|14349,14352
1|14353,14354
tablet|14355,14361
(|14361,14362
s|14362,14363
)|14363,14364
by|14365,14367
mouth|14368,14373
<EOL>|14374,14375
once|14375,14379
daily|14380,14385
Disp|14386,14390
#|14391,14392
*|14392,14393
30|14393,14395
Tablet|14396,14402
Refills|14403,14410
:|14410,14411
*|14411,14412
5|14412,14413
<EOL>|14414,14415
3.|14415,14417
Apixaban|14419,14427
2.5|14428,14431
mg|14432,14434
PO|14435,14437
BID|14438,14441
<EOL>|14443,14444
4.|14444,14446
Atenolol|14448,14456
50|14457,14459
mg|14460,14462
PO|14463,14465
DAILY|14466,14471
<EOL>|14473,14474
5.|14474,14476
LevoFLOXacin|14478,14490
500|14491,14494
mg|14495,14497
PO|14498,14500
Q24H|14501,14505
<EOL>|14507,14508
6.|14508,14510
Losartan|14512,14520
Potassium|14521,14530
50|14531,14533
mg|14534,14536
PO|14537,14539
DAILY|14540,14545
<EOL>|14547,14548
<EOL>|14548,14549
<EOL>|14550,14551
Discharge|14551,14560
Disposition|14561,14572
:|14572,14573
<EOL>|14573,14574
Home|14574,14578
With|14579,14583
Service|14584,14591
<EOL>|14591,14592
<EOL>|14593,14594
Facility|14594,14602
:|14602,14603
<EOL>|14603,14604
_|14604,14605
_|14605,14606
_|14606,14607
<EOL>|14607,14608
<EOL>|14609,14610
Discharge|14610,14619
Diagnosis|14620,14629
:|14629,14630
<EOL>|14630,14631
transient|14631,14640
dysarthria|14641,14651
not|14652,14655
secondary|14656,14665
to|14666,14668
TIA|14669,14672
or|14673,14675
stroke|14676,14682
<EOL>|14682,14683
Mild|14683,14687
Vitamin|14688,14695
B12|14696,14699
deficiency|14700,14710
<EOL>|14710,14711
<EOL>|14712,14713
Mental|14734,14740
Status|14741,14747
:|14747,14748
Clear|14749,14754
and|14755,14758
coherent|14759,14767
.|14767,14768
<EOL>|14768,14769
Level|14769,14774
of|14775,14777
Consciousness|14778,14791
:|14791,14792
Alert|14793,14798
and|14799,14802
interactive|14803,14814
.|14814,14815
<EOL>|14815,14816
Activity|14816,14824
Status|14825,14831
:|14831,14832
Ambulatory|14833,14843
-|14844,14845
requires|14846,14854
assistance|14855,14865
or|14866,14868
aid|14869,14872
(|14873,14874
walker|14874,14880
<EOL>|14881,14882
or|14882,14884
cane|14885,14889
)|14889,14890
.|14890,14891
<EOL>|14891,14892
<EOL>|14893,14894
Dear|14918,14922
Ms.|14923,14926
_|14927,14928
_|14928,14929
_|14929,14930
,|14930,14931
<EOL>|14931,14932
<EOL>|14932,14933
You|14933,14936
were|14937,14941
hospitalized|14942,14954
due|14955,14958
to|14959,14961
symptoms|14962,14970
of|14971,14973
slurred|14974,14981
speech|14982,14988
due|14989,14992
to|14993,14995
<EOL>|14996,14997
concern|14997,15004
for|15005,15008
an|15009,15011
ACUTE|15012,15017
ISCHEMIC|15018,15026
STROKE|15027,15033
,|15033,15034
a|15035,15036
condition|15037,15046
where|15047,15052
a|15053,15054
blood|15055,15060
<EOL>|15061,15062
vessel|15062,15068
providing|15069,15078
oxygen|15079,15085
and|15086,15089
nutrients|15090,15099
to|15100,15102
the|15103,15106
brain|15107,15112
is|15113,15115
blocked|15116,15123
by|15124,15126
<EOL>|15127,15128
a|15128,15129
clot|15130,15134
.|15134,15135
The|15136,15139
brain|15140,15145
is|15146,15148
the|15149,15152
part|15153,15157
of|15158,15160
your|15161,15165
body|15166,15170
that|15171,15175
controls|15176,15184
and|15185,15188
<EOL>|15189,15190
directs|15190,15197
all|15198,15201
the|15202,15205
other|15206,15211
parts|15212,15217
of|15218,15220
your|15221,15225
body|15226,15230
,|15230,15231
so|15232,15234
damage|15235,15241
to|15242,15244
the|15245,15248
brain|15249,15254
<EOL>|15255,15256
from|15256,15260
being|15261,15266
deprived|15267,15275
of|15276,15278
its|15279,15282
blood|15283,15288
supply|15289,15295
can|15296,15299
result|15300,15306
in|15307,15309
a|15310,15311
variety|15312,15319
<EOL>|15320,15321
of|15321,15323
symptoms|15324,15332
.|15332,15333
However|15334,15341
,|15341,15342
the|15343,15346
MRI|15347,15350
of|15351,15353
your|15354,15358
brain|15359,15364
did|15365,15368
not|15369,15372
show|15373,15377
<EOL>|15378,15379
evidence|15379,15387
of|15388,15390
stroke|15391,15397
or|15398,15400
TIA|15401,15404
.|15404,15405
Your|15406,15410
symptoms|15411,15419
could|15420,15425
have|15426,15430
been|15431,15435
related|15436,15443
<EOL>|15444,15445
to|15445,15447
blood|15448,15453
pressure|15454,15462
,|15462,15463
dehydration|15464,15475
,|15475,15476
alcohol|15477,15484
use|15485,15488
,|15488,15489
or|15490,15492
a|15493,15494
combination|15495,15506
of|15507,15509
<EOL>|15510,15511
these|15511,15516
factors|15517,15524
.|15524,15525
<EOL>|15525,15526
<EOL>|15526,15527
We|15527,15529
are|15530,15533
changing|15534,15542
your|15543,15547
medications|15548,15559
as|15560,15562
follows|15563,15570
:|15570,15571
<EOL>|15571,15572
Increase|15572,15580
apixaban|15581,15589
to|15590,15592
2.5|15593,15596
mg|15596,15598
twice|15599,15604
daily|15605,15610
<EOL>|15610,15611
Start|15611,15616
Vitamin|15617,15624
B12|15625,15628
daily|15629,15634
supplement|15635,15645
<EOL>|15645,15646
<EOL>|15646,15647
Please|15647,15653
take|15654,15658
your|15659,15663
other|15664,15669
medications|15670,15681
as|15682,15684
prescribed|15685,15695
.|15695,15696
<EOL>|15696,15697
<EOL>|15697,15698
Please|15698,15704
follow|15705,15711
up|15712,15714
with|15715,15719
your|15720,15724
primary|15725,15732
care|15733,15737
physician|15738,15747
as|15748,15750
listed|15751,15757
<EOL>|15758,15759
below|15759,15764
.|15764,15765
You|15766,15769
should|15770,15776
also|15777,15781
follow|15782,15788
up|15789,15791
with|15792,15796
your|15797,15801
cardiologist|15802,15814
as|15815,15817
you|15818,15821
<EOL>|15822,15823
were|15823,15827
noted|15828,15833
to|15834,15836
have|15837,15841
occasional|15842,15852
pauses|15853,15859
on|15860,15862
cardiac|15863,15870
monitoring|15871,15881
.|15881,15882
<EOL>|15882,15883
<EOL>|15883,15884
If|15884,15886
you|15887,15890
experience|15891,15901
any|15902,15905
of|15906,15908
the|15909,15912
symptoms|15913,15921
below|15922,15927
,|15927,15928
please|15929,15935
seek|15936,15940
<EOL>|15941,15942
emergency|15942,15951
medical|15952,15959
attention|15960,15969
by|15970,15972
calling|15973,15980
Emergency|15981,15990
Medical|15991,15998
<EOL>|15999,16000
Services|16000,16008
(|16009,16010
dialing|16010,16017
911|16018,16021
)|16021,16022
.|16022,16023
In|16024,16026
particular|16027,16037
,|16037,16038
please|16039,16045
pay|16046,16049
attention|16050,16059
to|16060,16062
<EOL>|16063,16064
the|16064,16067
sudden|16068,16074
onset|16075,16080
and|16081,16084
persistence|16085,16096
of|16097,16099
these|16100,16105
symptoms|16106,16114
:|16114,16115
<EOL>|16115,16116
-|16116,16117
Sudden|16118,16124
partial|16125,16132
or|16133,16135
complete|16136,16144
loss|16145,16149
of|16150,16152
vision|16153,16159
<EOL>|16159,16160
-|16160,16161
Sudden|16162,16168
loss|16169,16173
of|16174,16176
the|16177,16180
ability|16181,16188
to|16189,16191
speak|16192,16197
words|16198,16203
from|16204,16208
your|16209,16213
mouth|16214,16219
<EOL>|16219,16220
-|16220,16221
Sudden|16222,16228
loss|16229,16233
of|16234,16236
the|16237,16240
ability|16241,16248
to|16249,16251
understand|16252,16262
others|16263,16269
speaking|16270,16278
to|16279,16281
<EOL>|16282,16283
you|16283,16286
<EOL>|16286,16287
-|16287,16288
Sudden|16289,16295
weakness|16296,16304
of|16305,16307
one|16308,16311
side|16312,16316
of|16317,16319
the|16320,16323
body|16324,16328
<EOL>|16328,16329
-|16329,16330
Sudden|16331,16337
drooping|16338,16346
of|16347,16349
one|16350,16353
side|16354,16358
of|16359,16361
the|16362,16365
face|16366,16370
<EOL>|16370,16371
-|16371,16372
Sudden|16373,16379
loss|16380,16384
of|16385,16387
sensation|16388,16397
of|16398,16400
one|16401,16404
side|16405,16409
of|16410,16412
the|16413,16416
body|16417,16421
<EOL>|16421,16422
<EOL>|16422,16423
Sincerely|16423,16432
,|16432,16433
<EOL>|16433,16434
Your|16434,16438
_|16439,16440
_|16440,16441
_|16441,16442
Neurology|16443,16452
Team|16453,16457
<EOL>|16457,16458
<EOL>|16459,16460
Followup|16460,16468
Instructions|16469,16481
:|16481,16482
<EOL>|16482,16483
_|16483,16484
_|16484,16485
_|16485,16486
<EOL>|16486,16487

