 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|SIMPLE_SEGMENT|168,177|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|168,177|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|168,177|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Antibiotic|SIMPLE_SEGMENT|180,191|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|180,191|false|false|false|C0002645|amoxicillin|amoxicillin
Event|Event|SIMPLE_SEGMENT|180,191|false|false|false|||amoxicillin
Event|Event|SIMPLE_SEGMENT|194,203|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|194,203|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|212,227|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|218,227|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|218,227|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|218,227|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|229,237|false|false|false|||Weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|229,237|false|false|false|C0004093;C3714552|Asthenia;Weakness|Weakness
Event|Event|SIMPLE_SEGMENT|242,250|false|false|false|||lethargy
Finding|Sign or Symptom|SIMPLE_SEGMENT|242,250|false|false|false|C0023380|Lethargy|lethargy
Finding|Classification|SIMPLE_SEGMENT|254,259|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|260,268|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|272,290|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|281,290|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|281,290|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|281,290|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|281,290|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|281,290|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|300,307|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|300,307|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|300,307|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|300,307|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|300,310|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|300,326|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|300,326|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|311,318|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|311,318|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|311,326|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|319,326|false|false|false|C0221423|Illness (finding)|Illness
Finding|Body Substance|SIMPLE_SEGMENT|328,335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|328,335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|328,335|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|345,349|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|SIMPLE_SEGMENT|345,349|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|SIMPLE_SEGMENT|350,353|false|false|false|||old
Event|Event|SIMPLE_SEGMENT|366,373|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|366,376|false|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|377,384|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|377,384|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|377,384|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Location or Region|SIMPLE_SEGMENT|385,394|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|385,399|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|395,399|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|395,399|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|395,399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|395,399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|404,410|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|404,410|false|false|false|||anemia
Drug|Biologically Active Substance|SIMPLE_SEGMENT|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Drug|Organic Chemical|SIMPLE_SEGMENT|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|424,431|false|false|false|C0038636;C1161331|Saccharum officinale, sucrose, cane sugar, Homeopathic preparation;sucrose|sucrose
Event|Event|SIMPLE_SEGMENT|432,440|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|432,440|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|432,440|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|447,458|false|false|false|||complicated
Finding|Functional Concept|SIMPLE_SEGMENT|462,470|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|462,470|false|false|false|C0574032|Infusion procedures|infusion
Finding|Pathologic Function|SIMPLE_SEGMENT|462,479|false|false|false|C2368034|Infusion reaction|infusion reaction
Event|Event|SIMPLE_SEGMENT|471,479|false|false|false|||reaction
Finding|Functional Concept|SIMPLE_SEGMENT|471,479|false|false|false|C0443286|Reaction|reaction
Event|Event|SIMPLE_SEGMENT|481,489|false|false|false|||mottling
Finding|Finding|SIMPLE_SEGMENT|481,489|false|false|false|C0302133|Mottling|mottling
Event|Event|SIMPLE_SEGMENT|494,507|false|false|false|||discoloration
Finding|Finding|SIMPLE_SEGMENT|494,507|false|false|false|C0332572|Abnormal color|discoloration
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|511,515|false|false|false|C0016504|Foot|feet
Drug|Organic Chemical|SIMPLE_SEGMENT|524,532|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|524,532|false|false|false|C0038317|Steroids|steroids
Event|Event|SIMPLE_SEGMENT|524,532|false|false|false|||steroids
Event|Event|SIMPLE_SEGMENT|537,545|false|false|false|||presents
Event|Event|SIMPLE_SEGMENT|562,570|false|false|false|||lethargy
Finding|Sign or Symptom|SIMPLE_SEGMENT|562,570|false|false|false|C0023380|Lethargy|lethargy
Event|Event|SIMPLE_SEGMENT|575,583|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|575,583|false|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|586,593|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|586,593|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|602,609|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|602,609|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|602,609|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|SIMPLE_SEGMENT|622,626|false|false|false|||Aunt
Finding|Body Substance|SIMPLE_SEGMENT|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|630,637|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|645,652|false|false|false|||provide
Finding|Finding|SIMPLE_SEGMENT|653,657|false|false|false|C4281574|Much|much
Event|Event|SIMPLE_SEGMENT|658,665|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|658,665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|658,665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|658,665|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|700,704|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|700,704|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|726,733|false|false|false|||illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|726,733|true|false|false|C0221423|Illness (finding)|illness
Finding|Behavior|SIMPLE_SEGMENT|735,745|false|false|false|C0004927|Behavior|behavioral
Finding|Individual Behavior|SIMPLE_SEGMENT|735,752|false|false|false|C0542299|Behavioral change|behavioral change
Event|Event|SIMPLE_SEGMENT|746,752|false|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|746,752|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|746,752|false|false|false|C4319952|Change - procedure|change
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|764,768|false|false|false|C0009443;C0024117|Chronic Obstructive Airway Disease;Common Cold|cold
Drug|Organic Chemical|SIMPLE_SEGMENT|764,768|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|764,768|false|false|false|C0719425|Cold brand of chlorpheniramine-phenylpropanolamine|cold
Event|Event|SIMPLE_SEGMENT|764,768|false|false|false|||cold
Finding|Organism Function|SIMPLE_SEGMENT|764,768|false|false|false|C0234192|Cold Sensation|cold
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|764,768|false|false|false|C0009264|Cold Temperature|cold
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|764,768|false|false|false|C0010412|Cold Therapy|cold
Event|Event|SIMPLE_SEGMENT|777,784|false|false|false|||getting
Event|Event|SIMPLE_SEGMENT|810,814|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|810,814|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|830,841|false|false|false|||transfusion
Finding|Functional Concept|SIMPLE_SEGMENT|830,841|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|830,841|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Event|SIMPLE_SEGMENT|882,893|false|false|false|||accompanied
Event|Event|SIMPLE_SEGMENT|905,910|false|false|false|||visit
Finding|Social Behavior|SIMPLE_SEGMENT|905,910|false|false|false|C0545082|Visit|visit
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|924,927|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|SIMPLE_SEGMENT|924,927|false|false|false|C0082420|Endoglin, human|end
Event|Event|SIMPLE_SEGMENT|924,927|false|false|false|||end
Finding|Functional Concept|SIMPLE_SEGMENT|924,927|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|SIMPLE_SEGMENT|924,927|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Event|Event|SIMPLE_SEGMENT|935,943|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|935,943|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|935,943|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|949,958|false|false|false|||developed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|973,978|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|973,978|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|973,990|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|979,990|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1006,1012|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1006,1012|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1006,1012|false|false|false|C0027497|Nausea|nausea
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1014,1019|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1014,1019|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1014,1019|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Finding|SIMPLE_SEGMENT|1014,1026|false|false|false|C0039231|Tachycardia|heart racing
Event|Event|SIMPLE_SEGMENT|1020,1026|false|false|false|||racing
Finding|Intellectual Product|SIMPLE_SEGMENT|1020,1026|false|false|false|C1561444|Racing - Production Class Code|racing
Event|Event|SIMPLE_SEGMENT|1036,1040|false|false|false|||sent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1062,1065|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1062,1065|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1062,1065|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|1062,1065|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|1062,1065|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1062,1065|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|SIMPLE_SEGMENT|1081,1085|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|1081,1085|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1081,1085|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|1094,1101|false|false|false|||records
Finding|Idea or Concept|SIMPLE_SEGMENT|1094,1101|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|SIMPLE_SEGMENT|1094,1101|false|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Event|Event|SIMPLE_SEGMENT|1115,1124|false|false|false|||shivering
Finding|Finding|SIMPLE_SEGMENT|1115,1124|false|false|false|C0036973|Shivering|shivering
Event|Event|SIMPLE_SEGMENT|1136,1140|false|false|false|||open
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1145,1149|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1145,1149|false|false|false|C5848506||eyes
Finding|Finding|SIMPLE_SEGMENT|1152,1159|false|false|false|C0302133|Mottling|mottled
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1160,1165|false|false|false|C0018563|Hand|hands
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1170,1174|false|false|false|C0016504|Foot|feet
Event|Event|SIMPLE_SEGMENT|1190,1197|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|1190,1197|false|false|false|C2699424|Concern|concern
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1202,1213|false|false|false|C0231832|Respiratory rate|respiratory
Finding|Body Substance|SIMPLE_SEGMENT|1202,1213|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Functional Concept|SIMPLE_SEGMENT|1202,1213|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Intellectual Product|SIMPLE_SEGMENT|1202,1213|false|false|false|C0521346;C1314992;C1546767;C5442009|Respiratory attachment;Respiratory specimen;respiratory|respiratory
Finding|Sign or Symptom|SIMPLE_SEGMENT|1202,1222|false|false|false|C0476273|Respiratory distress|respiratory distress
Event|Event|SIMPLE_SEGMENT|1214,1222|false|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|1214,1222|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|1214,1222|false|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Event|Event|SIMPLE_SEGMENT|1232,1237|false|false|false|||given
Drug|Organic Chemical|SIMPLE_SEGMENT|1247,1255|false|false|false|C0700899|Benadryl|Benadryl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1247,1255|false|false|false|C0700899|Benadryl|Benadryl
Drug|Hormone|SIMPLE_SEGMENT|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Drug|Organic Chemical|SIMPLE_SEGMENT|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1267,1281|false|false|false|C0020268|hydrocortisone|hydrocortisone
Event|Event|SIMPLE_SEGMENT|1267,1281|false|false|false|||hydrocortisone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1267,1281|false|false|false|C0201968|Cortisol Measurement|hydrocortisone
Event|Event|SIMPLE_SEGMENT|1286,1294|false|false|false|||observed
Finding|Intellectual Product|SIMPLE_SEGMENT|1311,1315|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|1316,1326|false|false|false|||discharged
Finding|Finding|SIMPLE_SEGMENT|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1336,1340|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|1361,1370|false|false|false|||lethargic
Finding|Sign or Symptom|SIMPLE_SEGMENT|1361,1370|false|false|false|C0023380|Lethargy|lethargic
Event|Event|SIMPLE_SEGMENT|1372,1379|false|false|false|||meaning
Event|Event|SIMPLE_SEGMENT|1380,1388|false|false|false|||sleeping
Event|Event|SIMPLE_SEGMENT|1404,1408|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1404,1408|false|false|false|C1299581|Able (qualifier value)|able
Finding|Finding|SIMPLE_SEGMENT|1404,1415|false|false|false|C0560880|Able to sit|able to sit
Finding|Finding|SIMPLE_SEGMENT|1404,1418|false|false|false|C0560835|Able to sit up|able to sit up
Finding|Finding|SIMPLE_SEGMENT|1412,1415|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Gene or Genome|SIMPLE_SEGMENT|1412,1415|false|false|false|C0277814;C0728713;C1539668;C1539774|Does sit;HHAT gene;SIT1 gene;Sitting position|sit
Finding|Finding|SIMPLE_SEGMENT|1412,1418|false|false|false|C0560837|Does sit up|sit up
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1423,1427|false|false|false|C0080331|Walking (function)|walk
Event|Activity|SIMPLE_SEGMENT|1436,1441|false|false|false|C5966184|Issue (action)|issue
Event|Event|SIMPLE_SEGMENT|1436,1441|false|false|false|||issue
Finding|Finding|SIMPLE_SEGMENT|1436,1441|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|SIMPLE_SEGMENT|1436,1441|false|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|SIMPLE_SEGMENT|1448,1455|false|false|false|||arrived
Event|Event|SIMPLE_SEGMENT|1456,1460|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|1456,1460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|1456,1460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|1456,1460|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|1469,1473|false|false|false|||went
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1477,1480|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|1477,1480|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|1477,1480|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|1494,1496|false|false|false|||AM
Event|Event|SIMPLE_SEGMENT|1514,1519|false|false|false|||check
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1539,1544|false|false|false|C1410088|Still|still
Event|Event|SIMPLE_SEGMENT|1545,1553|false|false|false|||sleeping
Event|Event|SIMPLE_SEGMENT|1563,1572|false|false|false|||reporting
Event|Event|SIMPLE_SEGMENT|1575,1583|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|1575,1583|false|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|1595,1606|false|false|false|||transfusion
Finding|Functional Concept|SIMPLE_SEGMENT|1595,1606|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1595,1606|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Event|Activity|SIMPLE_SEGMENT|1607,1612|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|1607,1612|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|1607,1612|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|1607,1612|false|false|false|C1533810||place
Event|Event|SIMPLE_SEGMENT|1613,1617|false|false|false|||said
Event|Event|SIMPLE_SEGMENT|1624,1630|false|false|false|||happen
Event|Event|SIMPLE_SEGMENT|1644,1651|false|false|false|||mention
Event|Event|SIMPLE_SEGMENT|1658,1672|false|false|false|||characteristic
Event|Event|SIMPLE_SEGMENT|1684,1688|false|false|false|||gave
Drug|Organic Chemical|SIMPLE_SEGMENT|1693,1706|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1693,1706|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|SIMPLE_SEGMENT|1693,1706|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1693,1706|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Inorganic Chemical|SIMPLE_SEGMENT|1711,1716|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1711,1716|false|false|false|C0043047;C1550678|Water Specimen;water|water
Event|Event|SIMPLE_SEGMENT|1711,1716|false|false|false|||water
Finding|Intellectual Product|SIMPLE_SEGMENT|1711,1716|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1711,1716|false|false|false|C0020311|Hydrotherapy|water
Event|Event|SIMPLE_SEGMENT|1725,1729|false|false|false|||went
Drug|Organic Chemical|SIMPLE_SEGMENT|1738,1743|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1738,1743|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|SIMPLE_SEGMENT|1738,1743|false|false|false|||sleep
Finding|Organism Function|SIMPLE_SEGMENT|1738,1743|false|false|false|C0037313|Sleep|sleep
Finding|Idea or Concept|SIMPLE_SEGMENT|1754,1758|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|SIMPLE_SEGMENT|1774,1779|false|false|false|||heard
Finding|Finding|SIMPLE_SEGMENT|1784,1789|false|false|false|C0234422|Awake (finding)|awake
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1798,1803|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|1798,1803|false|false|false|||times
Event|Event|SIMPLE_SEGMENT|1808,1811|false|false|false|||use
Event|Event|SIMPLE_SEGMENT|1816,1824|false|false|false|||bathroom
Finding|Intellectual Product|SIMPLE_SEGMENT|1826,1830|false|false|false|C1720594|Then - dosing instruction fragment|Then
Event|Event|SIMPLE_SEGMENT|1837,1840|false|false|false|||got
Finding|Idea or Concept|SIMPLE_SEGMENT|1866,1869|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1866,1869|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1913,1919|false|false|false|||became
Event|Event|SIMPLE_SEGMENT|1920,1927|false|false|false|||worried
Finding|Finding|SIMPLE_SEGMENT|1920,1927|false|false|false|C0233481|Worried|worried
Event|Event|SIMPLE_SEGMENT|1933,1937|false|false|false|||told
Event|Event|SIMPLE_SEGMENT|1972,1976|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|1972,1976|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|1980,1982|false|false|false|||do
Event|Event|SIMPLE_SEGMENT|1999,2003|false|false|false|||said
Event|Event|SIMPLE_SEGMENT|2008,2017|false|false|false|||continued
Event|Event|SIMPLE_SEGMENT|2028,2036|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|2028,2036|false|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|2041,2045|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|2046,2052|false|false|false|||sleepy
Finding|Finding|SIMPLE_SEGMENT|2046,2052|false|false|false|C0013144|Drowsiness|sleepy
Event|Event|SIMPLE_SEGMENT|2062,2072|false|false|false|||instructed
Event|Event|SIMPLE_SEGMENT|2076,2078|false|false|false|||go
Event|Event|SIMPLE_SEGMENT|2096,2100|false|false|false|||went
Event|Event|SIMPLE_SEGMENT|2122,2132|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|2122,2132|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2122,2132|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|2213,2219|false|false|false|||drowsy
Finding|Finding|SIMPLE_SEGMENT|2213,2219|false|false|false|C0013144|Drowsiness|drowsy
Event|Event|SIMPLE_SEGMENT|2236,2241|false|false|false|||voice
Finding|Idea or Concept|SIMPLE_SEGMENT|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|SIMPLE_SEGMENT|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|SIMPLE_SEGMENT|2236,2241|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2244,2249|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2244,2249|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2244,2249|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|2244,2249|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2244,2249|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Finding|SIMPLE_SEGMENT|2250,2258|false|false|false|C1961028|Oriented to place|oriented
Event|Event|SIMPLE_SEGMENT|2259,2261|false|false|false|||x3
Finding|Idea or Concept|SIMPLE_SEGMENT|2264,2274|false|false|false|C0332290|Consistent with|consistent
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2275,2278|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2275,2278|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2275,2278|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2275,2278|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|2275,2278|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Event|Event|SIMPLE_SEGMENT|2279,2289|false|false|false|||fluttering
Finding|Pathologic Function|SIMPLE_SEGMENT|2279,2289|false|false|false|C0016385|Cardiac Flutter|fluttering
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2291,2297|false|false|false|C0034121|Pupil|pupils
Event|Event|SIMPLE_SEGMENT|2298,2306|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2298,2306|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|SIMPLE_SEGMENT|2298,2315|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2310,2315|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2310,2315|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|SIMPLE_SEGMENT|2310,2315|false|false|false|||light
Finding|Finding|SIMPLE_SEGMENT|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|2310,2315|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2310,2315|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2310,2315|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|SIMPLE_SEGMENT|2320,2331|false|false|false|C0241886|Extraocular|extraocular
Finding|Finding|SIMPLE_SEGMENT|2320,2345|false|false|false|C0702182|Extraocular eye movement|extraocular eye movements
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2332,2335|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2332,2335|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2332,2335|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2332,2335|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|2332,2335|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Physiologic Function|SIMPLE_SEGMENT|2332,2345|false|false|false|C0015413|Eye Movements|eye movements
Event|Event|SIMPLE_SEGMENT|2336,2345|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|2336,2345|false|false|false|C0026649|Movement|movements
Event|Event|SIMPLE_SEGMENT|2346,2350|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|2380,2384|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|2380,2384|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2380,2384|false|false|false|C0582103|Medical Examination|exam
Finding|Gene or Genome|SIMPLE_SEGMENT|2387,2390|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|SIMPLE_SEGMENT|2387,2390|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Event|SIMPLE_SEGMENT|2391,2395|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|2391,2395|false|false|false|C0043227|Work|work
Anatomy|Cell|SIMPLE_SEGMENT|2408,2411|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2417,2420|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2417,2420|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|2417,2420|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|2417,2420|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2417,2420|false|false|false|C0019029|Hemoglobin concentration|Hgb
Drug|Organic Chemical|SIMPLE_SEGMENT|2435,2441|false|false|false|C0074722|sodium bicarbonate|bicarb
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2435,2441|false|false|false|C0074722|sodium bicarbonate|bicarb
Event|Event|SIMPLE_SEGMENT|2435,2441|false|false|false|||bicarb
Event|Event|SIMPLE_SEGMENT|2469,2473|false|false|false|||LFTs
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2483,2491|false|false|false|C0015879|Ferritin|Ferritin
Event|Event|SIMPLE_SEGMENT|2483,2491|false|false|false|||Ferritin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2483,2491|false|false|false|C0373607|Ferritin measurement|Ferritin
Event|Event|SIMPLE_SEGMENT|2501,2503|false|false|false|||pH
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2514,2518|false|false|false|C0391839|Carbon dioxide, partial pressure|PCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2514,2518|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|PCO2
Anatomy|Cell|SIMPLE_SEGMENT|2559,2562|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|2571,2580|false|false|false|C0026473|Monocytes|monocytes
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2581,2588|false|false|false|C0017725|glucose|glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|2581,2588|false|false|false|C0017725|glucose|glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2581,2588|false|false|false|C0017725|glucose|glucose
Event|Event|SIMPLE_SEGMENT|2581,2588|false|false|false|||glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2581,2588|false|false|false|C5781949|Glucose^1.5H post dose glucagon|glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2581,2588|false|false|false|C0337438|Glucose measurement|glucose
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2593,2600|false|false|false|C0033684|Proteins|protein
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2593,2600|false|false|false|C0033684|Proteins|protein
Event|Event|SIMPLE_SEGMENT|2593,2600|false|false|false|||protein
Finding|Conceptual Entity|SIMPLE_SEGMENT|2593,2600|false|false|false|C1521746|Protein Info|protein
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2593,2600|false|false|false|C0202202|Protein measurement|protein
Event|Event|SIMPLE_SEGMENT|2608,2621|false|false|false|||xanthochromia
Finding|Finding|SIMPLE_SEGMENT|2608,2621|true|false|false|C0863146|Yellow color (finding)|xanthochromia
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2642,2645|false|false|false|C1609165|tocilizumab|MRA
Event|Event|SIMPLE_SEGMENT|2642,2645|false|false|false|||MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2642,2645|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2642,2645|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|2650,2653|false|false|false|C0876081|MRV|MRV
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2650,2653|false|false|false|C0876081|MRV|MRV
Event|Event|SIMPLE_SEGMENT|2650,2653|false|false|false|||MRV
Event|Event|SIMPLE_SEGMENT|2660,2666|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|2670,2678|false|false|false|||thrombus
Finding|Pathologic Function|SIMPLE_SEGMENT|2670,2678|true|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|SIMPLE_SEGMENT|2682,2689|false|false|false|||venoous
Event|Event|SIMPLE_SEGMENT|2690,2700|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|2690,2700|false|false|false|C0040053|Thrombosis|thrombosis
Event|Event|SIMPLE_SEGMENT|2710,2721|false|false|false|||transferred
Event|Event|SIMPLE_SEGMENT|2741,2751|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|2741,2751|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|2741,2751|false|false|false|C0376636|Disease Management|management
Event|Activity|SIMPLE_SEGMENT|2760,2769|false|false|false|C0021822|Interview|interview
Event|Event|SIMPLE_SEGMENT|2760,2769|false|false|false|||interview
Finding|Intellectual Product|SIMPLE_SEGMENT|2760,2769|false|false|false|C0935630|Published Interview|interview
Event|Event|SIMPLE_SEGMENT|2781,2788|false|false|false|||provide
Finding|Finding|SIMPLE_SEGMENT|2789,2793|false|true|false|C4281574|Much|much
Event|Event|SIMPLE_SEGMENT|2794,2801|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2794,2801|false|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2794,2801|false|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2794,2801|false|true|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|2817,2820|false|false|false|||say
Event|Event|SIMPLE_SEGMENT|2846,2851|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|2846,2851|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|2858,2863|false|false|false|||keeps
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2868,2872|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2868,2872|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|2873,2879|false|false|false|||closed
Event|Event|SIMPLE_SEGMENT|2888,2899|false|false|false|||questioning
Finding|Mental Process|SIMPLE_SEGMENT|2888,2899|false|false|false|C0876928|Sexual Orientation - Questioning|questioning
Event|Event|SIMPLE_SEGMENT|2905,2912|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|2913,2921|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|2913,2921|false|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|2933,2941|false|false|false|||describe
Event|Event|SIMPLE_SEGMENT|2958,2966|false|false|false|||features
Event|Event|SIMPLE_SEGMENT|2979,2990|false|false|false|||photophobia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2979,2990|false|false|false|C0085636|Photophobia|photophobia
Event|Event|SIMPLE_SEGMENT|2999,3005|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|2999,3005|false|false|false|C1299582|Unable|unable
Event|Activity|SIMPLE_SEGMENT|3010,3021|false|false|false|C5909499|Participate|participate
Event|Event|SIMPLE_SEGMENT|3031,3042|false|false|false|||questioning
Finding|Mental Process|SIMPLE_SEGMENT|3031,3042|false|false|false|C0876928|Sexual Orientation - Questioning|questioning
Finding|Intellectual Product|SIMPLE_SEGMENT|3044,3049|false|false|false|C4050225|Often - answer to question|often
Event|Event|SIMPLE_SEGMENT|3058,3065|false|false|false|||tearful
Finding|Finding|SIMPLE_SEGMENT|3058,3065|false|false|false|C0424109|Weepiness|tearful
Event|Event|SIMPLE_SEGMENT|3070,3076|false|false|false|||saying
Event|Event|SIMPLE_SEGMENT|3082,3091|false|false|false|||questions
Event|Event|SIMPLE_SEGMENT|3096,3100|false|false|false|||hard
Event|Event|SIMPLE_SEGMENT|3113,3119|false|false|false|||father
Finding|Conceptual Entity|SIMPLE_SEGMENT|3113,3119|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|3113,3119|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Event|Event|SIMPLE_SEGMENT|3141,3148|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|3141,3148|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|3141,3151|true|false|false|C0262926|Medical History|history of
Event|Event|SIMPLE_SEGMENT|3152,3160|false|false|false|||seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|3152,3160|true|false|false|C0036572|Seizures|seizures
Anatomy|Body System|SIMPLE_SEGMENT|3165,3168|false|false|false|C3714787|Central Nervous System|CNS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3169,3178|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|3169,3178|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|3169,3178|false|false|false|C3714514|Infection|infection
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3195,3205|false|false|false|C0006107|Brain Concussion|concussion
Event|Event|SIMPLE_SEGMENT|3195,3205|false|false|false|||concussion
Event|Event|SIMPLE_SEGMENT|3219,3222|false|false|false|||old
Finding|Finding|SIMPLE_SEGMENT|3227,3247|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|3232,3239|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|3232,3239|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|3232,3239|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|3232,3239|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3232,3239|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|3232,3247|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3240,3247|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3240,3247|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3240,3247|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3249,3255|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|3249,3255|false|false|false|||Anemia
Finding|Functional Concept|SIMPLE_SEGMENT|3259,3265|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|3259,3273|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|3266,3273|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3266,3273|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3266,3273|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3266,3273|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|3279,3285|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|3279,3285|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|3279,3285|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|3279,3285|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|3279,3293|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|3286,3293|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|3286,3293|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|3286,3293|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|3286,3293|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|3295,3301|false|false|false|||Mother
Finding|Idea or Concept|SIMPLE_SEGMENT|3295,3301|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3309,3315|false|false|false|C0007570|Celiac Disease|celiac
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3309,3323|false|false|false|C0007570|Celiac Disease|celiac disease
Finding|Gene or Genome|SIMPLE_SEGMENT|3309,3323|false|false|false|C1332802|CTLA4 gene|celiac disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3316,3323|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|3316,3323|false|false|false|||disease
Finding|Functional Concept|SIMPLE_SEGMENT|3328,3338|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Finding|Pathologic Function|SIMPLE_SEGMENT|3328,3338|false|false|false|C0443146;C4551524|Autoimmune;Autoimmune reaction|autoimmune
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3328,3353|false|false|false|C0342158|Hypothyroidism, Autoimmune|autoimmune hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3339,3353|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Event|Event|SIMPLE_SEGMENT|3339,3353|false|false|false|||hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3355,3358|false|false|false|C1262020|Diffuse alveolar damage|Dad
Event|Event|SIMPLE_SEGMENT|3355,3358|false|false|false|||Dad
Finding|Intellectual Product|SIMPLE_SEGMENT|3355,3358|false|false|false|C3641946|Disability Assessment for Dementia Questionnaire|Dad
Event|Event|SIMPLE_SEGMENT|3362,3369|false|false|false|||healthy
Event|Event|SIMPLE_SEGMENT|3381,3387|false|false|false|||cousin
Event|Event|SIMPLE_SEGMENT|3393,3401|false|false|false|||seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|3393,3401|false|false|false|C0036572|Seizures|seizures
Event|Event|SIMPLE_SEGMENT|3405,3413|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|3405,3413|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|3405,3413|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|3405,3413|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|3405,3418|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3405,3418|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|3414,3418|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|3414,3418|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3414,3418|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3420,3429|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|3430,3434|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|3430,3434|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3430,3434|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|3462,3469|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|3462,3469|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|3462,3469|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|3485,3493|false|false|false|||sleeping
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3506,3509|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3506,3509|false|false|false|C0015392;C0700042;C4266572|Eye;Head>Eye;Orbital region|eye
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3506,3509|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3506,3509|false|false|false|C0015397;C0154094|Carcinoma in situ of eye;Disorder of eye|eye
Finding|Body Substance|SIMPLE_SEGMENT|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Finding|SIMPLE_SEGMENT|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Finding|Intellectual Product|SIMPLE_SEGMENT|3506,3509|false|false|false|C0262477;C1546630;C1550636|Eye - Specimen Source Code;Eye Specimen;Eye problem|eye
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3506,3513|false|false|false|C2706046|Eye lid|eye lid
Event|Event|SIMPLE_SEGMENT|3514,3524|false|false|false|||fluttering
Finding|Pathologic Function|SIMPLE_SEGMENT|3514,3524|false|false|false|C0016385|Cardiac Flutter|fluttering
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3526,3529|false|false|false|C0023759|Lip structure|lip
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3526,3529|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3526,3529|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|lip
Finding|Gene or Genome|SIMPLE_SEGMENT|3526,3529|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|lip
Event|Event|SIMPLE_SEGMENT|3530,3539|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|3530,3539|false|false|false|C0026649|Movement|movements
Finding|Sign or Symptom|SIMPLE_SEGMENT|3552,3566|false|false|false|C0233565|Bradykinesia|slow movements
Event|Event|SIMPLE_SEGMENT|3557,3566|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|3557,3566|false|false|false|C0026649|Movement|movements
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3570,3574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3570,3574|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3570,3574|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|3570,3574|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3570,3574|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3593,3598|false|false|false|C1512338|HEENT|HEENT
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3603,3609|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|3603,3609|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|3603,3609|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|3614,3622|false|false|false|||jaundice
Finding|Finding|SIMPLE_SEGMENT|3614,3622|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|SIMPLE_SEGMENT|3614,3622|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|SIMPLE_SEGMENT|3627,3634|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|3627,3634|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3638,3648|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|3654,3657|false|false|false|||RRR
Event|Event|SIMPLE_SEGMENT|3663,3667|false|false|false|||Pulm
Procedure|Health Care Activity|SIMPLE_SEGMENT|3663,3667|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Event|Event|SIMPLE_SEGMENT|3669,3678|false|false|false|||breathing
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3698,3701|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3698,3701|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3698,3701|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3703,3709|false|false|false|||clammy
Finding|Finding|SIMPLE_SEGMENT|3703,3709|false|false|false|C0392162|Clammy skin|clammy
Event|Event|SIMPLE_SEGMENT|3711,3715|false|false|false|||warm
Finding|Finding|SIMPLE_SEGMENT|3711,3715|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3711,3715|false|false|false|C0687712|warming process|warm
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3723,3727|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|3723,3727|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|3723,3727|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|3723,3727|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Mental Process|SIMPLE_SEGMENT|3743,3749|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3743,3756|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|3743,3756|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3750,3756|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|3750,3756|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|3750,3756|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|3778,3783|false|false|false|||upset
Finding|Mental Process|SIMPLE_SEGMENT|3778,3783|false|false|false|C3887804|Feeling upset|upset
Event|Event|SIMPLE_SEGMENT|3791,3795|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|3791,3795|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3791,3795|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|3803,3810|false|false|false|||tearful
Finding|Finding|SIMPLE_SEGMENT|3803,3810|false|false|false|C0424109|Weepiness|tearful
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3814,3819|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Intellectual Product|SIMPLE_SEGMENT|3821,3825|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|3826,3832|false|false|false|||abulic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3842,3847|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|3842,3847|false|false|false|||times
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3849,3853|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3849,3853|false|false|false|C5848506||Eyes
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3849,3858|false|false|false|C0266574|Ablepharon|Eyes open
Event|Event|SIMPLE_SEGMENT|3854,3858|false|false|false|||open
Event|Event|SIMPLE_SEGMENT|3875,3880|false|false|false|||voice
Finding|Idea or Concept|SIMPLE_SEGMENT|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|SIMPLE_SEGMENT|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|SIMPLE_SEGMENT|3875,3880|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Event|Event|SIMPLE_SEGMENT|3889,3897|false|false|false|||oriented
Event|Event|SIMPLE_SEGMENT|3913,3917|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|3924,3929|false|false|false|||Knows
Finding|Idea or Concept|SIMPLE_SEGMENT|3943,3951|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Intellectual Product|SIMPLE_SEGMENT|3965,3969|true|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Event|Event|SIMPLE_SEGMENT|3975,3979|false|false|false|||says
Finding|Idea or Concept|SIMPLE_SEGMENT|3995,4003|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|4018,4023|false|false|false|||tired
Finding|Finding|SIMPLE_SEGMENT|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|SIMPLE_SEGMENT|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|SIMPLE_SEGMENT|4018,4023|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Event|Event|SIMPLE_SEGMENT|4033,4039|false|false|false|||unable
Finding|Finding|SIMPLE_SEGMENT|4033,4039|false|false|false|C1299582|Unable|unable
Drug|Food|SIMPLE_SEGMENT|4044,4051|false|false|false|C0359589|Provide (product)|provide
Event|Activity|SIMPLE_SEGMENT|4044,4051|false|false|false|C1999230|Providing (action)|provide
Event|Event|SIMPLE_SEGMENT|4044,4051|false|false|false|||provide
Event|Event|SIMPLE_SEGMENT|4052,4059|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4052,4059|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|4061,4067|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|4061,4067|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4061,4067|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|4075,4085|false|false|false|||dysarthric
Event|Event|SIMPLE_SEGMENT|4087,4091|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|4096,4101|false|false|false|||words
Event|Event|SIMPLE_SEGMENT|4107,4112|false|false|false|||asked
Event|Event|SIMPLE_SEGMENT|4113,4122|false|false|false|||questions
Finding|Functional Concept|SIMPLE_SEGMENT|4127,4138|true|false|false|C0205359|Spontaneous|spontaneous
Event|Event|SIMPLE_SEGMENT|4139,4145|false|false|false|||speech
Finding|Organism Function|SIMPLE_SEGMENT|4139,4145|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4139,4145|false|false|false|C0846595|Speech assessment|speech
Event|Event|SIMPLE_SEGMENT|4146,4152|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|4146,4152|true|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|4146,4152|true|false|false|C3251815|Measurement of fluid output|output
Event|Event|SIMPLE_SEGMENT|4154,4161|false|false|false|||Follows
Finding|Gene or Genome|SIMPLE_SEGMENT|4162,4168|false|false|false|C1424587|LITAF gene|simple
Event|Event|SIMPLE_SEGMENT|4169,4177|false|false|false|||commands
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4188,4192|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4188,4192|false|false|false|C5848506||eyes
Event|Activity|SIMPLE_SEGMENT|4194,4198|false|false|false|C0206244|Lifting|lift
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4199,4203|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4199,4203|false|false|false|C5781420||legs
Event|Event|SIMPLE_SEGMENT|4212,4216|false|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|4212,4216|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|4220,4224|false|false|false|||name
Finding|Intellectual Product|SIMPLE_SEGMENT|4220,4224|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Event|Event|SIMPLE_SEGMENT|4226,4229|false|false|false|||key
Finding|Conceptual Entity|SIMPLE_SEGMENT|4226,4229|false|false|false|C1554080;C1706198|Key - HL7UpdateMode;Key - value|key
Finding|Intellectual Product|SIMPLE_SEGMENT|4226,4229|false|false|false|C1554080;C1706198|Key - HL7UpdateMode;Key - value|key
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4236,4243|false|false|false|C0015731;C1744713|Feathers|feather
Drug|Immunologic Factor|SIMPLE_SEGMENT|4236,4243|false|false|false|C3486460|Feathers (allergen)|feather
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4248,4254|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|4248,4254|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|4248,4254|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4255,4259|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4255,4259|false|false|false|C0018799|Heart Diseases|card
Event|Event|SIMPLE_SEGMENT|4255,4259|false|false|false|||card
Finding|Intellectual Product|SIMPLE_SEGMENT|4255,4259|false|false|false|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4255,4259|false|false|false|C5202809|CaRD Regimen|card
Finding|Intellectual Product|SIMPLE_SEGMENT|4264,4268|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|4269,4274|false|false|false|||stops
Event|Event|SIMPLE_SEGMENT|4275,4281|false|false|false|||naming
Event|Event|SIMPLE_SEGMENT|4286,4292|false|false|false|||closes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4297,4301|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4297,4301|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|4307,4312|false|false|false|||reads
Event|Event|SIMPLE_SEGMENT|4323,4331|false|false|false|||sentence
Finding|Intellectual Product|SIMPLE_SEGMENT|4323,4331|false|false|false|C0876929|Sentence|sentence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4335,4341|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|4335,4341|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|4335,4341|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4342,4346|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4342,4346|false|false|false|C0018799|Heart Diseases|card
Event|Event|SIMPLE_SEGMENT|4342,4346|false|false|false|||card
Finding|Intellectual Product|SIMPLE_SEGMENT|4342,4346|false|false|false|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4342,4346|false|false|false|C5202809|CaRD Regimen|card
Finding|Intellectual Product|SIMPLE_SEGMENT|4351,4355|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|4368,4374|false|false|false|||closes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4379,4383|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4379,4383|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|4390,4395|false|false|false|||asked
Event|Event|SIMPLE_SEGMENT|4399,4407|false|false|false|||describe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4408,4414|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|4408,4414|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|4408,4414|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4415,4419|false|false|false|C2340164|Stratum radiatum|card
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4415,4419|false|false|true|C0018799|Heart Diseases|card
Event|Event|SIMPLE_SEGMENT|4415,4419|false|false|false|||card
Finding|Intellectual Product|SIMPLE_SEGMENT|4415,4419|false|false|true|C3275277|Card (document)|card
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4415,4419|false|false|true|C5202809|CaRD Regimen|card
Event|Event|SIMPLE_SEGMENT|4432,4436|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|4461,4472|false|false|false|||participate
Event|Event|SIMPLE_SEGMENT|4484,4488|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|4484,4488|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4484,4488|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4492,4499|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4492,4506|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4492,4506|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4500,4506|false|false|false|C0027740|Nerve|Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4527,4533|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|4546,4550|false|false|false|||EOMI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4559,4568|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|SIMPLE_SEGMENT|4559,4568|false|false|false|||nystagmus
Event|Event|SIMPLE_SEGMENT|4578,4591|false|false|false|||confrontation
Finding|Finding|SIMPLE_SEGMENT|4578,4591|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4578,4591|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4578,4591|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4594,4610|false|false|false|C0029090|Ophthalmoscopy|Fundoscopic exam
Event|Event|SIMPLE_SEGMENT|4606,4610|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|4606,4610|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4606,4610|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|4611,4619|false|false|false|||revealed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4623,4634|true|false|false|C0030353|Papilledema|papilledema
Event|Event|SIMPLE_SEGMENT|4623,4634|false|false|false|||papilledema
Event|Event|SIMPLE_SEGMENT|4636,4644|false|false|false|||exudates
Finding|Body Substance|SIMPLE_SEGMENT|4636,4644|false|false|false|C0015388|Exudate|exudates
Event|Event|SIMPLE_SEGMENT|4649,4660|false|false|false|||hemorrhages
Finding|Pathologic Function|SIMPLE_SEGMENT|4649,4660|false|false|false|C0019080|Hemorrhage|hemorrhages
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4663,4666|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|4663,4666|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4671,4677|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4671,4683|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|SIMPLE_SEGMENT|4671,4683|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|SIMPLE_SEGMENT|4678,4683|false|false|false|||droop
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4685,4691|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4692,4703|false|false|false|C1995013|Set of muscles|musculature
Event|Event|SIMPLE_SEGMENT|4704,4713|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|4704,4713|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|4704,4713|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|4720,4727|false|false|false|||grimace
Finding|Sign or Symptom|SIMPLE_SEGMENT|4720,4727|false|false|false|C0239779|Grimaces|grimace
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4730,4734|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|SIMPLE_SEGMENT|4730,4734|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|SIMPLE_SEGMENT|4730,4734|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|SIMPLE_SEGMENT|4736,4743|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|SIMPLE_SEGMENT|4736,4743|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|SIMPLE_SEGMENT|4744,4750|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|4744,4750|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|4754,4758|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|4754,4758|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|4754,4758|false|false|false|C0582103|Medical Examination|exam
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4767,4773|false|false|false|C0700374|Palate|Palate
Event|Event|SIMPLE_SEGMENT|4774,4782|false|false|false|||elevates
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4804,4810|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4804,4810|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Event|Event|SIMPLE_SEGMENT|4804,4810|false|false|false|||Tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|4804,4810|false|false|false|C0872394|Procedure on tongue|Tongue
Event|Event|SIMPLE_SEGMENT|4811,4820|false|false|false|||protrudes
Anatomy|Cell Component|SIMPLE_SEGMENT|4824,4831|false|false|false|C1660780|midline cell component|midline
Finding|Functional Concept|SIMPLE_SEGMENT|4835,4840|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4849,4853|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|4849,4853|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|SIMPLE_SEGMENT|4849,4853|false|false|false|||bulk
Event|Event|SIMPLE_SEGMENT|4855,4859|false|false|false|||tone
Event|Event|SIMPLE_SEGMENT|4876,4880|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|4892,4896|false|false|false|||move
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4901,4905|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4901,4905|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4901,4905|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|SIMPLE_SEGMENT|4901,4905|false|false|false|||arms
Finding|Gene or Genome|SIMPLE_SEGMENT|4901,4905|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|4901,4905|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4912,4916|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4912,4916|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4912,4916|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|SIMPLE_SEGMENT|4912,4916|false|false|false|||arms
Finding|Gene or Genome|SIMPLE_SEGMENT|4912,4916|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|4912,4916|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|SIMPLE_SEGMENT|4917,4923|false|false|false|||placed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4933,4937|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4933,4937|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4933,4937|false|false|false|C0362076|Problems with head|head
Event|Event|SIMPLE_SEGMENT|4933,4937|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4933,4937|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4943,4947|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4943,4947|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4943,4947|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|SIMPLE_SEGMENT|4943,4947|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|4943,4947|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4964,4968|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4964,4968|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|SIMPLE_SEGMENT|4964,4968|false|false|false|||face
Finding|Gene or Genome|SIMPLE_SEGMENT|4964,4968|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4980,4985|false|false|false|C0991568|Drops - Drug Form|drops
Event|Event|SIMPLE_SEGMENT|4980,4985|false|false|false|||drops
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4993,4996|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|4993,4996|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|4993,4996|false|false|false|C2346952|Bachelor of Education|bed
Finding|Finding|SIMPLE_SEGMENT|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Functional Concept|SIMPLE_SEGMENT|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Finding|Idea or Concept|SIMPLE_SEGMENT|5002,5012|false|false|false|C2587213;C2911690;C4761797|Control function;Controlled mark;Disease Controlled|controlled
Event|Event|SIMPLE_SEGMENT|5013,5020|false|false|false|||fashion
Event|Event|SIMPLE_SEGMENT|5032,5036|false|false|false|||lift
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5041,5045|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5041,5045|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5041,5045|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|SIMPLE_SEGMENT|5041,5045|false|false|false|||arms
Finding|Gene or Genome|SIMPLE_SEGMENT|5041,5045|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|5041,5045|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|SIMPLE_SEGMENT|5049,5053|false|false|false|||hold
Event|Event|SIMPLE_SEGMENT|5063,5068|false|false|false|||rails
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5076,5079|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|5076,5079|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|5076,5079|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|5099,5104|false|false|false|||lifts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5109,5113|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5109,5113|false|false|false|C5781420||legs
Event|Event|SIMPLE_SEGMENT|5114,5125|false|false|false|||antigravity
Event|Event|SIMPLE_SEGMENT|5176,5187|false|false|false|||withdrawals
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5191,5208|false|false|false|C1140618|Upper Extremity|upper extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5197,5208|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|5234,5245|false|false|false|||withdrawals
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5249,5254|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|5249,5254|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5249,5266|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5255,5266|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|5278,5285|false|false|false|||stimuli
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|5278,5285|false|false|false|C0234402|Stimulus|stimuli
Event|Event|SIMPLE_SEGMENT|5290,5294|false|false|false|||says
Event|Event|SIMPLE_SEGMENT|5304,5308|false|false|false|||DTRs
Finding|Gene or Genome|SIMPLE_SEGMENT|5317,5320|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|SIMPLE_SEGMENT|5317,5320|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5325,5328|false|false|false|C0030587|Paroxysmal atrial tachycardia|Pat
Drug|Organic Chemical|SIMPLE_SEGMENT|5325,5328|false|false|false|C2825250|Fenamole|Pat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5325,5328|false|false|false|C2825250|Fenamole|Pat
Event|Event|SIMPLE_SEGMENT|5325,5328|false|false|false|||Pat
Finding|Molecular Function|SIMPLE_SEGMENT|5325,5328|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|Pat
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5325,5328|false|false|false|C3897364|Thermoacoustic Computed Tomography|Pat
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5329,5332|false|false|false|C0001080|Achondroplasia|Ach
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Drug|Organic Chemical|SIMPLE_SEGMENT|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5329,5332|false|false|false|C0001041|acetylcholine|Ach
Event|Event|SIMPLE_SEGMENT|5329,5332|false|false|false|||Ach
Finding|Gene or Genome|SIMPLE_SEGMENT|5329,5332|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Finding|Sign or Symptom|SIMPLE_SEGMENT|5329,5332|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5380,5387|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|Plantar
Event|Event|SIMPLE_SEGMENT|5388,5396|false|false|false|||response
Finding|Finding|SIMPLE_SEGMENT|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|SIMPLE_SEGMENT|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|SIMPLE_SEGMENT|5388,5396|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5401,5407|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Event|Event|SIMPLE_SEGMENT|5423,5435|false|false|false|||Coordination
Finding|Functional Concept|SIMPLE_SEGMENT|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|5423,5435|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Body Substance|SIMPLE_SEGMENT|5437,5444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5437,5444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5437,5444|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5455,5466|false|false|false|||participate
Finding|Finding|SIMPLE_SEGMENT|5469,5473|false|false|false|C0016928|Gait|Gait
Event|Event|SIMPLE_SEGMENT|5485,5491|false|false|false|||assess
Finding|Body Substance|SIMPLE_SEGMENT|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5495,5502|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|5513,5516|false|false|false|||get
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5524,5527|false|true|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|5524,5527|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|5524,5527|false|true|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|5529,5538|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5529,5538|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5529,5538|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5529,5538|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5529,5538|false|false|false|C0030685|Patient Discharge|Discharge
Event|Event|SIMPLE_SEGMENT|5539,5543|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|5539,5543|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5539,5543|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|5545,5552|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|5545,5552|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|5545,5552|false|false|false|C3812897|General medical service|General
Event|Event|SIMPLE_SEGMENT|5554,5561|false|false|false|||sitting
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5583,5587|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5583,5587|false|false|false|C5848506||eyes
Event|Event|SIMPLE_SEGMENT|5588,5594|false|false|false|||closed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5595,5600|false|false|false|C1512338|HEENT|HEENT
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5605,5611|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|5605,5611|false|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|5605,5611|true|false|false|C0548346|Trauma assessment and care|trauma
Event|Event|SIMPLE_SEGMENT|5616,5624|false|false|false|||jaundice
Finding|Finding|SIMPLE_SEGMENT|5616,5624|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Finding|Sign or Symptom|SIMPLE_SEGMENT|5616,5624|true|false|false|C0022346;C2010848;C2203646|Icterus;jaundice;yellow skin or eyes (symptom)|jaundice
Event|Event|SIMPLE_SEGMENT|5629,5636|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|5629,5636|true|false|false|C0221198|Lesion|lesions
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5640,5650|false|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5656,5661|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5656,5661|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|5656,5661|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5656,5661|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|SIMPLE_SEGMENT|5656,5673|false|false|false|C0085610;C2108107;C5235162|Sinus Bradycardia by ECG Finding;Sinus bradycardia;continuous electrocardiogram sinus bradycardia|sinus bradycardia
Finding|Pathologic Function|SIMPLE_SEGMENT|5656,5673|false|false|false|C0085610;C2108107;C5235162|Sinus Bradycardia by ECG Finding;Sinus bradycardia;continuous electrocardiogram sinus bradycardia|sinus bradycardia
Event|Event|SIMPLE_SEGMENT|5662,5673|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|5662,5673|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|SIMPLE_SEGMENT|5684,5688|false|false|false|||Pulm
Procedure|Health Care Activity|SIMPLE_SEGMENT|5684,5688|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5719,5722|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|5719,5722|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|5719,5722|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|5724,5728|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|5724,5728|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5724,5728|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|5733,5737|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5738,5746|false|false|false|||perfused
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5751,5755|true|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|5751,5755|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|5751,5755|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|5751,5755|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Event|Event|SIMPLE_SEGMENT|5759,5767|false|false|false|||mottling
Finding|Finding|SIMPLE_SEGMENT|5759,5767|false|false|false|C0302133|Mottling|mottling
Finding|Mental Process|SIMPLE_SEGMENT|5783,5789|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5783,5796|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|5783,5796|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5790,5796|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|5790,5796|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|5790,5796|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|5808,5817|false|false|false|||questions
Event|Event|SIMPLE_SEGMENT|5834,5842|false|false|false|||sentence
Finding|Intellectual Product|SIMPLE_SEGMENT|5834,5842|false|false|false|C0876929|Sentence|sentence
Event|Event|SIMPLE_SEGMENT|5849,5854|false|false|false|||humor
Finding|Intellectual Product|SIMPLE_SEGMENT|5849,5854|false|false|false|C0020168|Humor|humor
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5849,5854|false|false|false|C0597811|Humor therapy|humor
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|5859,5866|false|false|false|C1704241|complex (molecular entity)|complex
Event|Event|SIMPLE_SEGMENT|5867,5876|false|false|false|||sentences
Finding|Intellectual Product|SIMPLE_SEGMENT|5867,5876|false|false|false|C0876929|Sentence|sentences
Event|Event|SIMPLE_SEGMENT|5877,5885|false|false|false|||observed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5893,5897|false|false|false|C0015392|Eye|Eyes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5893,5897|false|false|false|C5848506||Eyes
Event|Event|SIMPLE_SEGMENT|5913,5918|false|false|false|||close
Finding|Finding|SIMPLE_SEGMENT|5913,5918|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|SIMPLE_SEGMENT|5913,5918|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|SIMPLE_SEGMENT|5932,5939|false|false|false|||talking
Event|Event|SIMPLE_SEGMENT|5941,5947|false|false|false|||Speech
Finding|Organism Function|SIMPLE_SEGMENT|5941,5947|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5941,5947|false|false|false|C0846595|Speech assessment|Speech
Event|Event|SIMPLE_SEGMENT|5955,5965|false|false|false|||dysarthric
Finding|Functional Concept|SIMPLE_SEGMENT|5970,5981|true|false|false|C0205359|Spontaneous|spontaneous
Event|Event|SIMPLE_SEGMENT|5982,5988|false|false|false|||speech
Finding|Organism Function|SIMPLE_SEGMENT|5982,5988|true|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5982,5988|true|false|false|C0846595|Speech assessment|speech
Event|Event|SIMPLE_SEGMENT|5989,5995|false|false|false|||output
Finding|Conceptual Entity|SIMPLE_SEGMENT|5989,5995|true|false|false|C1709366|system output|output
Procedure|Health Care Activity|SIMPLE_SEGMENT|5989,5995|true|false|false|C3251815|Measurement of fluid output|output
Finding|Gene or Genome|SIMPLE_SEGMENT|6005,6011|false|false|false|C1424587|LITAF gene|simple
Event|Event|SIMPLE_SEGMENT|6012,6020|false|false|false|||commands
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6024,6031|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6024,6038|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6024,6038|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6032,6038|false|false|false|C0027740|Nerve|Nerves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6057,6063|false|false|false|C0034121|Pupil|Pupils
Event|Event|SIMPLE_SEGMENT|6076,6080|false|false|false|||EOMI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6089,6098|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|SIMPLE_SEGMENT|6089,6098|false|false|false|||nystagmus
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6104,6110|false|false|false|C0015450|Face|facial
Finding|Finding|SIMPLE_SEGMENT|6104,6120|false|false|false|C0517999|facial sensation|facial sensation
Event|Event|SIMPLE_SEGMENT|6111,6120|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|6111,6120|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6111,6120|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6111,6120|false|false|false|C2229507|sensory exam|sensation
Finding|Finding|SIMPLE_SEGMENT|6121,6127|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6139,6142|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|SIMPLE_SEGMENT|6139,6142|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6147,6153|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6147,6159|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|SIMPLE_SEGMENT|6147,6159|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|SIMPLE_SEGMENT|6154,6159|false|false|false|||droop
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6161,6167|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6168,6179|false|false|false|C1995013|Set of muscles|musculature
Event|Event|SIMPLE_SEGMENT|6180,6189|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|6180,6189|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|6180,6189|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Event|Event|SIMPLE_SEGMENT|6195,6202|false|false|false|||grimace
Finding|Sign or Symptom|SIMPLE_SEGMENT|6195,6202|false|false|false|C0239779|Grimaces|grimace
Finding|Functional Concept|SIMPLE_SEGMENT|6207,6214|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|SIMPLE_SEGMENT|6207,6214|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6215,6221|false|false|false|C0015450|Face|facial
Event|Event|SIMPLE_SEGMENT|6222,6231|false|false|false|||movements
Finding|Organism Function|SIMPLE_SEGMENT|6222,6231|false|false|false|C0026649|Movement|movements
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6245,6251|false|false|false|C0700374|Palate|palate
Event|Event|SIMPLE_SEGMENT|6252,6260|false|false|false|||elevates
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6276,6282|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6276,6282|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Procedure|Health Care Activity|SIMPLE_SEGMENT|6276,6282|false|false|false|C0872394|Procedure on tongue|tongue
Finding|Finding|SIMPLE_SEGMENT|6276,6290|false|false|false|C3693372|tongue midline|tongue midline
Anatomy|Cell Component|SIMPLE_SEGMENT|6283,6290|false|false|false|C1660780|midline cell component|midline
Finding|Functional Concept|SIMPLE_SEGMENT|6293,6298|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6307,6311|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|SIMPLE_SEGMENT|6307,6311|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|SIMPLE_SEGMENT|6307,6311|false|false|false|||bulk
Event|Event|SIMPLE_SEGMENT|6313,6317|false|false|false|||tone
Event|Activity|SIMPLE_SEGMENT|6330,6337|false|false|false|C0206244|Lifting|Lifting
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6338,6342|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6338,6342|false|false|false|C5782111||arms
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6338,6342|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|SIMPLE_SEGMENT|6338,6342|false|false|false|||arms
Finding|Gene or Genome|SIMPLE_SEGMENT|6338,6342|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|SIMPLE_SEGMENT|6338,6342|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6338,6351|false|false|false|C0015385|Limb structure|arms and legs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6347,6351|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6347,6351|false|false|false|C5781420||legs
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6360,6367|true|false|false|C0282189|Gravity (physical force)|gravity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6384,6394|true|false|false|C1442099|Resistance|resistance
Event|Event|SIMPLE_SEGMENT|6384,6394|false|false|false|||resistance
Finding|Mental Process|SIMPLE_SEGMENT|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Physiologic Function|SIMPLE_SEGMENT|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Finding|Social Behavior|SIMPLE_SEGMENT|6384,6394|true|false|false|C0237834;C0683598;C1514892|Resistance (Psychotherapeutic);Resistance Process;social resistance|resistance
Event|Event|SIMPLE_SEGMENT|6412,6421|false|false|false|||Sensation
Finding|Finding|SIMPLE_SEGMENT|6412,6421|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6412,6421|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|6412,6421|false|false|false|C2229507|sensory exam|Sensation
Event|Event|SIMPLE_SEGMENT|6422,6428|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|6422,6428|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|6432,6437|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|6432,6437|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|6432,6437|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6432,6437|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|6442,6453|false|false|false|||temperature
Procedure|Health Care Activity|SIMPLE_SEGMENT|6442,6453|false|false|false|C0886414|Body temperature measurement|temperature
Event|Event|SIMPLE_SEGMENT|6467,6471|false|false|false|||DTRs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6476,6484|false|false|false|C0030647|Patella|patellar
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6486,6492|false|false|false|C0559499|Biceps brachii muscle structure|biceps
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6494,6509|false|false|false|C0224264|Structure of brachioradialis muscle|brachioradialis
Event|Event|SIMPLE_SEGMENT|6523,6535|false|false|false|||Coordination
Finding|Functional Concept|SIMPLE_SEGMENT|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|SIMPLE_SEGMENT|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|SIMPLE_SEGMENT|6523,6535|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|SIMPLE_SEGMENT|6540,6549|false|false|false|||dysmetria
Finding|Finding|SIMPLE_SEGMENT|6540,6549|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Event|Event|SIMPLE_SEGMENT|6553,6559|false|false|false|||tremor
Finding|Sign or Symptom|SIMPLE_SEGMENT|6553,6559|true|false|false|C0040822|Tremor|tremor
Finding|Finding|SIMPLE_SEGMENT|6564,6568|false|false|false|C0016928|Gait|Gait
Finding|Finding|SIMPLE_SEGMENT|6580,6584|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|SIMPLE_SEGMENT|6618,6627|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6628,6632|false|false|false|C0587081|Laboratory test finding|labs
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6664,6671|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|6664,6671|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6664,6671|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6664,6671|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6675,6679|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|6675,6679|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6675,6679|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|6675,6679|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6675,6679|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6694,6700|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|6694,6700|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|6694,6700|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6694,6700|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6706,6715|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|6706,6715|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|6706,6715|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6706,6715|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6720,6728|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|6720,6728|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|6720,6728|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6720,6728|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6739,6742|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6739,6742|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|6739,6742|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|6739,6742|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|6739,6742|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6746,6751|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6746,6755|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6746,6755|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6746,6755|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6752,6755|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6752,6755|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|6752,6755|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|6752,6755|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6773,6776|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6773,6776|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|6773,6776|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|6773,6776|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|6773,6776|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6773,6776|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6777,6781|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|6777,6781|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|6777,6781|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|6777,6781|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6777,6781|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6785,6788|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6785,6788|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|6785,6788|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|6785,6788|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|6785,6788|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6789,6793|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|6789,6793|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|6789,6793|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|6789,6793|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6789,6793|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6798,6801|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|6798,6801|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|6798,6801|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|6798,6801|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|6798,6801|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6798,6806|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|6798,6806|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6798,6806|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|6802,6806|false|false|false|||PHOS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|6838,6845|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|6838,6845|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|6838,6845|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6838,6845|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6850,6859|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Event|Event|SIMPLE_SEGMENT|6850,6859|false|false|false|||PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6850,6859|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6864,6873|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6864,6873|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Drug|Enzyme|SIMPLE_SEGMENT|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6892,6895|false|false|false|C5565118|TGM2 protein, human|tTG
Event|Event|SIMPLE_SEGMENT|6892,6895|false|false|false|||tTG
Finding|Gene or Genome|SIMPLE_SEGMENT|6892,6895|false|false|false|C5575307|TGM2 wt Allele|tTG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Immunologic Factor|SIMPLE_SEGMENT|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6896,6899|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Event|Event|SIMPLE_SEGMENT|6896,6899|false|false|false|||IgA
Finding|Gene or Genome|SIMPLE_SEGMENT|6896,6899|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|IgA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6896,6899|false|false|false|C0202083|Immunoglobulin A measurement|IgA
Anatomy|Cell|SIMPLE_SEGMENT|6916,6919|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|6924,6927|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6924,6927|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6924,6927|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6934,6937|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6934,6937|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|6934,6937|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|6934,6937|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6934,6937|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|6943,6946|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6943,6946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6943,6946|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|6952,6955|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|6952,6955|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|6952,6955|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6952,6955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6952,6955|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|6960,6963|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6960,6963|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|6960,6963|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|6960,6963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|6960,6963|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6960,6963|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|6969,6973|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6969,6973|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|7013,7016|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7013,7016|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Body Substance|SIMPLE_SEGMENT|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7039,7044|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|SIMPLE_SEGMENT|7052,7058|false|false|false|||RANDOM
Finding|Body Substance|SIMPLE_SEGMENT|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7071,7076|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Classification|SIMPLE_SEGMENT|7082,7090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|7082,7090|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7082,7090|false|false|false|C5237010|Expression Negative|NEGATIVE
Finding|Body Substance|SIMPLE_SEGMENT|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7103,7108|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Event|Event|SIMPLE_SEGMENT|7119,7122|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7119,7122|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|7132,7135|false|false|false|C5848551|Neg - answer|NEG
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Organic Chemical|SIMPLE_SEGMENT|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7136,7143|false|false|false|C0221793;C0376196|Opiate Alkaloids;Opiates|opiates
Event|Event|SIMPLE_SEGMENT|7136,7143|false|false|false|||opiates
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7136,7143|false|false|false|C0242401|Opiate Measurement|opiates
Event|Event|SIMPLE_SEGMENT|7144,7147|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7144,7147|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7149,7156|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|SIMPLE_SEGMENT|7149,7156|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7149,7156|false|false|false|C0009170|cocaine|cocaine
Event|Event|SIMPLE_SEGMENT|7149,7156|false|false|false|||cocaine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7149,7156|false|false|false|C0202362|Cocaine measurement|cocaine
Event|Event|SIMPLE_SEGMENT|7157,7160|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7157,7160|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|7170,7173|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|SIMPLE_SEGMENT|7182,7185|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|7194,7197|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7194,7197|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7210,7215|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|7210,7222|false|false|false|C0278030|Color of urine|URINE  COLOR
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7217,7222|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7217,7222|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|COLOR
Event|Event|SIMPLE_SEGMENT|7217,7222|false|false|false|||COLOR
Drug|Organic Chemical|SIMPLE_SEGMENT|7223,7228|false|false|false|C4047917|Cereal plant straw|Straw
Event|Event|SIMPLE_SEGMENT|7236,7241|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|7236,7241|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|SIMPLE_SEGMENT|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7261,7266|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7261,7273|false|false|false|C0018965|Hematuria|URINE  BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7268,7273|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|7268,7273|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|7268,7273|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|SIMPLE_SEGMENT|7274,7276|false|false|false|||LG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7278,7285|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|NITRITE
Event|Event|SIMPLE_SEGMENT|7286,7289|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7286,7289|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7290,7297|false|false|false|C0033684|Proteins|PROTEIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7290,7297|false|false|false|C0033684|Proteins|PROTEIN
Event|Event|SIMPLE_SEGMENT|7290,7297|false|false|false|||PROTEIN
Finding|Conceptual Entity|SIMPLE_SEGMENT|7290,7297|false|false|false|C1521746|Protein Info|PROTEIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7290,7297|false|false|false|C0202202|Protein measurement|PROTEIN
Event|Event|SIMPLE_SEGMENT|7298,7301|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7298,7301|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7303,7310|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|7303,7310|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7303,7310|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7303,7310|false|false|false|C0337438|Glucose measurement|GLUCOSE
Event|Event|SIMPLE_SEGMENT|7311,7314|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7311,7314|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|SIMPLE_SEGMENT|7315,7321|false|false|false|C0022634|Ketones|KETONE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Organic Chemical|SIMPLE_SEGMENT|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7326,7335|false|false|false|C0005437;C5241078|Bilirubin;bilirubin preparation|BILIRUBIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7326,7335|false|false|false|C0201913;C0863174|Bilirubin, total measurement;blood bilirubin level test|BILIRUBIN
Event|Event|SIMPLE_SEGMENT|7336,7339|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7336,7339|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|7350,7353|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7350,7353|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|7367,7370|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|7367,7370|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|SIMPLE_SEGMENT|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7383,7388|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7383,7393|false|false|false|C0221752;C2188659|Red blood cells urine positive|URINE  RBC
Anatomy|Cell|SIMPLE_SEGMENT|7390,7393|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7390,7393|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7390,7393|false|false|false|C0014792|Erythrocytes|RBC
Anatomy|Cell|SIMPLE_SEGMENT|7397,7400|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|SIMPLE_SEGMENT|7403,7411|false|false|false|C1510439|bacteria aspects|BACTERIA
Event|Event|SIMPLE_SEGMENT|7412,7415|false|false|false|||FEW
Drug|Food|SIMPLE_SEGMENT|7417,7422|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Immunologic Factor|SIMPLE_SEGMENT|7417,7422|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|7417,7422|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7417,7422|false|false|false|C0043392;C0717551|Candida albicans allergenic extract;Yeast, Dried|YEAST
Event|Event|SIMPLE_SEGMENT|7423,7427|false|false|false|||NONE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7429,7432|false|false|false|C0267963|Exocrine pancreatic insufficiency|EPI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7429,7432|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7429,7432|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Hormone|SIMPLE_SEGMENT|7429,7432|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Organic Chemical|SIMPLE_SEGMENT|7429,7432|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7429,7432|false|false|false|C0014563;C4281721|Tissue Factor Pathway Inhibitor, human;epinephrine|EPI
Event|Event|SIMPLE_SEGMENT|7429,7432|false|false|false|||EPI
Finding|Gene or Genome|SIMPLE_SEGMENT|7429,7432|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Finding|Intellectual Product|SIMPLE_SEGMENT|7429,7432|false|false|false|C0451152;C1420705;C3273314|Eysenck personality inventory;TFPI gene;TFPI wt Allele|EPI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7429,7432|false|false|false|C0162734;C3641909|Echo-Planar Imaging;Electronic Portal Imaging|EPI
Finding|Body Substance|SIMPLE_SEGMENT|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|7447,7452|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|SIMPLE_SEGMENT|7447,7460|false|false|false|C0455910|Mucus in urine (finding)|URINE  MUCOUS
Finding|Body Substance|SIMPLE_SEGMENT|7454,7460|false|false|false|C0026727;C2753459|Mucus (substance);mucus layer|MUCOUS
Event|Event|SIMPLE_SEGMENT|7461,7465|false|false|false|||RARE
Finding|Gene or Genome|SIMPLE_SEGMENT|7461,7465|false|false|false|C1514917|Retinoic Acid Response Element|RARE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7485,7488|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|7485,7488|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7485,7488|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Anatomy|Cell|SIMPLE_SEGMENT|7512,7515|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|7512,7515|false|false|false|||WBC
Anatomy|Cell|SIMPLE_SEGMENT|7520,7523|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7520,7523|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7520,7523|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7529,7532|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7529,7532|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|7529,7532|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|7529,7532|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7529,7532|false|false|false|C0019029|Hemoglobin concentration|HGB
Event|Event|SIMPLE_SEGMENT|7538,7541|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7538,7541|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7538,7541|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|7547,7550|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|7547,7550|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7547,7550|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7547,7550|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7547,7550|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|7555,7558|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7555,7558|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|7555,7558|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|7555,7558|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|7555,7558|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7555,7558|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|7564,7568|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7564,7568|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|SIMPLE_SEGMENT|7608,7613|false|false|false|||NEUTS
Drug|Antibiotic|SIMPLE_SEGMENT|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|7623,7628|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7633,7636|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|7633,7636|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|7633,7636|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|SIMPLE_SEGMENT|7740,7743|false|false|false|||PLT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7740,7743|false|false|false|C0201617|Primed lymphocyte test|PLT
Finding|Classification|SIMPLE_SEGMENT|7772,7775|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|PO2
Finding|Molecular Function|SIMPLE_SEGMENT|7772,7775|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|PO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7772,7775|false|false|false|C1283004|PO2 measurement|PO2
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7780,7784|false|false|false|C0391839|Carbon dioxide, partial pressure|PCO2
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7780,7784|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|PCO2
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7804,7807|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7804,7807|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|SIMPLE_SEGMENT|7804,7807|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|7804,7807|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7811,7815|false|false|false|C2987514|Anatomical base|BASE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Chemical Viewed Functionally|SIMPLE_SEGMENT|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7811,7815|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|BASE
Finding|Gene or Genome|SIMPLE_SEGMENT|7811,7815|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Finding|Idea or Concept|SIMPLE_SEGMENT|7811,7815|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|BASE
Event|Event|SIMPLE_SEGMENT|7821,7829|false|false|false|||COMMENTS
Finding|Intellectual Product|SIMPLE_SEGMENT|7821,7829|false|false|false|C0282411;C0947611|Comment;Published Comment|COMMENTS
Event|Event|SIMPLE_SEGMENT|7836,7839|false|false|false|||TOP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7854,7861|false|false|false|C0017725|glucose|GLUCOSE
Event|Event|SIMPLE_SEGMENT|7854,7861|false|false|false|||GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7854,7861|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7854,7861|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7865,7869|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|7865,7869|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7865,7869|false|false|false|C0041942|urea|UREA
Event|Event|SIMPLE_SEGMENT|7865,7869|false|false|false|||UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7865,7869|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7884,7890|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Event|Event|SIMPLE_SEGMENT|7884,7890|false|false|false|||SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|7884,7890|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7884,7890|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7896,7905|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Event|Event|SIMPLE_SEGMENT|7896,7905|false|false|false|||POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|7896,7905|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7896,7905|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7910,7918|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Event|Event|SIMPLE_SEGMENT|7910,7918|false|false|false|||CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|7910,7918|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7910,7918|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7929,7932|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7929,7932|false|false|false|C0007012|carbon dioxide|CO2
Event|Event|SIMPLE_SEGMENT|7929,7932|false|false|false|||CO2
Finding|Finding|SIMPLE_SEGMENT|7929,7932|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|7929,7932|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7936,7941|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7936,7945|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7936,7945|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7936,7945|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7942,7945|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7942,7945|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Event|Event|SIMPLE_SEGMENT|7942,7945|false|false|false|||GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|7942,7945|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7995,7998|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7995,7998|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|7995,7998|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|7995,7998|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|7995,7998|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7995,7998|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7999,8003|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|7999,8003|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|7999,8003|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|7999,8003|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7999,8003|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8007,8010|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8007,8010|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|8007,8010|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|8007,8010|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|8007,8010|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8011,8015|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|8011,8015|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|8011,8015|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|8011,8015|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8011,8015|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8023,8026|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|SIMPLE_SEGMENT|8023,8026|false|false|false|C0010287|Creatine Kinase|CPK
Event|Event|SIMPLE_SEGMENT|8023,8026|false|false|false|||CPK
Finding|Gene or Genome|SIMPLE_SEGMENT|8023,8026|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8023,8026|false|false|false|C0201973|Creatine kinase measurement|CPK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8031,8034|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|8031,8034|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|8031,8034|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|8031,8034|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|8031,8034|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8071,8076|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|SIMPLE_SEGMENT|8071,8076|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|SIMPLE_SEGMENT|8071,8076|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8071,8076|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8094,8101|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|SIMPLE_SEGMENT|8094,8101|false|false|false|||ALBUMIN
Finding|Gene or Genome|SIMPLE_SEGMENT|8094,8101|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|SIMPLE_SEGMENT|8094,8101|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8094,8101|false|false|false|C0201838|Albumin measurement|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Drug|Vitamin|SIMPLE_SEGMENT|8106,8113|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|CALCIUM
Event|Event|SIMPLE_SEGMENT|8106,8113|false|false|false|||CALCIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|8106,8113|false|false|false|C4553026|Calcium metabolic function|CALCIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8106,8113|false|false|false|C0201925|Calcium measurement|CALCIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8118,8127|false|false|false|C0031603;C1601799|Phosphates;phosphate ion|PHOSPHATE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8118,8127|false|false|false|C0523826|Phosphate measurement|PHOSPHATE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8133,8142|false|false|false|C0024467;C3540792;C3714621|Magnesium Drug Class;Magnesium supplements, alimentary tract and metabolism;magnesium|MAGNESIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8133,8142|false|false|false|C0373675|Magnesium measurement|MAGNESIUM
Event|Event|SIMPLE_SEGMENT|8161,8164|false|false|false|||VIT
Finding|Gene or Genome|SIMPLE_SEGMENT|8161,8164|false|false|false|C1421454;C5401427;C5401428|AML Vitals Table;EWS Vitals Table;VIT gene|VIT
Finding|Intellectual Product|SIMPLE_SEGMENT|8161,8164|false|false|false|C1421454;C5401427;C5401428|AML Vitals Table;EWS Vitals Table;VIT gene|VIT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8161,8164|false|false|false|C1831721|VIT Regimen|VIT
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Organic Chemical|SIMPLE_SEGMENT|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Drug|Vitamin|SIMPLE_SEGMENT|8161,8168|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|VIT B12
Event|Event|SIMPLE_SEGMENT|8165,8168|false|false|false|||B12
Finding|Gene or Genome|SIMPLE_SEGMENT|8165,8168|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8188,8191|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8188,8191|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|8188,8191|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8188,8191|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8210,8213|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|SIMPLE_SEGMENT|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8210,8213|false|false|false|C0040160|thyrotropin|TSH
Event|Event|SIMPLE_SEGMENT|8210,8213|false|false|false|||TSH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8210,8213|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8250,8253|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Drug|Immunologic Factor|SIMPLE_SEGMENT|8250,8253|false|false|false|C0006560;C4048285|C-Reactive Protein, human;C-reactive protein|CRP
Event|Event|SIMPLE_SEGMENT|8250,8253|false|false|false|||CRP
Finding|Gene or Genome|SIMPLE_SEGMENT|8250,8253|false|false|false|C1413716;C1413766;C1826658;C1879974|CRP gene;CRP wt Allele;CSRP1 gene;PPIAP10 gene|CRP
Event|Event|SIMPLE_SEGMENT|8259,8264|false|false|false|||dsDNA
Event|Event|SIMPLE_SEGMENT|8265,8273|false|false|false|||NEGATIVE
Finding|Classification|SIMPLE_SEGMENT|8265,8273|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|8265,8273|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8265,8273|false|false|false|C5237010|Expression Negative|NEGATIVE
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8315,8318|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|8315,8318|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|8315,8318|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|8319,8322|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|8319,8322|false|false|false|C5848551|Neg - answer|NEG
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8323,8330|false|false|false|C0161679|Toxic effect of ethyl alcohol|ETHANOL
Drug|Organic Chemical|SIMPLE_SEGMENT|8323,8330|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8323,8330|false|false|false|C0001962;C3854029;C3854030|CNS depressants ethanol;antiseptics ethanol;ethanol|ETHANOL
Event|Event|SIMPLE_SEGMENT|8323,8330|false|false|false|||ETHANOL
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8323,8330|false|false|false|C0202304|Ethanol measurement|ETHANOL
Event|Event|SIMPLE_SEGMENT|8331,8334|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|8331,8334|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|8345,8348|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|8345,8348|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|8360,8363|false|false|false|||NEG
Finding|Finding|SIMPLE_SEGMENT|8360,8363|false|false|false|C5848551|Neg - answer|NEG
Event|Event|SIMPLE_SEGMENT|8365,8368|false|false|false|||EEG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8365,8368|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|SIMPLE_SEGMENT|8389,8399|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|8389,8399|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|8389,8399|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|8406,8415|false|false|false|||telemetry
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8406,8415|false|false|false|C0039451|Telemetry|telemetry
Event|Event|SIMPLE_SEGMENT|8416,8424|false|false|false|||captured
Event|Event|SIMPLE_SEGMENT|8439,8450|false|false|false|||activations
Event|Event|SIMPLE_SEGMENT|8457,8467|false|false|false|||background
Finding|Conceptual Entity|SIMPLE_SEGMENT|8457,8467|false|false|false|C1706907|Background|background
Event|Event|SIMPLE_SEGMENT|8468,8474|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|8482,8488|false|false|false|||waking
Finding|Physiologic Function|SIMPLE_SEGMENT|8482,8488|false|false|false|C0442696|Waking|waking
Drug|Organic Chemical|SIMPLE_SEGMENT|8493,8498|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8493,8498|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|SIMPLE_SEGMENT|8493,8498|false|false|false|C0037313|Sleep|sleep
Event|Event|SIMPLE_SEGMENT|8499,8507|false|false|false|||patterns
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|8530,8543|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|8530,8543|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|8530,8543|true|false|false|C0000769|teratologic|abnormalities
Event|Event|SIMPLE_SEGMENT|8558,8566|false|false|false|||features
Event|Event|SIMPLE_SEGMENT|8587,8595|false|false|false|||seizures
Finding|Sign or Symptom|SIMPLE_SEGMENT|8587,8595|false|false|false|C0036572|Seizures|seizures
Event|Event|SIMPLE_SEGMENT|8599,8610|false|false|false|||bradycardia
Finding|Finding|SIMPLE_SEGMENT|8599,8610|false|false|false|C0428977;C3812171|Bradycardia;Bradycardia by ECG Finding|bradycardia
Event|Event|SIMPLE_SEGMENT|8615,8620|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|8624,8631|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|8624,8631|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8624,8631|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|8642,8645|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|8642,8645|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8642,8645|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|8642,8645|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8642,8651|false|false|false|C4028269|Nuclear magnetic resonance imaging brain|MRI BRAIN
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8646,8651|false|false|false|C0006104;C4266577|Brain;Head>Brain|BRAIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8646,8651|false|false|false|C0006111|Brain Diseases|BRAIN
Event|Event|SIMPLE_SEGMENT|8646,8651|false|false|false|||BRAIN
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8665,8673|true|false|false|C0009924|Contrast Media|CONTRAST
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8679,8687|false|false|false|C2926606||FINDINGS
Event|Event|SIMPLE_SEGMENT|8679,8687|false|false|false|||FINDINGS
Finding|Functional Concept|SIMPLE_SEGMENT|8679,8687|false|false|false|C2607943|findings aspects|FINDINGS
Drug|Organic Chemical|SIMPLE_SEGMENT|8701,8706|false|false|false|C0309093|FLAIR (product)|FLAIR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8701,8706|false|false|false|C0309093|FLAIR (product)|FLAIR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8701,8706|false|false|false|C2826145|Fluid Attenuated Inversion Recovery|FLAIR
Event|Event|SIMPLE_SEGMENT|8707,8718|false|false|false|||hypointense
Finding|Idea or Concept|SIMPLE_SEGMENT|8726,8736|false|false|false|C1517605|Isointense|isointense
Event|Event|SIMPLE_SEGMENT|8737,8743|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|8737,8743|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|8737,8743|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Cell Component|SIMPLE_SEGMENT|8747,8754|false|false|false|C1660780|midline cell component|midline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8769,8777|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|8769,8777|false|false|false|||anterior
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8782,8791|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8782,8801|false|false|false|C0032009;C0447640|Pituitary Gland, Posterior;pars nervosa of hypophysis|posterior pituitary
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Hormone|SIMPLE_SEGMENT|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8782,8801|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8792,8801|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8792,8801|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|SIMPLE_SEGMENT|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|SIMPLE_SEGMENT|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8792,8801|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Event|Event|SIMPLE_SEGMENT|8792,8801|false|false|false|||pituitary
Event|Event|SIMPLE_SEGMENT|8805,8810|false|false|false|||noted
Event|Event|SIMPLE_SEGMENT|8824,8832|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|8824,8832|true|false|false|C3887511|Evidence|evidence
Event|Event|SIMPLE_SEGMENT|8838,8848|false|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|8838,8848|false|false|false|C0019080|Hemorrhage|hemorrhage
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8850,8855|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|8850,8855|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|8850,8855|false|false|false|C0013604|Edema|edema
Finding|Finding|SIMPLE_SEGMENT|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|SIMPLE_SEGMENT|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|SIMPLE_SEGMENT|8857,8861|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|SIMPLE_SEGMENT|8857,8868|false|false|false|C4086564|Mass Effect|mass effect
Event|Event|SIMPLE_SEGMENT|8862,8868|false|false|false|||effect
Anatomy|Cell Component|SIMPLE_SEGMENT|8870,8877|false|false|false|C1660780|midline cell component|midline
Finding|Finding|SIMPLE_SEGMENT|8870,8883|false|false|false|C4086580|Midline Shift|midline shift
Event|Event|SIMPLE_SEGMENT|8878,8883|false|false|false|||shift
Finding|Functional Concept|SIMPLE_SEGMENT|8878,8883|false|false|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|8878,8883|false|false|false|C2347509|Physical Shift|shift
Event|Event|SIMPLE_SEGMENT|8887,8897|false|false|false|||infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|8887,8897|false|false|false|C0021308|Infarction|infarction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8904,8914|false|false|false|C0018827|Heart Ventricle|ventricles
Event|Event|SIMPLE_SEGMENT|8919,8924|false|false|false|||sulci
Event|Event|SIMPLE_SEGMENT|8929,8935|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|8939,8946|false|false|false|||caliber
Event|Event|SIMPLE_SEGMENT|8951,8964|false|false|false|||configuration
Finding|Conceptual Entity|SIMPLE_SEGMENT|8951,8964|false|false|false|C2827597|Computer Configuration|configuration
Finding|Finding|SIMPLE_SEGMENT|8979,8987|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|SIMPLE_SEGMENT|8979,8987|true|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Event|Activity|SIMPLE_SEGMENT|8988,8999|true|false|false|C2349975|Enhance (action)|enhancement
Event|Event|SIMPLE_SEGMENT|8988,8999|false|false|false|||enhancement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8988,8999|true|false|false|C1627358|Refractive surgery enhancement|enhancement
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9006,9014|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|9015,9029|false|false|false|||administration
Event|Occupational Activity|SIMPLE_SEGMENT|9015,9029|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9015,9029|false|false|false|C1533734|Administration (procedure)|administration
Event|Event|SIMPLE_SEGMENT|9035,9045|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|9035,9045|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|9035,9045|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Drug|Organic Chemical|SIMPLE_SEGMENT|9059,9064|false|false|false|C0309093|FLAIR (product)|FLAIR
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9059,9064|false|false|false|C0309093|FLAIR (product)|FLAIR
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9059,9064|false|false|false|C2826145|Fluid Attenuated Inversion Recovery|FLAIR
Event|Event|SIMPLE_SEGMENT|9065,9076|false|false|false|||hypointense
Finding|Idea or Concept|SIMPLE_SEGMENT|9084,9094|false|false|false|C1517605|Isointense|isointense
Event|Event|SIMPLE_SEGMENT|9095,9101|false|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|9095,9101|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|9095,9101|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Cell Component|SIMPLE_SEGMENT|9105,9112|false|false|false|C1660780|midline cell component|midline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9127,9135|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|9127,9135|false|false|false|||anterior
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9140,9149|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9140,9159|false|false|false|C0032009;C0447640|Pituitary Gland, Posterior;pars nervosa of hypophysis|posterior pituitary
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Hormone|SIMPLE_SEGMENT|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9140,9159|false|false|false|C0032017;C3714635|Posterior Pituitary Hormone Drug Class;posterior pituitary hormones|posterior pituitary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9150,9159|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9150,9159|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|SIMPLE_SEGMENT|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|SIMPLE_SEGMENT|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9150,9159|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Finding|Finding|SIMPLE_SEGMENT|9160,9166|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9160,9166|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|9167,9177|false|false|false|||represents
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|9196,9200|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|9196,9200|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|9196,9200|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|9196,9200|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|SIMPLE_SEGMENT|9212,9222|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|9212,9222|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|9212,9222|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Event|Event|SIMPLE_SEGMENT|9226,9232|false|false|false|||needed
Event|Event|SIMPLE_SEGMENT|9234,9243|false|false|false|||dedicated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|9244,9253|false|false|false|C0032005|Pituitary Gland|pituitary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9244,9253|false|false|false|C0032002|Pituitary Diseases|pituitary
Drug|Hormone|SIMPLE_SEGMENT|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Organic Chemical|SIMPLE_SEGMENT|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9244,9253|false|false|false|C0304812|Pituitary hormone preparation|pituitary
Event|Event|SIMPLE_SEGMENT|9254,9256|false|false|false|||MR
Event|Event|SIMPLE_SEGMENT|9265,9273|false|false|false|||obtained
Finding|Intellectual Product|SIMPLE_SEGMENT|9282,9287|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|9288,9296|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9288,9303|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|9288,9303|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Intellectual Product|SIMPLE_SEGMENT|9309,9318|false|false|false|C2349155|Worksheet|worksheet
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9321,9332|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9321,9332|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|9321,9332|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|9321,9332|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|9321,9345|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|9336,9345|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9336,9345|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|9347,9357|false|false|false|C0015620|famotidine|famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9347,9357|false|false|false|C0015620|famotidine|famotidine
Event|Event|SIMPLE_SEGMENT|9347,9357|false|false|false|||famotidine
Finding|Finding|SIMPLE_SEGMENT|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Finding|Intellectual Product|SIMPLE_SEGMENT|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Finding|Organism Function|SIMPLE_SEGMENT|9370,9375|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|birth
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9370,9383|false|false|false|C0700589|Contraceptive methods|birth control
Drug|Organic Chemical|SIMPLE_SEGMENT|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|SIMPLE_SEGMENT|9376,9383|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|SIMPLE_SEGMENT|9376,9383|false|false|false|||control
Finding|Conceptual Entity|SIMPLE_SEGMENT|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|SIMPLE_SEGMENT|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|SIMPLE_SEGMENT|9376,9383|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|SIMPLE_SEGMENT|9435,9445|false|false|false|C0015620|famotidine|Famotidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9435,9445|false|false|false|C0015620|famotidine|Famotidine
Drug|Organic Chemical|SIMPLE_SEGMENT|9467,9477|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9467,9477|false|false|false|C0025859|metoprolol|Metoprolol
Event|Event|SIMPLE_SEGMENT|9467,9477|false|false|false|||Metoprolol
Drug|Organic Chemical|SIMPLE_SEGMENT|9467,9486|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9467,9486|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9478,9486|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9478,9486|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Organic Chemical|SIMPLE_SEGMENT|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|9510,9523|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|9510,9523|false|false|false|||Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|9526,9534|false|false|false|C0026162|Minerals|minerals
Event|Event|SIMPLE_SEGMENT|9526,9534|false|false|false|||minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9537,9540|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|9537,9540|false|false|false|||TAB
Finding|Intellectual Product|SIMPLE_SEGMENT|9614,9618|false|false|false|C1720092|Once - dosing instruction fragment|ONCE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9620,9629|false|false|false|C3854082||Prognosis
Event|Event|SIMPLE_SEGMENT|9620,9629|false|false|false|||Prognosis
Procedure|Health Care Activity|SIMPLE_SEGMENT|9620,9629|false|false|false|C0033325|Forecast of outcome|Prognosis
Finding|Idea or Concept|SIMPLE_SEGMENT|9631,9635|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|Good
Event|Activity|SIMPLE_SEGMENT|9666,9670|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|9666,9670|false|false|false|C2828567|PRSS30P gene|Disp
Event|Event|SIMPLE_SEGMENT|9680,9687|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|9680,9687|false|false|false|C0807726|refill|Refills
Event|Event|SIMPLE_SEGMENT|9695,9704|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9695,9704|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9695,9704|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9695,9716|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|9695,9716|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9705,9716|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|9705,9716|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|9705,9716|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|9718,9726|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|9718,9726|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|9718,9731|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|9727,9731|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|9727,9731|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|9727,9731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|9727,9731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|9734,9742|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|9734,9742|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|9750,9759|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9750,9759|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9750,9759|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|9750,9769|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9760,9769|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|9760,9769|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|9760,9769|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|9760,9769|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9760,9769|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Conceptual Entity|SIMPLE_SEGMENT|9771,9781|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Finding|Functional Concept|SIMPLE_SEGMENT|9771,9781|false|false|false|C0205245;C0542341;C2700217|Function (attribute);Functional;Functional Relationship|Functional
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9795,9803|false|false|false|C0039082|Syndrome|syndrome
Event|Event|SIMPLE_SEGMENT|9795,9803|false|false|false|||syndrome
Event|Event|SIMPLE_SEGMENT|9808,9817|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9808,9817|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9808,9817|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9808,9817|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9808,9817|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9818,9827|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9818,9827|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|9818,9827|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|9818,9827|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|9829,9835|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9829,9842|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|9829,9842|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9836,9842|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9836,9842|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9844,9849|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|9844,9849|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|9854,9862|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|9854,9862|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|9864,9869|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9864,9886|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|9864,9886|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|9873,9886|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|9873,9886|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|9873,9886|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Event|Event|SIMPLE_SEGMENT|9888,9897|false|false|false|||Lethargic
Finding|Sign or Symptom|SIMPLE_SEGMENT|9888,9897|false|false|false|C0023380|Lethargy|Lethargic
Event|Event|SIMPLE_SEGMENT|9902,9911|false|false|false|||arousable
Event|Activity|SIMPLE_SEGMENT|9913,9921|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|9913,9921|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|9913,9921|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9922,9928|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|9922,9928|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|9922,9928|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|9930,9940|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|9930,9940|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|9930,9940|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|9943,9954|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|9943,9954|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|9943,9954|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|9959,9968|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|9959,9968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9959,9968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9959,9968|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9959,9968|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9959,9981|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9959,9981|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|9959,9981|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|9969,9981|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|9969,9981|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|9969,9981|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|9983,9987|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|10007,10015|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|10007,10015|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|10007,10015|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|10023,10027|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|10023,10027|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|10023,10027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10023,10027|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|10023,10030|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|SIMPLE_SEGMENT|10065,10073|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10085,10093|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|10085,10093|false|false|false|C0018681|Headache|headache
Event|Event|SIMPLE_SEGMENT|10095,10103|false|false|false|||lethargy
Finding|Sign or Symptom|SIMPLE_SEGMENT|10095,10103|false|false|false|C0023380|Lethargy|lethargy
Event|Event|SIMPLE_SEGMENT|10110,10118|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10110,10118|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Drug|Biologically Active Substance|SIMPLE_SEGMENT|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10128,10132|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10128,10132|false|false|false|C0337439|Iron measurement|iron
Event|Event|SIMPLE_SEGMENT|10133,10141|false|false|false|||infusion
Finding|Functional Concept|SIMPLE_SEGMENT|10133,10141|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10133,10141|false|false|false|C0574032|Infusion procedures|infusion
Event|Event|SIMPLE_SEGMENT|10154,10160|false|false|false|||number
Finding|Idea or Concept|SIMPLE_SEGMENT|10154,10160|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Event|SIMPLE_SEGMENT|10164,10169|false|false|false|||tests
Finding|Intellectual Product|SIMPLE_SEGMENT|10164,10169|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10164,10169|false|false|false|C0022885|Laboratory Procedures|tests
Finding|Idea or Concept|SIMPLE_SEGMENT|10187,10195|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10216,10226|false|false|false|||reassuring
Procedure|Health Care Activity|SIMPLE_SEGMENT|10216,10226|false|false|false|C0557055|Reassuring (procedure)|reassuring
Event|Event|SIMPLE_SEGMENT|10231,10234|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|10231,10234|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10231,10234|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|10231,10234|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10243,10248|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10243,10248|false|false|false|C0006111|Brain Diseases|brain
Event|Event|SIMPLE_SEGMENT|10249,10255|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|10259,10267|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|10259,10267|true|false|false|C3887511|Evidence|evidence
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10272,10278|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|10272,10278|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|10272,10278|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|SIMPLE_SEGMENT|10282,10294|false|false|false|||inflammation
Finding|Pathologic Function|SIMPLE_SEGMENT|10282,10294|false|false|false|C0021368|Inflammation|inflammation
Event|Event|SIMPLE_SEGMENT|10299,10302|false|false|false|||EEG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10299,10302|false|false|false|C0013819|Electroencephalography|EEG
Event|Event|SIMPLE_SEGMENT|10306,10313|false|false|false|||monitor
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|10319,10324|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10319,10324|false|false|false|C0006111|Brain Diseases|brain
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|10319,10330|false|false|false|C0678909|Brain Waves|brain waves
Event|Event|SIMPLE_SEGMENT|10325,10330|false|false|false|||waves
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|10325,10330|false|false|false|C0678544||waves
Event|Event|SIMPLE_SEGMENT|10332,10338|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|10342,10350|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|10342,10350|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|10342,10353|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|10354,10361|false|false|false|||seizure
Finding|Sign or Symptom|SIMPLE_SEGMENT|10354,10361|true|false|false|C0036572|Seizures|seizure
Event|Event|SIMPLE_SEGMENT|10368,10376|false|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|10368,10376|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|SIMPLE_SEGMENT|10387,10395|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|10421,10436|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|10421,10436|false|false|false|C0019993|Hospitalization|hospitalization
Event|Event|SIMPLE_SEGMENT|10446,10454|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|10459,10466|false|false|false|||improve
Event|Event|SIMPLE_SEGMENT|10477,10482|false|false|false|||leave
Event|Event|SIMPLE_SEGMENT|10487,10495|false|false|false|||hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|10487,10495|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10505,10512|false|false|false|||leaving
Finding|Idea or Concept|SIMPLE_SEGMENT|10517,10525|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|10538,10546|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|10550,10554|false|false|false|||work
Event|Event|SIMPLE_SEGMENT|10559,10568|false|false|false|||improving
Event|Event|SIMPLE_SEGMENT|10574,10582|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|10574,10582|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|10592,10599|false|false|false|||improve
Event|Event|SIMPLE_SEGMENT|10615,10619|false|false|false|||work
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10644,10648|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|SIMPLE_SEGMENT|10644,10648|false|false|false|||best
Finding|Gene or Genome|SIMPLE_SEGMENT|10644,10648|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|SIMPLE_SEGMENT|10659,10663|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|10659,10663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|10659,10663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10659,10668|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|10659,10668|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|10671,10679|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10680,10692|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|10680,10692|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|10680,10692|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

