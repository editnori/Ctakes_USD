CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Has difficulty doing (qualifier value)|Finding|false|false||Difficultynull|Inspiration (function)|Finding|false|false||in breathingnull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|History of present illness (finding)|Finding|true|false||History of Present Illnessnull|null|Attribute|true|false||History of Present Illnessnull|Medical History|Finding|true|false||History ofnull|History of present illness (finding)|Finding|true|false||History
null|History of previous events|Finding|true|false||History
null|Historical aspects qualifier|Finding|true|false||History
null|Medical History|Finding|true|false||History
null|Concept History|Finding|true|false||Historynull|History|Subject|true|false||Historynull|Present illness|Finding|true|false||Present Illnessnull|Present|Finding|true|false||Present
null|Presentation|Finding|true|false||Presentnull|Illness (finding)|Finding|true|false||Illnessnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|null|Disorder|false|false||NSCLCnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Usual|Modifier|false|false||usualnull|personal health|Finding|false|false||state of healthnull|State|Finding|false|false||statenull|Geographic state|Entity|false|false||state
null|US State|Entity|false|false||statenull|Health|Finding|false|false||healthnull|Evening|Time|false|false||eveningnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Somewhat|Finding|false|false||somewhatnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Breath|Finding|false|false||breathnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Morning|Time|false|false||morningnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Illness (finding)|Finding|true|false||sicknull|Contacts|Procedure|true|false||contactsnull|Recent|Time|true|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Sedentary lifestyle|Finding|false|false||sedentary lifestylenull|Sedentary lifestyle|Finding|false|false||sedentarynull|Sedentary|Modifier|false|false||sedentarynull|Life Style|Finding|false|false||lifestylenull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Fever symptoms (finding)|Finding|true|false||fever
null|Fever|Finding|true|false||fevernull|Chills|Finding|true|false||chillsnull|Dizziness|Finding|false|false||dizziness
null|Vertigo|Finding|false|false||dizzinessnull|Lightheadedness|Finding|false|false||lightheadednessnull|Syncope|Finding|false|false||syncopenull|Syncope <Gastrophryninae>|Entity|false|false||syncopenull|Hypoxia|Finding|false|false||hypoxicnull|on room air|Finding|false|false||on room airnull|Room Air|Drug|false|false||room airnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|short-acting thyroid stimulator|Drug|false|false||sats
null|short-acting thyroid stimulator|Drug|false|false||satsnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Unsuccessful|Modifier|false|false||unsuccessfulnull|Apyrexial|Finding|false|false||afebrilenull|Leukocytes|Anatomy|false|false||WBCnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture (Anthropological)|Finding|false|false||culturesnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Injection of antibiotic|Procedure|false|false||antibiotic administrationnull|Antibiotics|Drug|false|false||antibioticnull|Administration (procedure)|Procedure|false|false||administrationnull|Administration occupational activities|Event|false|false||administrationnull|Plain chest X-ray|Procedure|true|false||CXRnull|Peptide Nucleic Acids|Drug|true|false||PNAnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Known|Modifier|false|false||knownnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|CAT scan of head|Procedure|true|false||CT headnull|null|Attribute|true|false||CT headnull|Problems with head|Disorder|true|false||headnull|Procedure on head|Procedure|true|false||headnull|Structure of head of caudate nucleus|Anatomy|true|false||head
null|Head|Anatomy|true|false||headnull|Head Device|Device|true|false||headnull|Metastatic malignant neoplasm|Disorder|true|false||metastases
null|Neoplasm Metastasis|Disorder|true|false||metastasesnull|Metastatic Lesion|Finding|true|false||metastasesnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Patient Transfer|Procedure|false|false||transfer, patientnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|null|Device|false|false||NRBnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Inventory of Callous-Unemotional Traits|Finding|false|false||ICUnull|Structure of intraculminate fissure|Anatomy|false|false||ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Feeling comfortable|Finding|false|false||comfortablenull|short-acting thyroid stimulator|Drug|false|false||Sats
null|short-acting thyroid stimulator|Drug|false|false||Satsnull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Flow|Phenomenon|false|false||flownull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Tent - Recreation Equipment|Device|false|false||tentnull|Reactive Oxygen Species|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|rosiglitazone|Drug|false|false||ROS
null|Reactive Oxygen Species|Drug|false|false||ROSnull|ROS1 wt Allele|Finding|false|false||ROS
null|ROS1 gene|Finding|false|false||ROSnull|Review of systems (procedure)|Procedure|false|false||ROSnull|rostral sulcus|Anatomy|false|false||ROSnull|Relationship modifier - Patient|Finding|true|false||patient
null|Specimen Type - Patient|Finding|true|false||patient
null|Mail Claim Party - Patient|Finding|true|false||patient
null|Report source - Patient|Finding|true|false||patient
null|null|Finding|true|false||patient
null|Disabled Person Code - Patient|Finding|true|false||patientnull|Patients|Subject|true|false||patientnull|Veterinary Patient|Entity|true|false||patientnull|Fever|Finding|true|false||feversnull|Chills|Finding|true|false||chillsnull|Body Weight Changes|Finding|true|false||weight changenull|infant weight for previous delivery (history)|Finding|true|false||weight
null|Weight symptom (finding)|Finding|true|false||weightnull|Weighing patient|Procedure|true|false||weightnull|null|Attribute|true|false||weightnull|Body Weight|Subject|true|false||weightnull|Importance Weight|Modifier|true|false||weightnull|Weight|LabModifier|true|false||weightnull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Abdominal Pain|Finding|false|false||abdominal painnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Constipation|Finding|false|false||constipationnull|Melena|Finding|false|false||melenanull|Hematochezia|Disorder|false|false||hematochezianull|Blood in stool|Finding|false|false||hematochezianull|Chest Pain|Finding|false|false||chest painnull|null|Attribute|false|false||chest painnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|sleeping upright or using specific number of extra pillows (orthopnea)|Finding|false|false||orthopnea
null|Orthopnea|Finding|false|false||orthopneanull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Peripheral edema|Finding|false|false||extremity edemanull|Limb structure|Anatomy|false|false||extremitynull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Increased frequency of micturition|Finding|false|false||urinary frequencynull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|Frequency|Finding|false|false||frequency
null|How Often|Finding|false|false||frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Urgent|Modifier|false|false||urgencynull|Dysuria|Finding|false|false||dysurianull|Lightheadedness|Finding|false|false||lightheadednessnull|Gait|Finding|false|false||gaitnull|General unsteadiness|Finding|false|false||unsteadinessnull|Focal|Modifier|false|false||focalnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Vision|Finding|false|false||visionnull|null|Attribute|false|false||visionnull|Specialized Stand Alone Plan - Vision|Entity|false|false||visionnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Headache|Finding|false|false||headachenull|Eruption of skin (disorder)|Disorder|true|false||rashnull|Skin rash|Finding|true|false||rash
null|Eruptions|Finding|true|false||rash
null|Exanthema|Finding|true|false||rashnull|Skin symptom change|Finding|false|false||skin changesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||skinnull|Skin Specimen Source Code|Finding|false|false||skin
null|Skin Specimen|Finding|false|false||skinnull|Skin, Human|Anatomy|false|false||skin
null|Skin|Anatomy|false|false||skinnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Cyclophosphamide/Doxorubicin/Vincristine|Drug|false|false||CVAnull|Acute ill-defined cerebrovascular disease|Disorder|false|false||CVA
null|Cerebrovascular accident|Disorder|false|false||CVAnull|Small|LabModifier|false|false||smallnull|Left posterior|Modifier|false|false||left posteriornull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Coronal (qualifier value)|Modifier|false|false||frontalnull|Infarction|Finding|false|false||infarctnull|Age related macular degeneration|Disorder|false|false||Macular Degeneration
null|Macular degeneration|Disorder|false|false||Macular Degenerationnull|macular|Modifier|false|false||Macularnull|biologic degeneration|Finding|false|false||Degeneration
null|Abnormal degeneration|Finding|false|false||Degenerationnull|null|Disorder|false|false||NSCLCnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Neoplasms|Disorder|false|false||oncologynull|oncology services|Procedure|false|false||oncologynull|oncology (field)|Title|false|false||oncologynull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Right sided|Modifier|false|false||right-sidednull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pulmonary (intended site)|Finding|false|false||pulmonarynull|Lung|Anatomy|false|false||pulmonarynull|null|Attribute|false|false||pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|Unrelated (finding)|Finding|false|false||unrelatednull|Unrelated to Intervention|Modifier|false|false||unrelatednull|Myocardial Infarction|Disorder|false|false||myocardial infarctionnull|null|Attribute|false|false||myocardial infarctionnull|Myocardium|Anatomy|false|false||myocardialnull|Myocardial|Modifier|false|false||myocardialnull|Infarction|Finding|false|false||infarctionnull|Adenocarcinoma|Disorder|false|false||adenocarcinoma
null|Malignant adenomatous neoplasm|Disorder|false|false||adenocarcinomanull|Patterns|Modifier|false|false||patternnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Participation Type - origin|Finding|false|false||origin
null|National origin|Finding|false|false||originnull|Beginning|Time|false|false||originnull|KRT7 wt Allele|Finding|false|false||CK7
null|KRT7 gene|Finding|false|false||CK7null|thyroid transcription factor 1|Drug|false|false||TTF-1
null|thyroid transcription factor 1|Drug|false|false||TTF-1
null|NKX2-1 protein, human|Drug|false|false||TTF-1
null|NKX2-1 protein, human|Drug|false|false||TTF-1
null|TTF1 protein, human|Drug|false|false||TTF-1
null|TTF1 protein, human|Drug|false|false||TTF-1null|NKX2-1 wt Allele|Finding|false|false||TTF-1
null|TTF1 wt Allele|Finding|false|false||TTF-1
null|NKX2-1 gene|Finding|false|false||TTF-1null|RHOH wt Allele|Finding|false|false||TTF
null|RHOH gene|Finding|false|false||TTFnull|Tumour treating fields therapy|Procedure|false|false||TTFnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Metastatic non-small cell lung cancer|Disorder|false|false||stage IV nonsmall cell lung cancernull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Numerous|LabModifier|false|false||multiplenull|Intrapulmonary Route of Administration|Finding|false|false||intrapulmonarynull|Intrapulmonary|Modifier|false|false||intrapulmonarynull|Lesion|Finding|false|false||lesionsnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Central Nervous System Involvement|Finding|true|false||central nervous system involvementnull|CENTRAL NERVOUS SYSTEM DIAGNOSTIC RADIOPHARMACEUTICALS|Drug|true|false||central nervous systemnull|Central Nervous System|Anatomy|true|false||central nervous systemnull|Central brand of multivitamin with minerals|Drug|true|false||central
null|Central brand of multivitamin with minerals|Drug|true|false||centralnull|Central Minus|Procedure|true|false||centralnull|Central|Modifier|true|false||centralnull|NERVOUS SYSTEM DRUGS|Drug|true|false||nervous systemnull|Nervous system structure|Anatomy|true|false||nervous systemnull|Nervous - anatomy qualifier|Finding|true|false||nervous
null|Nervousness|Finding|true|false||nervousnull|System (basic dose form)|Drug|false|false||systemnull|System, LOINC Axis 4|Finding|false|false||system
null|System|Finding|false|false||systemnull|Device system|Device|false|false||system
null|System - kit|Device|false|false||systemnull|System (unit of presentation)|LabModifier|false|false||systemnull|Involvement with|Finding|false|false||involvementnull|Neoplasm Metastasis|Disorder|false|false||metastasis
null|Metastatic malignant neoplasm|Disorder|false|false||metastasisnull|Metastasis|Finding|false|false||metastasis
null|Metastatic Lesion|Finding|false|false||metastasisnull|Status post|Time|false|false||Status post
null|Post|Time|false|false||Status postnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|event cycle|Time|false|false||cyclesnull|pemetrexed|Drug|false|false||pemetrexed
null|pemetrexed|Drug|false|false||pemetrexednull|mg/m2|LabModifier|false|false||mg/m2null|Course|Time|false|false||coursenull|Cytopenia|Disorder|false|false||cytopeniasnull|Cytopenia (finding)|Finding|false|false||cytopeniasnull|Growth and Development function|Finding|false|false||development
null|development aspects|Finding|false|false||development
null|biological development|Finding|false|false||development
null|Development|Finding|false|false||developmentnull|Creatinine increased|Finding|false|false||increased creatinine
null|Serum creatinine raised|Finding|false|false||increased creatininenull|Finding of creatinine level|Finding|false|false||creatinine levelsnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Levels (qualifier value)|Modifier|false|false||levelsnull|Chest CT|Procedure|false|false||Chest CTnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|ITMIG MRECIST Partial Response|Finding|false|false||partial response
null|irPR (Immune-Related Response Criteria)|Finding|false|false||partial response
null|IMWG Partial Response|Finding|false|false||partial response
null|partial response|Finding|false|false||partial response
null|RECIL PR|Finding|false|false||partial responsenull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Communication Response|Finding|false|false||response
null|Disease Response|Finding|false|false||response
null|Answer (statement)|Finding|false|false||responsenull|Response process|Subject|false|false||responsenull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Improvement|Finding|false|false||improvementnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Upper|Modifier|false|false||superiornull|Anatomical segmentation|Modifier|false|false||segmentnull|Structure of right lower lobe of lung|Anatomy|false|false||right lower lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|density|LabModifier|false|false||densitiesnull|Structure of left lower lobe of lung|Anatomy|false|false||left lower lobenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Still|Disorder|false|false||Stillnull|bacitracin|Drug|false|false||BAC
null|bacitracin|Drug|false|false||BACnull|Bronchioloalveolar Adenocarcinoma|Disorder|false|false||BACnull|Blood alcohol concentration|Finding|false|false||BACnull|BAC Regimen|Procedure|false|false||BACnull|polyhedral organelle|Anatomy|false|false||BACnull|Bacterial Artificial Chromosomes|Device|false|false||BACnull|Chest CT|Procedure|false|false||CT Chestnull|null|Attribute|false|false||CT Chestnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Density above reference range|Finding|false|false||increased density
null|Decreased translucency|Finding|false|false||increased densitynull|density|LabModifier|false|false||densitynull|Structure of right lower lobe of lung|Anatomy|false|false||right lower lobenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glassnull|Chromosome 2q32-Q33 Deletion Syndrome|Disorder|false|false||glassnull|Glass Packaging Device|Device|false|false||glass
null|Glass (substance)|Device|false|false||glassnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacities
null|Decreased translucency|Finding|false|false||opacitiesnull|Lingula of cerebellum|Anatomy|false|false||lingula
null|Lingula|Anatomy|false|false||lingula
null|Lingula of left lung|Anatomy|false|false||lingulanull|Lingula <Lingulidae>|Entity|false|false||lingulanull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Much|Finding|false|false||muchnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Chest CT|Procedure|false|false||Chest CTnull|Chest problem|Finding|false|false||Chestnull|Chest|Anatomy|false|false||Chest
null|Anterior thoracic region|Anatomy|false|false||Chestnull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|Parameterized Data Type - Interval|Finding|true|false||intervalnull|Interval|Time|true|false||intervalnull|Disease Progression|Finding|true|false||progression
null|Progression|Finding|true|false||progressionnull|Known|Modifier|true|false||knownnull|Disease|Disorder|true|false||diseasenull|Query Status Code - new|Finding|true|false||new
null|Act Status - new|Finding|true|false||newnull|Newar Language|Entity|true|false||newnull|New|Modifier|true|false||newnull|Site|Modifier|true|false||sitesnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Indirect exposure mechanism - Father|Finding|false|false||father
null|Relationship - Father|Finding|false|false||father
null|Father - courtesy title|Finding|false|false||fathernull|Father (person)|Subject|false|false||fathernull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Relationship - Mother|Finding|false|false||mothernull|Mother (person)|Subject|false|false||mothernull|Neoplasm of uncertain or unknown behavior of stomach|Disorder|false|false||stomach
null|Stomach Diseases|Disorder|false|false||stomach
null|Benign neoplasm of stomach|Disorder|false|false||stomach
null|Carcinoma in situ of stomach|Disorder|false|false||stomachnull|Stomach problem|Finding|false|false||stomachnull|Procedure on stomach|Procedure|false|false||stomachnull|Stomach structure|Anatomy|false|false||stomach
null|Abdomen>Stomach|Anatomy|false|false||stomach
null|Stomach|Anatomy|false|false||stomachnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Osteosarcoma of bone|Disorder|false|false||osteosarcoma
null|Osteosarcoma|Disorder|false|false||osteosarcomanull|RB1 gene|Finding|false|false||osteosarcomanull|Medical History|Finding|true|false||history ofnull|History of present illness (finding)|Finding|true|false||history
null|History of previous events|Finding|true|false||history
null|Historical aspects qualifier|Finding|true|false||history
null|Medical History|Finding|true|false||history
null|Concept History|Finding|true|false||historynull|History|Subject|true|false||historynull|Malignant neoplasm of lung|Disorder|true|false||lung cancer
null|Carcinoma of lung|Disorder|true|false||lung cancernull|Lung diseases|Disorder|true|false||lungnull|Lung Problem|Finding|true|false||lungnull|Chest>Lung|Anatomy|true|false||lung
null|Lung|Anatomy|true|false||lungnull|Malignant tumor of colon|Disorder|true|false||cancer, colonnull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|true|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Malignant tumor of colon|Disorder|true|false||colon cancer
null|Malignant neoplasm of large intestine|Disorder|true|false||colon cancer
null|Colon Carcinoma|Disorder|true|false||colon cancernull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false||colon
null|Colonic Diseases|Disorder|true|false||colon
null|Carcinoma in situ of colon|Disorder|true|false||colonnull|COLON PROBLEM|Finding|true|false||colonnull|Colon structure (body structure)|Anatomy|true|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|true|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|Malignant Neoplasms|Disorder|true|false||cancernull|Specialty Type - cancer|Title|true|false||cancernull|Cancer <Cancridae>|Entity|true|false||cancernull|Malignant neoplasm of breast|Disorder|false|false||breast cancer
null|Breast Carcinoma|Disorder|false|false||breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|On admission|Time|false|false||On Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|Face tent oxygen delivery device|Device|false|false||face tentnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false||facenull|FANCE wt Allele|Finding|false|false||face
null|FANCE gene|Finding|false|false||face
null|ELOVL6 gene|Finding|false|false||facenull|Head>Face|Anatomy|false|false||face
null|Face|Anatomy|false|false||facenull|Face (spatial concept)|Modifier|false|false||facenull|Tent - Recreation Equipment|Device|false|false||tentnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GEN
null|GEN1 wt Allele|Finding|false|false||GEN
null|GEN1 gene|Finding|false|false||GENnull|Well (answer to question)|Finding|true|false||Wellnull|Well (container)|Device|true|false||Wellnull|Microplate Well|Modifier|true|false||Well
null|Good|Modifier|true|false||Well
null|Healthy|Modifier|true|false||Wellnull|Females|Subject|true|false||female
null|Woman|Subject|true|false||femalenull|Female, Self-Report|Modifier|true|false||female
null|Female Phenotype|Modifier|true|false||femalenull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|true|false||HEENTnull|Pupil equal round and reacting to light|Finding|false|false||PERRLnull|Scleral Diseases|Disorder|false|false||scleranull|examination of sclera|Procedure|false|false||scleranull|Sclera|Anatomy|false|false||scleranull|Anicteric|Finding|false|false||anictericnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Passive joint movement of neck (finding)|Finding|false|false||NECK
null|Neck problem|Finding|false|false||NECKnull|dendritic spine neck|Anatomy|false|false||NECK
null|Neck|Anatomy|false|false||NECKnull|Jugular venous engorgement|Finding|true|false||JVDnull|Cervical lymphadenopathy|Disorder|true|false||cervical lymphadenopathynull|Swollen lymph nodes in the neck|Finding|true|false||cervical lymphadenopathynull|Neck|Anatomy|true|false||cervicalnull|Cervical|Modifier|true|false||cervicalnull|Lymphadenopathy|Disorder|true|false||lymphadenopathynull|Swollen Lymph Node|Finding|true|false||lymphadenopathynull|Carcinoma in situ of trachea|Disorder|true|false||trachea
null|Benign neoplasm of trachea|Disorder|true|false||trachea
null|Tracheal Diseases|Disorder|true|false||tracheanull|trachea findings|Finding|true|false||tracheanull|Procedure on trachea|Procedure|true|false||tracheanull|Neck+Chest>Trachea|Anatomy|true|false||trachea
null|Trachea|Anatomy|true|false||tracheanull|Trachea <Xyleninae>|Entity|true|false||tracheanull|midline cell component|Anatomy|true|false||midlinenull|Midline (qualifier value)|Modifier|true|false||midlinenull|cordycepin|Drug|true|false||COR
null|cordycepin|Drug|true|false||CORnull|Heart|Anatomy|true|false||CORnull|Cornish language|Entity|true|false||CORnull|Regular|Modifier|true|false||Regularnull|Amount type - Rate|Finding|true|false||ratenull|Rating (action)|Event|true|false||ratenull|Rate|LabModifier|true|false||ratenull|Rhythm|Finding|true|false||rhythm
null|rhythmic process (biological)|Finding|true|false||rhythmnull|Pulmonary ventilator management|Procedure|false|false||PULMnull|Decreased breath sounds|Finding|false|false||Decreased breath soundsnull|null|Attribute|false|false||breath sounds
null|Respiratory Sounds|Attribute|false|false||breath soundsnull|Breath|Finding|false|false||breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Faint - appearance|Finding|false|false||faint
null|Syncope|Finding|false|false||faintnull|Basilar Rales|Finding|false|false||crackles
null|Rales|Finding|false|false||cracklesnull|Language Ability Proficiency - Good|Finding|false|false||Good
null|Language Proficiency - Good|Finding|false|false||Goodnull|Specimen Quality - Good|Modifier|false|false||Good
null|Good|Modifier|false|false||Goodnull|Exertion|Finding|false|false||effortnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false||ABDnull|ABD (body structure)|Anatomy|false|false||ABD
null|Abdomen|Anatomy|false|false||ABDnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|LRRC4B gene|Finding|true|false||HSMnull|Hereditary Multiple Exostoses|Disorder|true|false||EXTnull|EXT1 wt Allele|Finding|true|false||EXT
null|EXT1 gene|Finding|true|false||EXTnull|Neurology speciality|Title|true|false||NEUROnull|Neurologic (qualifier value)|Modifier|true|false||NEUROnull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to person|Finding|false|false||oriented to personnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||SKIN
null|Skin and subcutaneous tissue disorders|Disorder|false|false||SKINnull|Skin Specimen Source Code|Finding|false|false||SKIN
null|Skin Specimen|Finding|false|false||SKINnull|Skin, Human|Anatomy|false|false||SKIN
null|Skin|Anatomy|false|false||SKINnull|yellow skin or eyes (symptom)|Finding|true|false||jaundice
null|Icterus|Finding|true|false||jaundice
null|jaundice|Finding|true|false||jaundicenull|Cyanosis|Finding|true|false||cyanosisnull|Gross (qualifier value)|Modifier|true|false||grossnull|Dermatitis|Disorder|true|false||dermatitisnull|Ecchymosis|Finding|true|false||ecchymosesnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||HGB
null|Hemoglobin|Drug|false|false||HGBnull|CYGB gene|Finding|false|false||HGBnull|Hemoglobin concentration|Lab|false|false||HGBnull|Hemopoietic stem cell transplant|Procedure|false|false||HCT
null|Hematocrit Measurement|Procedure|false|false||HCTnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Primed lymphocyte test|Procedure|false|false||PLTnull|Count Dosing Unit|LabModifier|false|false||COUNT
null|Count|LabModifier|false|false||COUNTnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Bands|Device|false|false||BANDSnull|Lymph|Finding|false|false||LYMPHSnull|Monos|Drug|false|false||MONOS
null|Mono-S|Drug|false|false||MONOS
null|Monos|Drug|false|false||MONOSnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||EOS
null|Familial eosinophilia|Disorder|false|false||EOSnull|PRSS33 gene|Finding|false|false||EOS
null|IKZF4 gene|Finding|false|false||EOSnull|Eos <Loriini>|Entity|false|false||EOSnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Tears (substance)|Finding|false|false||TEARDROPnull|Rukia ruki (organism)|Entity|false|false||TEARDROPnull|Tear Shape|Modifier|false|false||TEARDROPnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREA
null|urea|Drug|false|false||UREAnull|Urea measurement|Procedure|false|false||UREAnull|Sodium supplements|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|sodium|Drug|false|false||SODIUM
null|Sodium Drug Class|Drug|false|false||SODIUMnull|Sodium metabolic function|Finding|false|false||SODIUMnull|Sodium measurement|Procedure|false|false||SODIUMnull|Potassium Drug Class|Drug|false|false||POTASSIUM
null|Dietary Potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|potassium|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUM
null|Potassium supplement|Drug|false|false||POTASSIUMnull|Potassium metabolic function|Finding|false|false||POTASSIUMnull|Potassium measurement|Procedure|false|false||POTASSIUMnull|chloride ion|Drug|false|false||CHLORIDE
null|Chlorides|Drug|false|false||CHLORIDEnull|Chloride metabolic function|Finding|false|false||CHLORIDEnull|Chloride measurement|Procedure|false|false||CHLORIDEnull|Total|Modifier|false|false||TOTALnull|carbon dioxide|Drug|false|false||CO2
null|carbon dioxide|Drug|false|false||CO2null|MT-CO2 gene|Finding|false|false||CO2
null|null|Finding|false|false||CO2
null|C2 wt Allele|Finding|false|false||CO2null|blood anion gap (lab test)|Procedure|false|false||ANION GAP
null|Anion gap measurement|Procedure|false|false||ANION GAPnull|Anion Gap|Attribute|false|false||ANION GAPnull|Anion gap result|Lab|false|false||ANION GAPnull|Anions|Drug|false|false||ANIONnull|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|Ras GTPase-Activating Protein 1, Human|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAP
null|GTPase-Activating Proteins|Drug|false|false||GAPnull|RASA1 wt Allele|Finding|false|false||GAP
null|RASA1 gene|Finding|false|false||GAPnull|Gap (space)|Modifier|false|false||GAPnull|lactate|Drug|false|false||LACTATE
null|lactate|Drug|false|false||LACTATE
null|Lactates|Drug|false|false||LACTATEnull|Lactic acid measurement|Procedure|false|false||LACTATEnull|Mandibular right first molar mesial prosthesis|Device|false|false||30PMnull|Color of urine|Finding|false|false||URINE  COLORnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||COLOR
null|Coloring Excipient|Drug|false|false||COLORnull|color - solid dosage form|Modifier|false|false||COLOR
null|Color|Modifier|false|false||COLORnull|Color quantity|LabModifier|false|false||COLORnull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE  BLOODnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|Nitrites|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITE
null|nitrite ion|Drug|false|false||NITRITEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||PROTEIN
null|Proteins|Drug|false|false||PROTEINnull|Protein Info|Finding|false|false||PROTEINnull|Protein measurement|Procedure|false|false||PROTEINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSE
null|glucose|Drug|false|false||GLUCOSEnull|Glucose measurement|Procedure|false|false||GLUCOSEnull|Glucose^1.5H post dose glucagon|Lab|false|false||GLUCOSEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Ketones|Drug|false|false||KETONEnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|bilirubin preparation|Drug|false|false||BILIRUBIN
null|bilirubin preparation|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBIN
null|Bilirubin|Drug|false|false||BILIRUBINnull|Bilirubin, total measurement|Procedure|false|false||BILIRUBIN
null|blood bilirubin level test|Procedure|false|false||BILIRUBINnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Micro (prefix)|Finding|false|false||Micro
null|Microbiology - Laboratory Class|Finding|false|false||Micronull|Microbiology procedure|Procedure|false|false||Micronull|Unit Of Measure Prefix - micro|LabModifier|false|false||Micronull|Legionella urinary antigen|Procedure|false|false||Legionella Urinary Antigennull|Legionella|Entity|false|false||Legionellanull|Urinary tract|Anatomy|false|false||Urinarynull|urinary|Modifier|false|false||Urinarynull|Antigens|Drug|false|false||Antigennull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Negative|Finding|false|false||NEGATIVE FORnull|Rh Negative Blood Group|Finding|false|false||NEGATIVE
null|Negative|Finding|false|false||NEGATIVE
null|Negative Finding|Finding|false|false||NEGATIVEnull|Expression Negative|Lab|false|false||NEGATIVEnull|Negative - qualifier|Modifier|false|false||NEGATIVE
null|Negative Charge|Modifier|false|false||NEGATIVEnull|Negative Number|LabModifier|false|false||NEGATIVEnull|Legionella|Entity|true|false||LEGIONELLAnull|Serogroup|Finding|true|false||SEROGROUPnull|Antigens|Drug|true|false||ANTIGENnull|Portion of urine|Finding|false|false||Urine
null|null|Finding|false|false||Urine
null|Urine|Finding|false|false||Urine
null|In Urine|Finding|false|false||Urine
null|Urine specimen|Finding|false|false||Urinenull|Urine culture|Procedure|false|false||URINE CULTUREnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Scientific Study|Procedure|false|false||Studiesnull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Sinus rhythm|Finding|false|false||Sinus rhythm
null|null|Finding|false|false||Sinus rhythmnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false||Sinusnull|pathologic fistula|Disorder|false|false||Sinusnull|Sinus - general anatomical term|Anatomy|false|false||Sinus
null|Nasal sinus|Anatomy|false|false||Sinusnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Bilateral Prophylactic Mastectomy|Procedure|false|false||bpmnull|breaths per minute|LabModifier|false|false||bpm
null|beats per minute|LabModifier|false|false||bpmnull|Fracture of second cervical vertebra|Disorder|false|false||axisnull|Axis vertebra|Anatomy|false|false||axisnull|Genus Axis|Entity|false|false||axisnull|Axis|Modifier|false|false||axisnull|Interval|Time|false|false||intervalsnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|WASF1 gene|Finding|false|false||wavenull|null|Phenomenon|false|false||wavenull|Mental Depression|Disorder|false|false||depressionsnull|Plain chest X-ray|Procedure|false|false||CXRnull|Marital Status - Single|Finding|false|false||SINGLE
null|Unmarried|Finding|false|false||SINGLEnull|Singular|LabModifier|false|false||SINGLEnull|Views AP|Modifier|false|false||AP VIEWnull|View|Modifier|false|false||VIEWnull|Chest problem|Finding|false|false||CHESTnull|Chest|Anatomy|false|false||CHEST
null|Anterior thoracic region|Anatomy|false|false||CHESTnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Median (qualifier value)|Modifier|false|false||median
null|Midline (qualifier value)|Modifier|false|false||mediannull|Statistical Median|LabModifier|false|false||median
null|Population Median|LabModifier|false|false||median
null|Sample Median|LabModifier|false|false||mediannull|Sternotomy (procedure)|Procedure|false|false||sternotomynull|Cardiac attachment|Finding|false|false||cardiacnull|Heart|Anatomy|false|false||cardiacnull|Cardiac - anatomy qualifier|Modifier|false|false||cardiacnull|Mediastinum|Anatomy|false|false||mediastinalnull|Mediastinal|Modifier|false|false||mediastinalnull|Hilar|Modifier|false|false||hilarnull|Contour form|Modifier|false|false||contoursnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Disease|Disorder|false|false||diseasenull|Increased (finding)|Finding|false|false||increased
null|Increase|Finding|false|false||increasednull|Increased|LabModifier|false|false||increasednull|Extent|Modifier|false|false||extent ofnull|Extent|Modifier|false|false||extentnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacity
null|Decreased translucency|Finding|false|false||opacitynull|Structure of base of right lung|Anatomy|false|false||right lung basenull|Right lung|Anatomy|false|false||right lungnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Basal segment of lung|Anatomy|false|false||lung basenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|nitrogenous base|Drug|false|false||base
null|Base|Drug|false|false||base
null|Dental Base|Drug|false|false||base
null|base - RoleClass|Drug|false|false||basenull|Base - General Qualifier|Finding|false|false||base
null|BPIFA4P gene|Finding|false|false||base
null|Base - RX Component Type|Finding|false|false||basenull|Anatomical base|Anatomy|false|false||basenull|Base - unit of product usage|LabModifier|false|false||basenull|Malaise|Finding|false|false||Illnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacities
null|Decreased translucency|Finding|false|false||opacitiesnull|Lingula of left lung|Anatomy|false|false||lingula
null|Lingula of cerebellum|Anatomy|false|false||lingula
null|Lingula|Anatomy|false|false||lingulanull|Lingula <Lingulidae>|Entity|false|false||lingulanull|Structure of left lower lobe of lung|Anatomy|false|false||left lower lobenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Similarity|Modifier|false|false||similarnull|null|Time|false|false||priornull|Small|LabModifier|false|false||Smallnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pleural effusion (disorder)|Finding|false|false||pleural effusion
null|Pleural effusion fluid|Finding|false|false||pleural effusion
null|null|Finding|false|false||pleural effusionnull|Pleural Diseases|Disorder|false|false||pleuralnull|Pleura|Anatomy|false|false||pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Hyperdistention|Disorder|false|false||hyperinflationnull|Lung|Anatomy|false|false||lungsnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|false|false||Evidence ofnull|Evidence|Finding|false|false||Evidencenull|Disease Progression|Finding|false|false||disease progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|true|false||progression
null|Progression|Finding|true|false||progressionnull|CAT scan of head|Procedure|false|false||CT Headnull|null|Attribute|false|false||CT Headnull|Problems with head|Disorder|false|false||Headnull|Procedure on head|Procedure|false|false||Headnull|Structure of head of caudate nucleus|Anatomy|false|false||Head
null|Head|Anatomy|false|false||Headnull|Head Device|Device|false|false||Headnull|findings aspects|Finding|false|false||FINDINGSnull|null|Attribute|false|false||FINDINGSnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Acute hemorrhage|Finding|true|false||acute hemorrhagenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Hemorrhage|Finding|true|false||hemorrhagenull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|Mass of body structure|Finding|true|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false||mass
null|null|Finding|true|false||mass
null|FBN1 wt Allele|Finding|true|false||mass
null|FBN1 gene|Finding|true|false||mass
null|Mass of body region|Finding|true|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Recent|Time|false|false||recentnull|Infarction|Finding|false|false||infarctionnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Encephalomalacia|Disorder|false|false||encephalomalacianull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|malignant neoplasm of frontal lobe|Disorder|false|false||frontal lobenull|frontal lobe|Anatomy|false|false||frontal lobenull|Coronal (qualifier value)|Modifier|false|false||frontalnull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Consistent with|Finding|false|false||compatible withnull|Compatible|Modifier|false|false||compatible withnull|Consistent with|Finding|false|false||compatiblenull|Compatible|Modifier|false|false||compatiblenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Infarction|Finding|false|false||infarctnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Heart Ventricle|Anatomy|false|false||ventriclesnull|Atrophic|Finding|false|false||atrophynull|bifrontal|Modifier|false|false||bifrontalnull|Areas <Spilosomini>|Entity|false|false||Areasnull|Area|Modifier|false|false||Areasnull|Periventricular|Modifier|false|false||periventricularnull|Subcortical|Anatomy|false|false||subcorticalnull|White matter|Anatomy|false|false||white matternull|White (population group)|Subject|false|false||white
null|Caucasian|Subject|false|false||white
null|Caucasians|Subject|false|false||whitenull|White color|Modifier|false|false||whitenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Sequela of disorder|Finding|false|false||sequelanull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Small|LabModifier|false|false||smallnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Ischemic|Finding|false|false||ischemicnull|Disease|Disorder|false|false||diseasenull|Bone Tissue, Human|Anatomy|true|false||osseous
null|Skeletal bone|Anatomy|true|false||osseousnull|Lesion|Finding|true|false||lesion
null|null|Finding|true|false||lesionnull|Pathologic calcification, calcified structure|Finding|false|false||calcifications
null|Physiologic calcification|Finding|false|false||calcificationsnull|Calcified (qualifier value)|Modifier|false|false||calcificationsnull|Bilateral|Modifier|false|false||bilateralnull|Carotid Arteries|Anatomy|false|false||carotidnull|Nasal sinus|Anatomy|false|false||paranasal sinusesnull|pathologic fistula|Disorder|false|false||sinusesnull|Head>Sinuses|Anatomy|false|false||sinuses
null|Nasal sinus|Anatomy|false|false||sinusesnull|null|Modifier|false|false||unremarkablenull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Intracranial Route of Administration|Finding|true|false||intracranialnull|Intracranial|Anatomy|true|false||intracranialnull|Process Pharmacologic Substance|Drug|true|false||processnull|Process (qualifier value)|Finding|true|false||processnull|bony process|Anatomy|true|false||processnull|Process|Phenomenon|true|false||processnull|Mass of body structure|Finding|true|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|true|false||mass
null|null|Finding|true|false||mass
null|FBN1 wt Allele|Finding|true|false||mass
null|FBN1 gene|Finding|true|false||mass
null|Mass of body region|Finding|true|false||massnull|Mass, a measure of quantity of matter|LabModifier|true|false||mass
null|Molecular Mass|LabModifier|true|false||massnull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Chest CT|Procedure|false|false||CT chestnull|null|Attribute|false|false||CT chestnull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|impression (attitude)|Finding|false|false||IMPRESSION
null|EKG impression|Finding|false|false||IMPRESSIONnull|Parameterized Data Type - Interval|Finding|false|false||Intervalnull|Interval|Time|false|false||Intervalnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Diffuse|Modifier|false|false||diffusenull|Bilateral|Modifier|false|false||bilateralnull|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glass
null|methamphetamine|Drug|false|false||glassnull|Chromosome 2q32-Q33 Deletion Syndrome|Disorder|false|false||glassnull|Glass Packaging Device|Device|false|false||glass
null|Glass (substance)|Device|false|false||glassnull|Abnormally opaque structure (morphologic abnormality)|Finding|false|false||opacities
null|Decreased translucency|Finding|false|false||opacitiesnull|Bronchioles|Anatomy|false|false||bronchiolarnull|Dense|Modifier|false|false||densenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Lingula of cerebellum|Anatomy|false|false||lingula
null|Lingula|Anatomy|false|false||lingula
null|Lingula of left lung|Anatomy|false|false||lingulanull|Lingula <Lingulidae>|Entity|false|false||lingulanull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of middle lobe of right lung|Anatomy|false|false||middle lobenull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Review of|Finding|false|false||review ofnull|Review (Publication Type)|Finding|false|false||review
null|Act Class - review|Finding|false|false||reviewnull|Numerous|LabModifier|false|false||multiplenull|Recent|Time|false|false||recentnull|null|Time|false|false||priornull|Chest problem|Finding|false|false||chestnull|Chest|Anatomy|false|false||chest
null|Anterior thoracic region|Anatomy|false|false||chestnull|X-rays, Homeopathic Preparations|Drug|false|false||x-raysnull|Plain x-ray|Procedure|false|false||x-rays
null|Diagnostic radiologic examination|Procedure|false|false||x-raysnull|Roentgen Rays|Phenomenon|false|false||x-raysnull|Cancer/Testis Antigen|Drug|false|false||CTsnull|Carpal Tunnel Syndrome|Disorder|false|false||CTsnull|TTR wt Allele|Finding|false|false||CTs
null|TTR gene|Finding|false|false||CTsnull|Concatenated Tag Sequencing|Procedure|false|false||CTsnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Patient Outcome - Worsening|Finding|false|false||worseningnull|Worsening (qualifier value)|Modifier|false|false||worseningnull|Bronchioloalveolar Adenocarcinoma|Disorder|true|false||bronchioalveolar carcinomanull|Carcinoma|Disorder|true|false||carcinomanull|Absent|Finding|true|false||absence ofnull|Absence (morphologic abnormality)|Disorder|true|false||absencenull|Absent|Finding|true|false||absencenull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|true|false||change
null|Changed status|LabModifier|true|false||changenull|Rapid|Modifier|true|false||rapidnull|Pneumonia|Disorder|true|false||pneumonianull|Course|Time|false|false||coursenull|Pneumonia|Disorder|false|false||pneumonianull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Unrecognized|Modifier|false|false||unrecognizednull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Basis|Drug|false|false||basisnull|Basis - conceptual entity|Finding|false|false||basisnull|Signs and Symptoms|Finding|false|false||clinical findingsnull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Patient Condition Code - Stable|Finding|false|false||Stablenull|Stable status|Modifier|false|false||Stablenull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Cardiomegaly|Finding|false|false||cardiomegalynull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Pulmonary Emphysema|Disorder|false|false||emphysemanull|Pathological accumulation of air in tissues|Finding|false|false||emphysemanull|Cholelithiasis|Disorder|true|false||Cholelithiasisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Cholecystitis|Disorder|true|false||cholecystitisnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|null|Disorder|false|false||NSCLCnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Hypoxia, CTCAE|Finding|false|false||hypoxia
null|Hypoxia|Finding|false|false||hypoxianull|Hypoxia, CTCAE|Finding|false|false||Hypoxia
null|Hypoxia|Finding|false|false||Hypoxianull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Complaint (finding)|Finding|false|false||complaintsnull|Progressive|Finding|false|false||progressivenull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Home oxygen supply|Finding|true|false||home oxygennull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|oxygen|Drug|true|false||oxygen
null|oxygen|Drug|true|false||oxygen
null|oxygen|Drug|true|false||oxygennull|Oxygen Therapy Care|Procedure|true|false||oxygennull|Oxygen Equipment Location|Modifier|true|false||oxygennull|Requirement|Finding|true|false||requirementnull|BaseLine dental cement|Drug|true|false||baselinenull|baseline - TableCellVerticalAlign|Finding|true|false||baselinenull|Baseline|LabModifier|true|false||baselinenull|On admission|Time|false|false||On admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|null|Device|false|false||NRBnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Saturated|Phenomenon|false|false||saturationsnull|Saturated|Phenomenon|false|false||saturationsnull|Admission activity|Procedure|true|false||Admission
null|Hospital admission|Procedure|true|false||Admissionnull|Plain chest X-ray|Procedure|true|false||CXRnull|Definite|Modifier|true|false||definite
null|Definitely Related to Intervention|Modifier|true|false||definitenull|Administration Method - Infiltrate|Finding|true|false||infiltrate
null|null|Finding|true|false||infiltrate
null|Infiltration|Finding|true|false||infiltratenull|Concern|Finding|false|false||concernnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Known|Modifier|false|false||knownnull|Lung diseases|Disorder|false|false||lung diseasenull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Disease|Disorder|false|false||diseasenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Leukocytes|Anatomy|false|false||WBCnull|Concern|Finding|false|false||concernnull|INFECTIOUS PROCESS|Finding|false|false||infectious processnull|Communicable Diseases|Disorder|false|false||infectiousnull|infectious - Entity Risk|Modifier|false|false||infectiousnull|Process Pharmacologic Substance|Drug|false|false||processnull|Process (qualifier value)|Finding|false|false||processnull|bony process|Anatomy|false|false||processnull|Process|Phenomenon|false|false||processnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|vancomycin|Drug|false|false||vancomycin
null|vancomycin|Drug|false|false||vancomycinnull|Vancomycin measurement|Procedure|false|false||vancomycinnull|Single Agent Therapy|Procedure|false|false||monotherapynull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|Late|Time|false|false||laternull|Plain chest X-ray|Procedure|false|false||CXRnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Additional|Finding|false|false||Additionalnull|Hypoxia, CTCAE|Finding|false|false||hypoxia
null|Hypoxia|Finding|false|false||hypoxianull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Biological Markers|Attribute|true|false||biomarkersnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Unable|Finding|false|false||unablenull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Due to|Finding|false|false||due
null|Due|Finding|false|false||duenull|Chronic Kidney Diseases|Disorder|false|false||chronic kidney diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Kidney Diseases|Disorder|false|false||kidney diseasenull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|Disease|Disorder|false|false||diseasenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Room Air|Drug|false|false||room airnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Endoglin, human|Drug|false|false||end
null|Endoglin, human|Drug|false|false||endnull|end - ActRelationshipCheckpoint|Finding|false|false||end
null|ENG gene|Finding|false|false||end
null|ENG wt Allele|Finding|false|false||endnull|Stop (qualifier value)|Time|false|false||endnull|End|Modifier|false|false||endnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|exercise induced|Finding|false|false||exertionalnull|Hypoxia, CTCAE|Finding|false|false||hypoxia
null|Hypoxia|Finding|false|false||hypoxianull|Usually asymptomatic|Finding|false|false||usually asymptomaticnull|Usually|Finding|false|false||usuallynull|Usual|Modifier|false|false||usuallynull|Asymptomatic diagnosis of|Finding|false|false||asymptomatic
null|Asymptomatic (finding)|Finding|false|false||asymptomaticnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Pneumonia|Disorder|false|false||pneumonianull|Lung consolidation|Disorder|false|false||Consolidationnull|Consolidation|Modifier|false|false||Consolidationnull|Structure of left lower lobe of lung|Anatomy|false|false||left lower lobenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Structure of lower lobe of lung|Anatomy|false|false||lower lobenull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|AKT1S1 wt Allele|Finding|false|false||lobe
null|AKT1S1 gene|Finding|false|false||lobenull|lobe|Anatomy|false|false||lobenull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Disease|Disorder|false|false||diseasenull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Time course|Time|false|false||time coursenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Course|Time|false|false||coursenull|Administration Method - Infiltrate|Finding|false|false||infiltrate
null|null|Finding|false|false||infiltrate
null|Infiltration|Finding|false|false||infiltratenull|Growth and Development function|Finding|false|false||development
null|development aspects|Finding|false|false||development
null|biological development|Finding|false|false||development
null|Development|Finding|false|false||developmentnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Procedure Practitioner Identifier Code Type - Radiologist|Finding|false|false||radiologistnull|radiologist|Subject|false|false||radiologistnull|Opposite|Modifier|false|false||oppositenull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|null|Disorder|false|false||NSCLCnull|Pneumonia|Disorder|true|false||pneumonianull|Course|Time|false|false||coursenull|ceftriaxone|Drug|false|false||ceftriaxone
null|ceftriaxone|Drug|false|false||ceftriaxonenull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Living Alone|Finding|false|false||alonenull|alone - group size|Subject|false|false||alonenull|Singular|LabModifier|false|false||alonenull|Blood culture|Procedure|true|false||Blood culturesnull|Blood and lymphatic system disorders|Disorder|true|false||Bloodnull|peripheral blood|Finding|true|false||Blood
null|Blood|Finding|true|false||Blood
null|In Blood|Finding|true|false||Bloodnull|Culture (Anthropological)|Finding|true|false||culturesnull|Growth & development aspects|Finding|true|false||growth
null|Tissue Growth|Finding|true|false||growth
null|Growth|Finding|true|false||growth
null|growth aspects|Finding|true|false||growthnull|Growth action|Phenomenon|true|false||growthnull|Numerous|LabModifier|false|false||Multiplenull|Specimen Type - Sputum|Finding|false|false||sputum
null|null|Finding|false|false||sputum
null|Sputum|Finding|false|false||sputumnull|Culture (Anthropological)|Finding|false|false||culturesnull|Oral Microbiome|Entity|false|false||oral flora
null|oral bacteria|Entity|false|false||oral floranull|Oral Dosage Form|Drug|false|false||oralnull|Oral Route of Administration|Finding|false|false||oral
null|Oral (intended site)|Finding|false|false||oralnull|Oral cavity|Anatomy|false|false||oralnull|Oral|Modifier|false|false||oralnull|Portion of urine|Finding|true|false||Urine
null|null|Finding|true|false||Urine
null|Urine|Finding|true|false||Urine
null|In Urine|Finding|true|false||Urine
null|Urine specimen|Finding|true|false||Urinenull|Legionella|Entity|false|false||legionellanull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Course|Time|false|false||coursenull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|null|Disorder|false|false||NSCLCnull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Current (present time)|Time|true|false||currentlynull|pharmacotherapeutic|Finding|true|false||chemotherapynull|Chemotherapy Regimen|Procedure|true|false||chemotherapy
null|Pharmacotherapy|Procedure|true|false||chemotherapy
null|Chemotherapy|Procedure|true|false||chemotherapynull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|Oncologists|Subject|false|false||oncologistnull|Continuous|Finding|false|false||continuednull|surveillance aspects|Finding|false|false||surveillancenull|Medical Surveillance|Procedure|false|false||surveillancenull|legal surveillance|Event|false|false||surveillancenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Further|Modifier|false|false||furthernull|Palliative care service|Entity|false|false||palliativenull|Palliative|Modifier|false|false||palliativenull|Systemic Route of Administration|Finding|false|false||systemic
null|Systemic|Finding|false|false||systemicnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Symptomatic|Finding|false|false||symptomaticnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Glycogen Storage Disease Type VI|Disorder|false|false||her diseasenull|Disease|Disorder|false|false||diseasenull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Disease Progression|Finding|false|false||disease progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Further|Modifier|false|false||furthernull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Risk|Finding|false|false||risksnull|Benefit|LabModifier|false|false||benefitsnull|Additional|Finding|false|false||additionalnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Abnormal renal function|Finding|false|false||kidney dysfunctionnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Comorbidity|Finding|false|false||comorbiditiesnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Further|Modifier|false|false||furthernull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Disease Progression|Finding|false|false||disease progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Relationship modifier - Patient|Finding|true|false||Patient
null|Specimen Type - Patient|Finding|true|false||Patient
null|Mail Claim Party - Patient|Finding|true|false||Patient
null|Report source - Patient|Finding|true|false||Patient
null|null|Finding|true|false||Patient
null|Disabled Person Code - Patient|Finding|true|false||Patientnull|Patients|Subject|true|false||Patientnull|Veterinary Patient|Entity|true|false||Patientnull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Electrocardiogram image|Finding|false|false||EKG
null|Electrocardiogram|Finding|false|false||EKGnull|Electrocardiography|Procedure|false|false||EKGnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Mental Depression|Disorder|false|false||depressionsnull|Biological Markers|Attribute|false|false||Biomarkersnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Adrenergic beta-Antagonists|Drug|false|false||beta-blockernull|Greek letter beta|Finding|false|false||betanull|Beta <eudicots>|Entity|false|false||betanull|Beta Distribution|LabModifier|false|false||betanull|Decreasing|Finding|false|false||decreased
null|Reduced|Finding|false|false||decreasednull|Decreased|LabModifier|false|false||decreasednull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Living Arrangement - Relative|Finding|false|false||relativenull|null|Attribute|false|false||relativenull|Relative (related person)|Subject|false|false||relativenull|Relative|Modifier|false|false||relativenull|Hypotension|Finding|false|false||hypotensionnull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Plavix|Drug|false|false||plavix
null|Plavix|Drug|false|false||plavixnull|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statin
null|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Drug|false|false||statinnull|EEF1A2 gene|Finding|false|false||statinnull|3-hydroxy-3-methylglutaryl-coenzyme A reductase inhibitor (disposition)|Modifier|false|false||statinnull|Chronic systolic heart failure|Disorder|false|false||chronic systolic CHFnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|systolic congestive heart failure|Disorder|false|false||systolic CHFnull|Systole|Finding|false|false||systolicnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|LVEF (procedure)|Procedure|false|false||LVEFnull|Left ventricular ejection fraction|Attribute|false|false||LVEFnull|Transthoracic echocardiography|Procedure|false|false||TTEnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Living Arrangement - Relative|Finding|false|false||relativenull|null|Attribute|false|false||relativenull|Relative (related person)|Subject|false|false||relativenull|Relative|Modifier|false|false||relativenull|Hypotension|Finding|false|false||hypotensionnull|Exertional tachycardia|Finding|false|false||exertional tachycardianull|exercise induced|Finding|false|false||exertionalnull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|creatinine|Drug|false|false||Creatinine
null|creatinine|Drug|false|false||Creatininenull|Creatinine metabolic function|Finding|false|false||Creatininenull|Creatinine measurement|Procedure|false|false||Creatininenull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Inventory of Callous-Unemotional Traits|Finding|false|false||ICUnull|Structure of intraculminate fissure|Anatomy|false|false||ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|monitoring of urine output for fluid balance|Procedure|false|false||urine outputnull|null|Attribute|false|false||urine output
null|null|Attribute|false|false||urine outputnull|Urine volume finding|LabModifier|false|false||urine outputnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Microcytic anemia|Disorder|false|false||Microcytic anemianull|microcytic|Finding|false|false||Microcyticnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Presentation|Finding|false|false||presentationnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Hemorrhage|Finding|true|false||bleedingnull|Exam|Finding|true|false||examnull|Medical Examination|Procedure|true|false||examnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Appropriate|Modifier|false|false||appropriatenull|Elevation procedure|Procedure|false|false||elevationnull|Elevation|Modifier|false|false||elevationnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|Steady|Modifier|false|false||steadynull|Course|Time|false|false||coursenull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|guaiac|Drug|false|false||guaiac
null|guaiac|Drug|false|false||guaiacnull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Further|Modifier|false|false||furthernull|Work-up|Procedure|false|false||work-upnull|Work|Event|false|false||worknull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|most likely|Finding|false|false||most likelynull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Secondary to|Modifier|false|false||secondary tonull|Neoplasm Metastasis|Disorder|false|false||secondarynull|metastatic qualifier|Finding|false|false||secondarynull|Secondary to|Modifier|false|false||secondarynull|second (number)|LabModifier|false|false||secondarynull|Acute inflammation|Finding|false|false||acute inflammationnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Inflammation|Finding|false|false||inflammationnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Underlying|Finding|false|false||underlyingnull|Chronic disease|Disorder|false|false||chronic diseasenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Disease|Disorder|false|false||diseasenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|amlodipine|Drug|false|false||amlodipine
null|amlodipine|Drug|false|false||amlodipinenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one dailynull|Daily|Time|false|false||dailynull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Lipitor|Drug|false|false||Lipitor
null|Lipitor|Drug|false|false||Lipitornull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Calcitriol Drug Class|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|Calcitriol Drug Class|Drug|false|false||calcitriolnull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once A Day|Drug|false|false||once a daynull|Once daily|Time|false|false||once a daynull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|Plavix|Drug|false|false||Plavix
null|Plavix|Drug|false|false||Plavixnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acidnull|Folic acid measurement|Procedure|false|false||folic acidnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one dailynull|Daily|Time|false|false||dailynull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|loperamide|Drug|false|false||loperamide
null|loperamide|Drug|false|false||loperamidenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Twice a day|Time|false|false||twice dailynull|Daily|Time|false|false||dailynull|lorazepam|Drug|false|false||lorazepam
null|lorazepam|Drug|false|false||lorazepamnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Hour|Time|false|false||hoursnull|Nausea|Finding|false|false||Nauseanull|null|Attribute|false|false||Nauseanull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Lopressor|Drug|false|false||Lopressor
null|Lopressor|Drug|false|false||Lopressornull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|trazodone|Drug|false|false||trazodone
null|trazodone|Drug|false|false||trazodonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one dailynull|Daily|Time|false|false||dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one dailynull|Daily|Time|false|false||dailynull|ranitidine hydrochloride|Drug|false|false||ranitidine HCl
null|ranitidine hydrochloride|Drug|false|false||ranitidine HClnull|ranitidine|Drug|false|false||ranitidine
null|ranitidine|Drug|false|false||ranitidinenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Acid Control|Drug|false|false||Acid Control
null|Acid Control|Drug|false|false||Acid Controlnull|Control brand of phenylpropanolamine|Drug|false|false||Control
null|CONTROL veterinary product|Drug|false|false||Control
null|control substance|Drug|false|false||Control
null|Control brand of phenylpropanolamine|Drug|false|false||Controlnull|Control - Relationship modifier|Finding|false|false||Control
null|Control function|Finding|false|false||Control
null|Scientific Control|Finding|false|false||Controlnull|Control Groups|Subject|false|false||Controlnull|True Control Status|Modifier|false|false||Control
null|control aspects|Modifier|false|false||Controlnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one daily
null|One Daily|Drug|false|false||one dailynull|Daily|Time|false|false||dailynull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Continuous|Finding|false|false||continuousnull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|portability|Modifier|false|false||portabilitynull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|levofloxacin|Drug|false|false||levofloxacin
null|levofloxacin|Drug|false|false||levofloxacinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Every - dosing instruction fragment|Finding|false|false||everynull|Every (qualifier)|Modifier|false|false||everynull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Last|Modifier|false|false||lastnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|atorvastatin|Drug|false|false||atorvastatin
null|atorvastatin|Drug|false|false||atorvastatinnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|metoprolol tartrate|Drug|false|false||metoprolol tartrate
null|metoprolol tartrate|Drug|false|false||metoprolol tartratenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|tartrate|Drug|false|false||tartrate
null|Tartrates|Drug|false|false||tartrate
null|tartrate|Drug|false|false||tartratenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Changing|Finding|false|false||CHANGEnull|Change - procedure|Procedure|false|false||CHANGEnull|Delta (difference)|LabModifier|false|false||CHANGE
null|Changed status|LabModifier|false|false||CHANGEnull|Act Relationship Subset - previous|Time|false|false||PREVIOUS
null|Previous|Time|false|false||PREVIOUSnull|Evening|Time|false|false||EVENINGnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Hold - dosing instruction fragment|Finding|false|false||hold
null|hold - Data Operation|Finding|false|false||holdnull|Hold (action)|Event|false|false||holdnull|Loose stool|Finding|false|false||loose stools
null|Diarrhea|Finding|false|false||loose stoolsnull|Loose|Modifier|false|false||loosenull|Feces|Finding|false|false||stoolsnull|null|Attribute|false|false||stoolsnull|Stool seat|Device|false|false||stoolsnull|trazodone|Drug|false|false||trazodone
null|trazodone|Drug|false|false||trazodonenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Once a day, at bedtime|Time|false|false||at bedtimenull|Once a day, at bedtime|Time|false|false||bedtime
null|Bedtime (qualifier value)|Time|false|false||bedtimenull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|clopidogrel|Drug|false|false||clopidogrel
null|clopidogrel|Drug|false|false||clopidogrelnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|ranitidine hydrochloride|Drug|false|false||ranitidine HCl
null|ranitidine hydrochloride|Drug|false|false||ranitidine HClnull|ranitidine|Drug|false|false||ranitidine
null|ranitidine|Drug|false|false||ranitidinenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Calcitriol Drug Class|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|calcitriol|Drug|false|false||calcitriol
null|Calcitriol Drug Class|Drug|false|false||calcitriolnull|microgram|LabModifier|false|false||mcgnull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|capsule (pharmacologic)|Drug|false|false||Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false||Capsule
null|Structure of organ capsule|Anatomy|false|false||Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acid
null|folic acid|Drug|false|false||folic acidnull|Folic acid measurement|Procedure|false|false||folic acidnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|aspirin|Drug|false|false||aspirin
null|aspirin|Drug|false|false||aspirinnull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Receptors, Antigen, B-Cell|Drug|false|false||Sig
null|Receptors, Antigen, B-Cell|Drug|false|false||Signull|Receptors, Antigen, B-Cell|Finding|false|false||Signull|Short insular gyrus|Anatomy|false|false||Signull|Surveillance Implementation Group|Entity|false|false||Sig
null|Staphylococcus intermedius group|Entity|false|false||Signull|Chewable Tablet|Drug|false|false||Tablet, Chewablenull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|Daily|Time|false|false||DAILYnull|Daily|Time|false|false||Dailynull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Pneumonia|Disorder|false|false||pneumonianull|stage, small cell lung cancer|Disorder|false|false||small cell lung cancer stagenull|Small cell carcinoma of lung|Disorder|false|false||small cell lung cancernull|Small|LabModifier|false|false||smallnull|CELP gene|Finding|false|false||cell
null|CEL gene|Finding|false|false||cellnull|Cells|Anatomy|false|false||cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Stage IV Lung Cancer AJCC v7|Disorder|false|false||lung cancer stage IVnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Diagnostic Neoplasm Staging|Procedure|false|false||cancer stagenull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Stage level 4|Finding|false|false||stage IVnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Progressive|Finding|false|false||progressingnull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis|Procedure|false|false||DIAGNOSESnull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Acute inflammation|Finding|false|false||acute inflammationnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Inflammation|Finding|false|false||inflammationnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Chronic systolic heart failure|Disorder|false|false||chronic systolic CHFnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|systolic congestive heart failure|Disorder|false|false||systolic CHFnull|Systole|Finding|false|false||systolicnull|Congestive heart failure|Disorder|false|false||CHFnull|Choroidal fissure|Anatomy|false|false||CHFnull|Hypertensive disease|Disorder|false|false||HTNnull|Chronic Kidney Diseases|Disorder|false|false||CKDnull|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Levels (qualifier value)|Modifier|false|false||levelsnull|Room type - Intensive care unit|Finding|false|false||Intensive Care Unitnull|intensive care unit|Device|false|false||Intensive Care Unitnull|intensive care unit|Entity|false|false||Intensive Care Unitnull|intensive care|Procedure|false|false||Intensive Carenull|Specialty Type - Intensive care|Title|false|false||Intensive Carenull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Malignant neoplasm of lung|Disorder|false|false||lung cancer
null|Carcinoma of lung|Disorder|false|false||lung cancernull|Lung diseases|Disorder|false|false||lungnull|Lung Problem|Finding|false|false||lungnull|Chest>Lung|Anatomy|false|false||lung
null|Lung|Anatomy|false|false||lungnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Probable diagnosis|Finding|false|false||probablenull|Probability|LabModifier|false|false||probablenull|Pneumonia|Disorder|false|false||pneumonianull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygen
null|oxygen|Drug|false|false||oxygennull|Oxygen Therapy Care|Procedure|false|false||oxygennull|Oxygen Equipment Location|Modifier|false|false||oxygennull|Levels (qualifier value)|Modifier|false|false||levelsnull|Primary Oncologist|Subject|false|false||primary oncologistnull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|Oncologists|Subject|false|false||oncologistnull|Risks and Benefits|Modifier|false|false||risks and benefitsnull|Risk|Finding|false|false||risksnull|Benefit|LabModifier|false|false||benefitsnull|Additional|Finding|false|false||additionalnull|pharmacotherapeutic|Finding|false|false||chemotherapynull|Chemotherapy Regimen|Procedure|false|false||chemotherapy
null|Pharmacotherapy|Procedure|false|false||chemotherapy
null|Chemotherapy|Procedure|false|false||chemotherapynull|Abnormal renal function|Finding|false|false||kidney dysfunctionnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||kidney
null|Benign neoplasm of kidney|Disorder|false|false||kidneynull|Kidney problem|Finding|false|false||kidneynull|examination of kidney|Procedure|false|false||kidney
null|Procedures on Kidney|Procedure|false|false||kidneynull|Kidney|Anatomy|false|false||kidney
null|Both kidneys|Anatomy|false|false||kidneynull|DYSFUNCTION - SKIN DISORDERS|Disorder|false|false||dysfunctionnull|Dysfunction|Finding|false|false||dysfunction
null|physiopathological|Finding|false|false||dysfunction
null|Functional disorder|Finding|false|false||dysfunctionnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Problems - What subject filter|Finding|false|false||problemsnull|X-Ray Computed Tomography|Procedure|false|false||CT scannull|Radionuclide Imaging|Procedure|false|false||scan
null|Scanning|Procedure|false|false||scannull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Further|Modifier|false|false||furthernull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Disease Progression|Finding|false|false||disease progressionnull|Disease|Disorder|false|false||diseasenull|Disease Progression|Finding|false|false||progression
null|Progression|Finding|false|false||progressionnull|Congestive heart failure|Disorder|false|false||congestive heart failurenull|Congestive|Modifier|false|false||congestivenull|Congestive heart failure|Disorder|false|false||heart failure
null|Heart failure|Disorder|false|false||heart failurenull|Malignant neoplasm of heart|Disorder|false|false||heart
null|benign neoplasm of heart|Disorder|false|false||heartnull|HEART PROBLEM|Finding|false|false||heartnull|Chest>Heart|Anatomy|false|false||heart
null|Heart|Anatomy|false|false||heartnull|Failure (biologic function)|Finding|false|false||failure
null|Failure|Finding|false|false||failure
null|Personal failure|Finding|false|false||failurenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Lasix|Drug|false|false||lasix
null|Lasix|Drug|false|false||lasixnull|amlodipine|Drug|false|false||amlodipine
null|amlodipine|Drug|false|false||amlodipinenull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Evening|Time|false|false||eveningnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Usual|Modifier|false|false||usualnull|Every morning|Time|false|false||every morningnull|Morning|Time|false|false||morningnull|Call - dosing instruction fragment|Finding|false|false||call
null|Call (Instruction)|Finding|false|false||call
null|Decision|Finding|false|false||call
null|CHL1 gene|Finding|false|false||callnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions