 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
F|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
NEUROSURGERY|158,170
<EOL>|170,171
<EOL>|172,173
Allergies|173,182
:|182,183
<EOL>|184,185
No|185,187
Known|188,193
Allergies|194,203
/|204,205
Adverse|206,213
Drug|214,218
Reactions|219,228
<EOL>|228,229
<EOL>|230,231
Attending|231,240
:|240,241
_|242,243
_|243,244
_|244,245
.|245,246
<EOL>|246,247
<EOL>|248,249
Chief|249,254
Complaint|255,264
:|264,265
<EOL>|265,266
Headaches|266,275
<EOL>|275,276
<EOL>|277,278
Major|278,283
Surgical|284,292
or|293,295
Invasive|296,304
Procedure|305,314
:|314,315
<EOL>|315,316
_|316,317
_|317,318
_|318,319
-|320,321
Suboccipital|322,334
craniotomy|335,345
for|346,349
resection|350,359
of|360,362
cerebellar|363,373
<EOL>|374,375
lesion|375,381
<EOL>|381,382
<EOL>|382,383
<EOL>|384,385
History|385,392
of|393,395
Present|396,403
Illness|404,411
:|411,412
<EOL>|412,413
_|413,414
_|414,415
_|415,416
is|417,419
a|420,421
_|422,423
_|423,424
_|424,425
female|426,432
with|433,437
hx|438,440
cerebral|441,449
aneurysm|450,458
<EOL>|459,460
clipping|460,468
in|469,471
_|472,473
_|473,474
_|474,475
who|476,479
presents|480,488
from|489,493
OSH|494,497
with|498,502
left|503,507
cerebellar|508,518
<EOL>|519,520
hypodensity|520,531
concerning|532,542
for|543,546
underlying|547,557
lesion|558,564
.|564,565
Patient|566,573
reports|574,581
<EOL>|582,583
that|583,587
three|588,593
weeks|594,599
ago|600,603
she|604,607
started|608,615
having|616,622
headaches|623,632
,|632,633
which|634,639
is|640,642
<EOL>|643,644
abnormal|644,652
for|653,656
her|657,660
.|660,661
She|662,665
describes|666,675
the|676,679
headaches|680,689
to|690,692
be|693,695
global|696,702
and|703,706
<EOL>|707,708
resolve|708,715
with|716,720
Tylenol|721,728
,|728,729
but|730,733
at|734,736
the|737,740
worst|741,746
was|747,750
an|751,753
_|754,755
_|755,756
_|756,757
.|757,758
She|759,762
also|763,767
<EOL>|768,769
reports|769,776
having|777,783
difficulty|784,794
walking|795,802
,|802,803
which|804,809
also|810,814
started|815,822
about|823,828
<EOL>|829,830
three|830,835
weeks|836,841
ago|842,845
.|845,846
She|847,850
describes|851,860
her|861,864
walking|865,872
as|873,875
"|876,877
staggering|877,887
side|888,892
<EOL>|893,894
to|894,896
side|897,901
.|901,902
"|902,903
She|904,907
denies|908,914
any|915,918
vision|919,925
changes|926,933
,|933,934
nausea|935,941
,|941,942
vomiting|943,951
,|951,952
<EOL>|953,954
confusion|954,963
,|963,964
or|965,967
word|968,972
finding|973,980
difficulty|981,991
.|991,992
She|993,996
saw|997,1000
her|1001,1004
eye|1005,1008
doctor|1009,1015
<EOL>|1016,1017
this|1017,1021
morning|1022,1029
for|1030,1033
routine|1034,1041
visit|1042,1047
,|1047,1048
who|1049,1052
referred|1053,1061
her|1062,1065
to|1066,1068
the|1069,1072
ED|1073,1075
for|1076,1079
<EOL>|1080,1081
evaluation|1081,1091
of|1092,1094
these|1095,1100
symptoms|1101,1109
.|1109,1110
OSH|1111,1114
CT|1115,1117
showed|1118,1124
an|1125,1127
area|1128,1132
of|1133,1135
<EOL>|1136,1137
hypodensity|1137,1148
in|1149,1151
the|1152,1155
left|1156,1160
cerebellum|1161,1171
,|1171,1172
concerning|1173,1183
for|1184,1187
underlying|1188,1198
<EOL>|1199,1200
lesion|1200,1206
.|1206,1207
She|1208,1211
was|1212,1215
subsequently|1216,1228
transferred|1229,1240
to|1241,1243
_|1244,1245
_|1245,1246
_|1246,1247
.|1247,1248
<EOL>|1249,1250
<EOL>|1250,1251
Of|1251,1253
note|1254,1258
,|1258,1259
patient|1260,1267
reports|1268,1275
her|1276,1279
aneurysm|1280,1288
clip|1289,1293
is|1294,1296
not|1297,1300
MRI|1301,1304
<EOL>|1305,1306
compatible|1306,1316
.|1316,1317
<EOL>|1317,1318
<EOL>|1318,1319
<EOL>|1320,1321
Past|1321,1325
Medical|1326,1333
History|1334,1341
:|1341,1342
<EOL>|1342,1343
-|1343,1344
_|1345,1346
_|1346,1347
_|1347,1348
<EOL>|1349,1350
-|1350,1351
Hypertension|1352,1364
<EOL>|1365,1366
-|1366,1367
S|1368,1369
/|1369,1370
p|1370,1371
aneurysm|1372,1380
clipping|1381,1389
_|1390,1391
_|1391,1392
_|1392,1393
at|1394,1396
_|1397,1398
_|1398,1399
_|1399,1400
by|1401,1403
Dr.|1404,1407
_|1408,1409
_|1409,1410
_|1410,1411
<EOL>|1411,1412
<EOL>|1413,1414
Social|1414,1420
History|1421,1428
:|1428,1429
<EOL>|1429,1430
_|1430,1431
_|1431,1432
_|1432,1433
<EOL>|1433,1434
Family|1434,1440
History|1441,1448
:|1448,1449
<EOL>|1449,1450
No|1450,1452
known|1453,1458
history|1459,1466
of|1467,1469
stroke|1470,1476
,|1476,1477
cancer|1478,1484
,|1484,1485
aneurysm|1486,1494
.|1494,1495
<EOL>|1496,1497
<EOL>|1497,1498
<EOL>|1499,1500
Physical|1500,1508
Exam|1509,1513
:|1513,1514
<EOL>|1514,1515
ON|1515,1517
ADMISSION|1518,1527
:|1527,1528
<EOL>|1529,1530
O|1530,1531
:|1531,1532
T|1533,1534
:|1534,1535
97.9|1536,1540
BP|1542,1544
:|1544,1545
130|1546,1549
/|1549,1550
62|1550,1552
HR|1555,1557
:|1557,1558
64|1559,1561
R|1565,1566
16|1567,1569
O2Sats|1574,1580
98|1581,1583
%|1583,1584
RA|1585,1587
<EOL>|1587,1588
Gen|1588,1591
:|1591,1592
WD|1593,1595
/|1595,1596
WN|1596,1598
,|1598,1599
comfortable|1600,1611
,|1611,1612
NAD|1613,1616
.|1616,1617
<EOL>|1617,1618
HEENT|1618,1623
:|1623,1624
Pupils|1625,1631
:|1631,1632
L|1633,1634
_|1635,1636
_|1636,1637
_|1637,1638
,|1638,1639
R|1640,1641
_|1642,1643
_|1643,1644
_|1644,1645
EOMs|1653,1657
full|1658,1662
<EOL>|1662,1663
Neck|1663,1667
:|1667,1668
Supple|1669,1675
.|1675,1676
<EOL>|1676,1677
Extrem|1677,1683
:|1683,1684
Warm|1685,1689
and|1690,1693
well|1694,1698
-|1698,1699
perfused|1699,1707
.|1707,1708
<EOL>|1708,1709
<EOL>|1709,1710
Neuro|1710,1715
:|1715,1716
<EOL>|1716,1717
Mental|1717,1723
status|1724,1730
:|1730,1731
Awake|1732,1737
and|1738,1741
alert|1742,1747
,|1747,1748
cooperative|1749,1760
with|1761,1765
exam|1766,1770
,|1770,1771
normal|1772,1778
<EOL>|1778,1779
affect|1779,1785
.|1785,1786
<EOL>|1786,1787
Orientation|1787,1798
:|1798,1799
Oriented|1800,1808
to|1809,1811
person|1812,1818
,|1818,1819
place|1820,1825
,|1825,1826
and|1827,1830
date|1831,1835
.|1835,1836
<EOL>|1836,1837
Language|1837,1845
:|1845,1846
Speech|1847,1853
fluent|1854,1860
with|1861,1865
good|1866,1870
comprehension|1871,1884
and|1885,1888
repetition|1889,1899
.|1899,1900
<EOL>|1900,1901
Naming|1901,1907
intact|1908,1914
.|1914,1915
No|1916,1918
dysarthria|1919,1929
or|1930,1932
paraphasic|1933,1943
errors|1944,1950
.|1950,1951
<EOL>|1951,1952
<EOL>|1952,1953
Cranial|1953,1960
Nerves|1961,1967
:|1967,1968
<EOL>|1968,1969
I|1969,1970
:|1970,1971
Not|1972,1975
tested|1976,1982
<EOL>|1982,1983
II|1983,1985
:|1985,1986
Left|1987,1991
pupil|1992,1997
5|1998,1999
-|1999,2000
4mm|2000,2003
,|2003,2004
right|2005,2010
4|2011,2012
-|2012,2013
3mm|2013,2016
,|2016,2017
both|2018,2022
equally|2023,2030
reactive|2031,2039
to|2040,2042
<EOL>|2042,2043
light|2043,2048
.|2048,2049
<EOL>|2050,2051
III|2051,2054
,|2054,2055
IV|2056,2058
,|2058,2059
VI|2060,2062
:|2062,2063
Extraocular|2064,2075
movements|2076,2085
intact|2086,2092
bilaterally|2093,2104
without|2105,2112
<EOL>|2112,2113
nystagmus|2113,2122
.|2122,2123
<EOL>|2123,2124
V|2124,2125
,|2125,2126
VII|2127,2130
:|2130,2131
Facial|2132,2138
strength|2139,2147
and|2148,2151
sensation|2152,2161
intact|2162,2168
and|2169,2172
symmetric|2173,2182
.|2182,2183
<EOL>|2183,2184
XI|2184,2186
:|2186,2187
Sternocleidomastoid|2188,2207
and|2208,2211
trapezius|2212,2221
normal|2222,2228
bilaterally|2229,2240
.|2240,2241
<EOL>|2241,2242
XII|2242,2245
:|2245,2246
Tongue|2247,2253
midline|2254,2261
without|2262,2269
fasciculations|2270,2284
.|2284,2285
<EOL>|2285,2286
<EOL>|2286,2287
Motor|2287,2292
:|2292,2293
Normal|2294,2300
bulk|2301,2305
and|2306,2309
tone|2310,2314
bilaterally|2315,2326
.|2326,2327
No|2328,2330
abnormal|2331,2339
movements|2340,2349
,|2349,2350
<EOL>|2350,2351
tremors|2351,2358
.|2358,2359
Strength|2360,2368
full|2369,2373
power|2374,2379
_|2380,2381
_|2381,2382
_|2382,2383
throughout|2384,2394
.|2394,2395
Slight|2396,2402
left|2403,2407
upward|2408,2414
<EOL>|2415,2416
drift|2416,2421
<EOL>|2421,2422
<EOL>|2422,2423
Sensation|2423,2432
:|2432,2433
Intact|2434,2440
to|2441,2443
light|2444,2449
touch|2450,2455
<EOL>|2455,2456
<EOL>|2456,2457
Coordination|2457,2469
:|2469,2470
normal|2471,2477
on|2478,2480
finger|2481,2487
-|2487,2488
nose|2488,2492
-|2492,2493
finger|2493,2499
and|2500,2503
heel|2504,2508
to|2509,2511
shin|2512,2516
<EOL>|2516,2517
<EOL>|2517,2518
=|2518,2519
=|2519,2520
=|2520,2521
=|2521,2522
=|2522,2523
=|2523,2524
=|2524,2525
=|2525,2526
=|2526,2527
=|2527,2528
=|2528,2529
=|2529,2530
=|2530,2531
=|2531,2532
=|2532,2533
=|2533,2534
=|2534,2535
=|2535,2536
=|2536,2537
=|2537,2538
=|2538,2539
=|2539,2540
=|2540,2541
=|2541,2542
=|2542,2543
=|2543,2544
=|2544,2545
=|2545,2546
=|2546,2547
=|2547,2548
=|2548,2549
=|2549,2550
=|2550,2551
=|2551,2552
=|2552,2553
=|2553,2554
=|2554,2555
=|2555,2556
=|2556,2557
=|2557,2558
=|2558,2559
=|2559,2560
=|2560,2561
=|2561,2562
=|2562,2563
=|2563,2564
=|2564,2565
=|2565,2566
=|2566,2567
=|2567,2568
=|2568,2569
=|2569,2570
=|2570,2571
=|2571,2572
<EOL>|2572,2573
<EOL>|2573,2574
ON|2574,2576
DISCHARGE|2577,2586
:|2586,2587
<EOL>|2588,2589
Exam|2589,2593
:|2593,2594
<EOL>|2594,2595
<EOL>|2595,2596
Opens|2596,2601
eyes|2602,2606
:|2606,2607
[|2608,2609
x|2609,2610
]|2610,2611
Spontaneous|2611,2622
[|2623,2624
]|2625,2626
To|2626,2628
voice|2629,2634
[|2635,2636
]|2637,2638
To|2638,2640
noxious|2641,2648
<EOL>|2648,2649
<EOL>|2649,2650
Orientation|2650,2661
:|2661,2662
[|2663,2664
x|2664,2665
]|2665,2666
Person|2666,2672
[|2673,2674
x|2674,2675
]|2675,2676
Place|2676,2681
[|2682,2683
x|2683,2684
]|2684,2685
Time|2685,2689
<EOL>|2689,2690
<EOL>|2690,2691
Follows|2691,2698
commands|2699,2707
:|2707,2708
[|2709,2710
]|2711,2712
Simple|2712,2718
[|2719,2720
x|2720,2721
]|2721,2722
Complex|2722,2729
[|2730,2731
]|2732,2733
None|2733,2737
<EOL>|2737,2738
<EOL>|2738,2739
Pupils|2739,2745
:|2745,2746
Right|2748,2753
4|2755,2756
-|2756,2757
3mm|2757,2760
Left|2766,2770
5|2771,2772
-|2772,2773
4mm|2773,2776
-|2777,2778
chronic|2779,2786
<EOL>|2786,2787
<EOL>|2787,2788
EOM|2788,2791
:|2791,2792
[|2793,2794
]|2795,2796
Full|2796,2800
[|2801,2802
x|2802,2803
]|2803,2804
Restricted|2804,2814
-|2815,2816
chronic|2817,2824
,|2824,2825
most|2826,2830
prominent|2831,2840
left|2841,2845
<EOL>|2846,2847
lateral|2847,2854
<EOL>|2854,2855
<EOL>|2855,2856
Face|2856,2860
Symmetric|2861,2870
:|2870,2871
[|2872,2873
x|2873,2874
]|2874,2875
Yes|2875,2878
[|2879,2880
]|2881,2882
NoTongue|2882,2890
Midline|2891,2898
:|2898,2899
[|2900,2901
x|2901,2902
]|2902,2903
Yes|2903,2906
[|2907,2908
]|2909,2910
No|2910,2912
<EOL>|2912,2913
<EOL>|2913,2914
Pronator|2914,2922
Drift|2923,2928
:|2928,2929
[|2930,2931
]|2932,2933
Yes|2933,2936
[|2937,2938
x|2938,2939
]|2939,2940
No|2940,2942
Speech|2946,2952
Fluent|2953,2959
:|2959,2960
[|2961,2962
x|2962,2963
]|2963,2964
Yes|2964,2967
[|2968,2969
]|2970,2971
No|2971,2973
<EOL>|2973,2974
<EOL>|2974,2975
Comprehension|2975,2988
Intact|2989,2995
:|2995,2996
[|2997,2998
x|2998,2999
]|2999,3000
Yes|3000,3003
[|3004,3005
]|3006,3007
No|3007,3009
<EOL>|3009,3010
<EOL>|3010,3011
Motor|3011,3016
:|3016,3017
<EOL>|3017,3018
TrapDeltoid|3018,3029
BicepTricepGrip|3031,3046
<EOL>|3046,3047
Right|3047,3052
5|3053,3054
5|3063,3064
5|3070,3071
5|3079,3080
5|3086,3087
<EOL>|3087,3088
Left|3088,3092
5|3093,3094
5|3103,3104
5|3110,3111
5|3119,3120
5|3126,3127
<EOL>|3127,3128
<EOL>|3128,3129
IPQuadHamATEHLGast|3129,3147
<EOL>|3147,3148
Right5|3148,3154
5|3162,3163
5|3170,3171
5|3177,3178
5|3186,3187
5|3195,3196
<EOL>|3196,3197
Left5|3197,3202
5|3210,3211
5|3218,3219
5|3225,3226
5|3234,3235
5|3243,3244
<EOL>|3244,3245
<EOL>|3245,3246
[|3246,3247
x|3247,3248
]|3248,3249
Sensation|3249,3258
intact|3259,3265
to|3266,3268
light|3269,3274
touch|3275,3280
<EOL>|3280,3281
<EOL>|3281,3282
<EOL>|3283,3284
Pertinent|3284,3293
Results|3294,3301
:|3301,3302
<EOL>|3302,3303
Please|3303,3309
see|3310,3313
OMR|3314,3317
for|3318,3321
pertinent|3322,3331
lab|3332,3335
and|3336,3339
imaging|3340,3347
results|3348,3355
.|3355,3356
<EOL>|3356,3357
<EOL>|3358,3359
Brief|3359,3364
Hospital|3365,3373
Course|3374,3380
:|3380,3381
<EOL>|3381,3382
#|3382,3383
Brain|3383,3388
lesion|3389,3395
<EOL>|3395,3396
Patient|3396,3403
was|3404,3407
found|3408,3413
to|3414,3416
have|3417,3421
cerebellar|3422,3432
hypodensity|3433,3444
on|3445,3447
NCHCT|3448,3453
from|3454,3458
<EOL>|3459,3460
OSH|3460,3463
.|3463,3464
CT|3465,3467
w|3468,3469
/|3469,3470
wo|3470,3472
contrast|3473,3481
was|3482,3485
obtained|3486,3494
while|3495,3500
in|3501,3503
the|3504,3507
ED|3508,3510
at|3511,3513
_|3514,3515
_|3515,3516
_|3516,3517
<EOL>|3518,3519
which|3519,3524
was|3525,3528
concerning|3529,3539
for|3540,3543
underlying|3544,3554
mass|3555,3559
lesion|3560,3566
and|3567,3570
<EOL>|3571,3572
hydrocephalus|3572,3585
.|3585,3586
(|3587,3588
Of|3588,3590
note|3591,3595
,|3595,3596
she|3597,3600
was|3601,3604
unable|3605,3611
to|3612,3614
get|3615,3618
MRI|3619,3622
due|3623,3626
to|3627,3629
<EOL>|3630,3631
reportedly|3631,3641
having|3642,3648
a|3649,3650
non-compatible|3651,3665
aneurysm|3666,3674
clip|3675,3679
that|3680,3684
was|3685,3688
placed|3689,3695
<EOL>|3696,3697
in|3697,3699
_|3700,3701
_|3701,3702
_|3702,3703
at|3704,3706
_|3707,3708
_|3708,3709
_|3709,3710
.|3710,3711
Patient|3712,3719
was|3720,3723
admitted|3724,3732
to|3733,3735
the|3736,3739
_|3740,3741
_|3741,3742
_|3742,3743
for|3744,3747
close|3748,3753
<EOL>|3754,3755
monitoring|3755,3765
and|3766,3769
surgical|3770,3778
planning|3779,3787
.|3787,3788
She|3789,3792
was|3793,3796
started|3797,3804
on|3805,3807
<EOL>|3808,3809
dexamethasone|3809,3822
4mg|3823,3826
Q6hr|3827,3831
for|3832,3835
mass|3836,3840
effect|3841,3847
.|3847,3848
CT|3849,3851
torso|3852,3857
was|3858,3861
obtained|3862,3870
<EOL>|3871,3872
which|3872,3877
showed|3878,3884
two|3885,3888
lung|3889,3893
nodules|3894,3901
,|3901,3902
see|3903,3906
below|3907,3912
for|3913,3916
more|3917,3921
information|3922,3933
.|3933,3934
<EOL>|3935,3936
Neuro|3936,3941
and|3942,3945
radiation|3946,3955
oncology|3956,3964
were|3965,3969
consulted|3970,3979
.|3979,3980
Plan|3981,3985
was|3986,3989
made|3990,3994
for|3995,3998
<EOL>|3999,4000
surgical|4000,4008
resection|4009,4018
of|4019,4021
the|4022,4025
lesion|4026,4032
.|4032,4033
On|4034,4036
_|4037,4038
_|4038,4039
_|4039,4040
,|4040,4041
it|4042,4044
was|4045,4048
determined|4049,4059
<EOL>|4060,4061
that|4061,4065
her|4066,4069
aneurysm|4070,4078
clip|4079,4083
was|4084,4087
MRI|4088,4091
compatible|4092,4102
and|4103,4106
she|4107,4110
was|4111,4114
able|4115,4119
to|4120,4122
<EOL>|4123,4124
have|4124,4128
a|4129,4130
MRI|4131,4134
Brain|4135,4140
for|4141,4144
surgical|4145,4153
planning|4154,4162
.|4162,4163
She|4164,4167
went|4168,4172
to|4173,4175
the|4176,4179
OR|4180,4182
the|4183,4186
<EOL>|4187,4188
evening|4188,4195
of|4196,4198
_|4199,4200
_|4200,4201
_|4201,4202
for|4203,4206
a|4207,4208
suboccipital|4209,4221
craniotomy|4222,4232
for|4233,4236
resection|4237,4246
of|4247,4249
<EOL>|4250,4251
her|4251,4254
cerebellar|4255,4265
lesion|4266,4272
.|4272,4273
Postoperatively|4274,4289
she|4290,4293
was|4294,4297
monitored|4298,4307
in|4308,4310
<EOL>|4311,4312
Neuro|4312,4317
ICU|4318,4321
,|4321,4322
where|4323,4328
she|4329,4332
remained|4333,4341
neurologically|4342,4356
and|4357,4360
hemodynamically|4361,4376
<EOL>|4377,4378
stable|4378,4384
.|4384,4385
She|4386,4389
was|4390,4393
transferred|4394,4405
to|4406,4408
the|4409,4412
_|4413,4414
_|4414,4415
_|4415,4416
on|4417,4419
POD|4420,4423
#|4423,4424
2|4424,4425
and|4426,4429
made|4430,4434
floor|4435,4440
<EOL>|4441,4442
status|4442,4448
.|4448,4449
Her|4450,4453
Dexamethasone|4454,4467
was|4468,4471
ordered|4472,4479
to|4480,4482
taper|4483,4488
down|4489,4493
to|4494,4496
a|4497,4498
<EOL>|4499,4500
maintenance|4500,4511
dose|4512,4516
of|4517,4519
2mg|4520,4523
BID|4524,4527
over|4528,4532
the|4533,4536
course|4537,4543
of|4544,4546
one|4547,4550
week|4551,4555
.|4555,4556
Her|4557,4560
<EOL>|4561,4562
pathology|4562,4571
finalized|4572,4581
as|4582,4584
small|4585,4590
cell|4591,4595
lung|4596,4600
carcinoma|4601,4610
.|4610,4611
<EOL>|4612,4613
<EOL>|4613,4614
#|4614,4615
Lung|4615,4619
lesions|4620,4627
<EOL>|4627,4628
CT|4628,4630
torso|4631,4636
was|4637,4640
obtained|4641,4649
which|4650,4655
showed|4656,4662
two|4663,4666
lung|4667,4671
nodules|4672,4679
,|4679,4680
one|4681,4684
in|4685,4687
the|4688,4691
<EOL>|4692,4693
left|4693,4697
paramedian|4698,4708
abutting|4709,4717
the|4718,4721
aortic|4722,4728
arch|4729,4733
and|4734,4737
the|4738,4741
other|4742,4747
in|4748,4750
the|4751,4754
<EOL>|4755,4756
right|4756,4761
upper|4762,4767
lobe|4768,4772
.|4772,4773
Pulmonary|4774,4783
was|4784,4787
consulted|4788,4797
and|4798,4801
stated|4802,4808
that|4809,4813
no|4814,4816
<EOL>|4817,4818
further|4818,4825
intervention|4826,4838
was|4839,4842
indicated|4843,4852
until|4853,4858
final|4859,4864
pathology|4865,4874
was|4875,4878
<EOL>|4879,4880
back|4880,4884
.|4884,4885
Heme|4886,4890
-|4890,4891
Onc|4891,4894
was|4895,4898
also|4899,4903
consulted|4904,4913
,|4913,4914
and|4915,4918
made|4919,4923
recommendations|4924,4939
that|4940,4944
<EOL>|4945,4946
no|4946,4948
further|4949,4956
lung|4957,4961
imaging|4962,4969
or|4970,4972
separate|4973,4981
lung|4982,4986
biopsy|4987,4993
was|4994,4997
needed|4998,5004
.|5004,5005
Both|5006,5010
<EOL>|5011,5012
Pulmonary|5012,5021
and|5022,5025
Heme|5026,5030
-|5030,5031
Onc|5031,5034
stated|5035,5041
that|5042,5046
staging|5047,5054
and|5055,5058
treatment|5059,5068
could|5069,5074
<EOL>|5075,5076
be|5076,5078
determined|5079,5089
based|5090,5095
on|5096,5098
the|5099,5102
tissue|5103,5109
pathology|5110,5119
from|5120,5124
resection|5125,5134
of|5135,5137
<EOL>|5138,5139
the|5139,5142
brain|5143,5148
lesion|5149,5155
.|5155,5156
Her|5157,5160
final|5161,5166
pathology|5167,5176
came|5177,5181
back|5182,5186
as|5187,5189
small|5190,5195
cell|5196,5200
<EOL>|5201,5202
lung|5202,5206
carcinoma|5207,5216
.|5216,5217
She|5218,5221
will|5222,5226
follow|5227,5233
-|5233,5234
up|5234,5236
with|5237,5241
the|5242,5245
thoracic|5246,5254
oncologist|5255,5265
<EOL>|5266,5267
on|5267,5269
_|5270,5271
_|5271,5272
_|5272,5273
.|5273,5274
<EOL>|5275,5276
<EOL>|5276,5277
#|5277,5278
Steroid|5278,5285
-|5285,5286
induced|5286,5293
hyperglycemia|5294,5307
<EOL>|5307,5308
Throughout|5308,5318
her|5319,5322
admission|5323,5332
,|5332,5333
the|5334,5337
patient|5338,5345
intermittently|5346,5360
required|5361,5369
<EOL>|5370,5371
sliding|5371,5378
scale|5379,5384
Insulin|5385,5392
for|5393,5396
elevated|5397,5405
blood|5406,5411
sugars|5412,5418
while|5419,5424
on|5425,5427
<EOL>|5428,5429
Dexamethasone|5429,5442
.|5442,5443
She|5444,5447
was|5448,5451
evaluated|5452,5461
by|5462,5464
the|5465,5468
_|5469,5470
_|5470,5471
_|5471,5472
inpatient|5473,5482
team|5483,5487
on|5488,5490
<EOL>|5491,5492
_|5492,5493
_|5493,5494
_|5494,5495
,|5495,5496
who|5497,5500
decided|5501,5508
that|5509,5513
she|5514,5517
did|5518,5521
not|5522,5525
need|5526,5530
to|5531,5533
go|5534,5536
home|5537,5541
on|5542,5544
Insulin|5545,5552
.|5552,5553
<EOL>|5554,5555
They|5555,5559
recommended|5560,5571
discharging|5572,5583
her|5584,5587
with|5588,5592
a|5593,5594
glucometer|5595,5605
so|5606,5608
that|5609,5613
she|5614,5617
<EOL>|5618,5619
could|5619,5624
check|5625,5630
her|5631,5634
blood|5635,5640
sugars|5641,5647
daily|5648,5653
with|5654,5658
a|5659,5660
goal|5661,5665
blood|5666,5671
sugar|5672,5677
less|5678,5682
<EOL>|5683,5684
than|5684,5688
200|5689,5692
.|5692,5693
She|5694,5697
was|5698,5701
advised|5702,5709
to|5710,5712
record|5713,5719
her|5720,5723
readings|5724,5732
and|5733,5736
follow|5737,5743
-|5743,5744
up|5744,5746
<EOL>|5747,5748
with|5748,5752
her|5753,5756
PCP|5757,5760
and|5761,5764
_|5765,5766
_|5766,5767
_|5767,5768
.|5768,5769
<EOL>|5770,5771
<EOL>|5771,5772
#|5772,5773
Bradycardia|5773,5784
<EOL>|5784,5785
She|5785,5788
was|5789,5792
due|5793,5796
to|5797,5799
transfer|5800,5808
out|5809,5812
to|5813,5815
the|5816,5819
_|5820,5821
_|5821,5822
_|5822,5823
on|5824,5826
POD1|5827,5831
,|5831,5832
however|5833,5840
was|5841,5844
<EOL>|5845,5846
kept|5846,5850
in|5851,5853
the|5854,5857
ICU|5858,5861
for|5862,5865
asymptomatic|5866,5878
bradycardia|5879,5890
to|5891,5893
the|5894,5897
_|5898,5899
_|5899,5900
_|5900,5901
.|5901,5902
She|5903,5906
<EOL>|5907,5908
remained|5908,5916
asymptomatic|5917,5929
,|5929,5930
and|5931,5934
her|5935,5938
heartrate|5939,5948
improved|5949,5957
with|5958,5962
fluids|5963,5969
,|5969,5970
<EOL>|5971,5972
and|5972,5975
administration|5976,5990
of|5991,5993
her|5994,5997
levothyroxine|5998,6011
.|6011,6012
She|6013,6016
intermittently|6017,6031
<EOL>|6032,6033
dipped|6033,6039
to|6040,6042
the|6043,6046
_|6047,6048
_|6048,6049
_|6049,6050
,|6050,6051
however|6052,6059
remained|6060,6068
asymptomatic|6069,6081
.|6081,6082
<EOL>|6082,6083
<EOL>|6083,6084
#|6084,6085
Bell|6085,6089
's|6089,6091
palsy|6092,6097
<EOL>|6097,6098
The|6098,6101
patient|6102,6109
was|6110,6113
resumed|6114,6121
on|6122,6124
her|6125,6128
home|6129,6133
Valacyclovir|6134,6146
and|6147,6150
Prenisolone|6151,6162
<EOL>|6163,6164
gtts|6164,6168
.|6168,6169
<EOL>|6170,6171
<EOL>|6171,6172
#|6172,6173
Urinary|6173,6180
urgency|6181,6188
<EOL>|6188,6189
On|6189,6191
POD|6192,6195
2|6196,6197
,|6197,6198
the|6199,6202
patient|6203,6210
complained|6211,6221
of|6222,6224
urinary|6225,6232
urgency|6233,6240
and|6241,6244
<EOL>|6245,6246
increased|6246,6255
frequency|6256,6265
.|6265,6266
U|6267,6268
/|6268,6269
A|6269,6270
was|6271,6274
negative|6275,6283
and|6284,6287
culture|6288,6295
was|6296,6299
negative|6300,6308
.|6308,6309
<EOL>|6310,6311
Her|6311,6314
symptoms|6315,6323
had|6324,6327
resolved|6328,6336
at|6337,6339
the|6340,6343
time|6344,6348
of|6349,6351
discharge|6352,6361
.|6361,6362
<EOL>|6362,6363
<EOL>|6363,6364
#|6364,6365
Dispo|6365,6370
<EOL>|6371,6372
The|6372,6375
patient|6376,6383
was|6384,6387
evaluated|6388,6397
by|6398,6400
_|6401,6402
_|6402,6403
_|6403,6404
and|6405,6408
OT|6409,6411
who|6412,6415
cleared|6416,6423
her|6424,6427
for|6428,6431
home|6432,6436
<EOL>|6437,6438
with|6438,6442
services|6443,6451
.|6451,6452
She|6453,6456
was|6457,6460
discharged|6461,6471
on|6472,6474
_|6475,6476
_|6476,6477
_|6477,6478
in|6479,6481
stable|6482,6488
condition|6489,6498
.|6498,6499
<EOL>|6500,6501
She|6501,6504
will|6505,6509
follow|6510,6516
up|6517,6519
in|6520,6522
_|6523,6524
_|6524,6525
_|6525,6526
on|6527,6529
_|6530,6531
_|6531,6532
_|6532,6533
.|6533,6534
<EOL>|6535,6536
<EOL>|6537,6538
Medications|6538,6549
on|6550,6552
Admission|6553,6562
:|6562,6563
<EOL>|6563,6564
-|6564,6565
ASA|6566,6569
81mg|6570,6574
<EOL>|6574,6575
-|6575,6576
Alendronate|6577,6588
70mg|6589,6593
weekly|6594,6600
<EOL>|6600,6601
-|6601,6602
Vitamin|6603,6610
D3|6611,6613
_|6614,6615
_|6615,6616
_|6616,6617
units|6618,6623
daily|6624,6629
<EOL>|6629,6630
-|6630,6631
Levothyroxine|6632,6645
88mcg|6646,6651
daily|6652,6657
<EOL>|6657,6658
-|6658,6659
Lisinopril|6660,6670
20mg|6671,6675
daily|6676,6681
<EOL>|6681,6682
<EOL>|6682,6683
<EOL>|6684,6685
Discharge|6685,6694
Medications|6695,6706
:|6706,6707
<EOL>|6707,6708
1.|6708,6710
Acetaminophen|6712,6725
650|6726,6729
mg|6730,6732
PO|6733,6735
Q6H|6736,6739
:|6739,6740
PRN|6740,6743
Pain|6744,6748
-|6749,6750
Mild|6751,6755
/|6755,6756
Fever|6756,6761
<EOL>|6763,6764
2.|6764,6766
Bisacodyl|6768,6777
10|6778,6780
mg|6781,6783
PO|6784,6786
/|6786,6787
PR|6787,6789
DAILY|6790,6795
<EOL>|6797,6798
3.|6798,6800
Dexamethasone|6802,6815
3|6816,6817
mg|6818,6820
PO|6821,6823
Q8H|6824,6827
Duration|6828,6836
:|6836,6837
6|6838,6839
Doses|6840,6845
<EOL>|6846,6847
start|6847,6852
_|6853,6854
_|6854,6855
_|6855,6856
:|6856,6857
3tabsq8hrs|6858,6868
x2|6869,6871
,|6871,6872
2tabsq8hrs|6873,6883
x6|6884,6886
,|6886,6887
2tabsq12hrs|6888,6899
<EOL>|6900,6901
maintenance|6901,6912
dose|6913,6917
.|6917,6918
<EOL>|6920,6921
This|6921,6925
is|6926,6928
dose|6929,6933
#|6934,6935
2|6936,6937
of|6938,6940
3|6941,6942
tapered|6943,6950
doses|6951,6956
<EOL>|6956,6957
RX|6957,6959
*|6960,6961
dexamethasone|6961,6974
1|6975,6976
mg|6977,6979
3|6980,6981
tablet|6982,6988
(|6988,6989
s|6989,6990
)|6990,6991
by|6992,6994
mouth|6995,7000
every|7001,7006
eight|7007,7012
(|7013,7014
8|7014,7015
)|7015,7016
<EOL>|7017,7018
hours|7018,7023
Disp|7024,7028
#|7029,7030
*|7030,7031
120|7031,7034
Tablet|7035,7041
Refills|7042,7049
:|7049,7050
*|7050,7051
1|7051,7052
<EOL>|7053,7054
4.|7054,7056
Docusate|7058,7066
Sodium|7067,7073
100|7074,7077
mg|7078,7080
PO|7081,7083
BID|7084,7087
<EOL>|7089,7090
5.|7090,7092
Famotidine|7094,7104
20|7105,7107
mg|7108,7110
PO|7111,7113
Q24H|7114,7118
<EOL>|7119,7120
RX|7120,7122
*|7123,7124
famotidine|7124,7134
20|7135,7137
mg|7138,7140
1|7141,7142
tablet|7143,7149
(|7149,7150
s|7150,7151
)|7151,7152
by|7153,7155
mouth|7156,7161
twice|7162,7167
a|7168,7169
day|7170,7173
Disp|7174,7178
#|7179,7180
*|7180,7181
60|7181,7183
<EOL>|7184,7185
Tablet|7185,7191
Refills|7192,7199
:|7199,7200
*|7200,7201
1|7201,7202
<EOL>|7203,7204
6.|7204,7206
Polyethylene|7208,7220
Glycol|7221,7227
17|7228,7230
g|7231,7232
PO|7233,7235
DAILY|7236,7241
:|7241,7242
PRN|7242,7245
Constipation|7246,7258
-|7259,7260
First|7261,7266
<EOL>|7267,7268
Line|7268,7272
<EOL>|7274,7275
7.|7275,7277
Senna|7279,7284
17.2|7285,7289
mg|7290,7292
PO|7293,7295
HS|7296,7298
<EOL>|7300,7301
8.|7301,7303
Levothyroxine|7305,7318
Sodium|7319,7325
88|7326,7328
mcg|7329,7332
PO|7333,7335
DAILY|7336,7341
<EOL>|7343,7344
9.|7344,7346
Lisinopril|7348,7358
20|7359,7361
mg|7362,7364
PO|7365,7367
DAILY|7368,7373
<EOL>|7375,7376
10.|7376,7379
PrednisoLONE|7381,7393
Acetate|7394,7401
1|7402,7403
%|7403,7404
Ophth|7405,7410
.|7410,7411
Susp.|7412,7417
1|7418,7419
DROP|7420,7424
LEFT|7425,7429
EYE|7430,7433
QID|7434,7437
<EOL>|7439,7440
11.|7440,7443
ValACYclovir|7445,7457
1000|7458,7462
mg|7463,7465
PO|7466,7468
Q8H|7469,7472
<EOL>|7474,7475
12.|7475,7478
Vitamin|7480,7487
D|7488,7489
_|7490,7491
_|7491,7492
_|7492,7493
UNIT|7494,7498
PO|7499,7501
DAILY|7502,7507
<EOL>|7509,7510
13.|7510,7513
HELD|7514,7518
-|7518,7519
Alendronate|7520,7531
Sodium|7532,7538
70|7539,7541
mg|7542,7544
PO|7545,7547
1X|7548,7550
/|7550,7551
WEEK|7551,7555
(|7556,7557
_|7557,7558
_|7558,7559
_|7559,7560
)|7560,7561
This|7563,7567
<EOL>|7568,7569
medication|7569,7579
was|7580,7583
held|7584,7588
.|7588,7589
Do|7590,7592
not|7593,7596
restart|7597,7604
Alendronate|7605,7616
Sodium|7617,7623
until|7624,7629
POD|7630,7633
<EOL>|7634,7635
_|7635,7636
_|7636,7637
_|7637,7638
-|7639,7640
_|7641,7642
_|7642,7643
_|7643,7644
<EOL>|7644,7645
14.|7645,7648
HELD|7649,7653
-|7653,7654
Aspirin|7655,7662
81|7663,7665
mg|7666,7668
PO|7669,7671
DAILY|7672,7677
This|7679,7683
medication|7684,7694
was|7695,7698
held|7699,7703
.|7703,7704
Do|7705,7707
<EOL>|7708,7709
not|7709,7712
restart|7713,7720
Aspirin|7721,7728
until|7729,7734
POD|7735,7738
14|7739,7741
-|7742,7743
_|7744,7745
_|7745,7746
_|7746,7747
<EOL>|7747,7748
_|7748,7749
_|7749,7750
_|7750,7751
glucometer|7752,7762
<EOL>|7762,7763
_|7763,7764
_|7764,7765
_|7765,7766
Freestyle|7767,7776
glucometer|7777,7787
.|7787,7788
Check|7789,7794
blood|7795,7800
sugars|7801,7807
_|7808,7809
_|7809,7810
_|7810,7811
hours|7812,7817
after|7818,7823
a|7824,7825
<EOL>|7826,7827
starchy|7827,7834
meal|7835,7839
.|7839,7840
Record|7841,7847
numbers|7848,7855
and|7856,7859
show|7860,7864
to|7865,7867
your|7868,7872
Oncologist|7873,7883
.|7883,7884
<EOL>|7885,7886
_|7886,7887
_|7887,7888
_|7888,7889
test|7890,7894
strips|7895,7901
<EOL>|7901,7902
#|7902,7903
50|7903,7905
.|7905,7906
Check|7907,7912
blood|7913,7918
sugars|7919,7925
QD.|7926,7929
3|7930,7931
refills|7932,7939
.|7939,7940
<EOL>|7942,7943
_|7943,7944
_|7944,7945
_|7945,7946
Lancets|7947,7954
<EOL>|7954,7955
#|7955,7956
50|7956,7958
.|7958,7959
Check|7960,7965
blood|7966,7971
sugars|7972,7978
QD.|7979,7982
3|7983,7984
refills|7985,7992
.|7992,7993
<EOL>|7994,7995
<EOL>|7995,7996
<EOL>|7997,7998
Discharge|7998,8007
Disposition|8008,8019
:|8019,8020
<EOL>|8020,8021
Home|8021,8025
With|8026,8030
Service|8031,8038
<EOL>|8038,8039
<EOL>|8040,8041
Facility|8041,8049
:|8049,8050
<EOL>|8050,8051
_|8051,8052
_|8052,8053
_|8053,8054
<EOL>|8054,8055
<EOL>|8056,8057
Discharge|8057,8066
Diagnosis|8067,8076
:|8076,8077
<EOL>|8077,8078
Brain|8078,8083
tumor|8084,8089
<EOL>|8089,8090
<EOL>|8090,8091
<EOL>|8092,8093
Discharge|8093,8102
Condition|8103,8112
:|8112,8113
<EOL>|8113,8114
Mental|8114,8120
Status|8121,8127
:|8127,8128
Clear|8129,8134
and|8135,8138
coherent|8139,8147
.|8147,8148
<EOL>|8148,8149
Level|8149,8154
of|8155,8157
Consciousness|8158,8171
:|8171,8172
Alert|8173,8178
and|8179,8182
interactive|8183,8194
.|8194,8195
<EOL>|8195,8196
Activity|8196,8204
Status|8205,8211
:|8211,8212
Ambulatory|8213,8223
-|8224,8225
requires|8226,8234
assistance|8235,8245
or|8246,8248
aid|8249,8252
.|8252,8253
<EOL>|8253,8254
<EOL>|8254,8255
<EOL>|8256,8257
Discharge|8257,8266
Instructions|8267,8279
:|8279,8280
<EOL>|8280,8281
Surgery|8281,8288
:|8288,8289
<EOL>|8289,8290
<EOL>|8290,8291
-|8291,8292
You|8293,8296
underwent|8297,8306
surgery|8307,8314
to|8315,8317
remove|8318,8324
a|8325,8326
brain|8327,8332
lesion|8333,8339
from|8340,8344
your|8345,8349
<EOL>|8350,8351
brain|8351,8356
.|8356,8357
<EOL>|8358,8359
<EOL>|8359,8360
-|8360,8361
A|8362,8363
sample|8364,8370
of|8371,8373
tissue|8374,8380
from|8381,8385
the|8386,8389
lesion|8390,8396
in|8397,8399
your|8400,8404
brain|8405,8410
was|8411,8414
sent|8415,8419
to|8420,8422
<EOL>|8423,8424
pathology|8424,8433
for|8434,8437
testing|8438,8445
.|8445,8446
<EOL>|8447,8448
<EOL>|8448,8449
-|8449,8450
Please|8451,8457
keep|8458,8462
your|8463,8467
incision|8468,8476
dry|8477,8480
until|8481,8486
your|8487,8491
sutures|8492,8499
are|8500,8503
removed|8504,8511
.|8511,8512
<EOL>|8513,8514
<EOL>|8514,8515
-|8515,8516
You|8517,8520
may|8521,8524
shower|8525,8531
at|8532,8534
this|8535,8539
time|8540,8544
but|8545,8548
keep|8549,8553
your|8554,8558
incision|8559,8567
dry|8568,8571
.|8571,8572
<EOL>|8572,8573
<EOL>|8573,8574
-|8574,8575
It|8576,8578
is|8579,8581
best|8582,8586
to|8587,8589
keep|8590,8594
your|8595,8599
incision|8600,8608
open|8609,8613
to|8614,8616
air|8617,8620
but|8621,8624
it|8625,8627
is|8628,8630
ok|8631,8633
to|8634,8636
<EOL>|8637,8638
cover|8638,8643
it|8644,8646
when|8647,8651
outside|8652,8659
.|8659,8660
<EOL>|8661,8662
<EOL>|8662,8663
-|8663,8664
Call|8665,8669
your|8670,8674
surgeon|8675,8682
if|8683,8685
there|8686,8691
are|8692,8695
any|8696,8699
signs|8700,8705
of|8706,8708
infection|8709,8718
like|8719,8723
<EOL>|8724,8725
redness|8725,8732
,|8732,8733
fever|8734,8739
,|8739,8740
or|8741,8743
drainage|8744,8752
.|8752,8753
<EOL>|8754,8755
<EOL>|8755,8756
Activity|8756,8764
:|8764,8765
<EOL>|8765,8766
<EOL>|8766,8767
-|8767,8768
We|8769,8771
recommend|8772,8781
that|8782,8786
you|8787,8790
avoid|8791,8796
heavy|8797,8802
lifting|8803,8810
,|8810,8811
running|8812,8819
,|8819,8820
climbing|8821,8829
,|8829,8830
<EOL>|8831,8832
or|8832,8834
other|8835,8840
strenuous|8841,8850
exercise|8851,8859
until|8860,8865
your|8866,8870
follow|8871,8877
-|8877,8878
up|8878,8880
appointment|8881,8892
.|8892,8893
<EOL>|8893,8894
<EOL>|8894,8895
-|8895,8896
You|8897,8900
make|8901,8905
take|8906,8910
leisurely|8911,8920
walks|8921,8926
and|8927,8930
slowly|8931,8937
increase|8938,8946
your|8947,8951
<EOL>|8952,8953
activity|8953,8961
at|8962,8964
your|8965,8969
own|8970,8973
pace|8974,8978
once|8979,8983
you|8984,8987
are|8988,8991
symptom|8992,8999
free|9000,9004
at|9005,9007
rest|9008,9012
.|9012,9013
<EOL>|9014,9015
_|9015,9016
_|9016,9017
_|9017,9018
try|9019,9022
to|9023,9025
do|9026,9028
too|9029,9032
much|9033,9037
all|9038,9041
at|9042,9044
once|9045,9049
.|9049,9050
<EOL>|9050,9051
<EOL>|9051,9052
-|9052,9053
No|9054,9056
driving|9057,9064
while|9065,9070
taking|9071,9077
any|9078,9081
narcotic|9082,9090
or|9091,9093
sedating|9094,9102
medication|9103,9113
.|9113,9114
<EOL>|9115,9116
<EOL>|9116,9117
-|9117,9118
If|9119,9121
you|9122,9125
experienced|9126,9137
a|9138,9139
seizure|9140,9147
while|9148,9153
admitted|9154,9162
,|9162,9163
you|9164,9167
are|9168,9171
NOT|9172,9175
<EOL>|9176,9177
allowed|9177,9184
to|9185,9187
drive|9188,9193
by|9194,9196
law|9197,9200
.|9200,9201
<EOL>|9202,9203
<EOL>|9203,9204
-|9204,9205
No|9206,9208
contact|9209,9216
sports|9217,9223
until|9224,9229
cleared|9230,9237
by|9238,9240
your|9241,9245
neurosurgeon|9246,9258
.|9258,9259
You|9260,9263
<EOL>|9264,9265
should|9265,9271
avoid|9272,9277
contact|9278,9285
sports|9286,9292
for|9293,9296
6|9297,9298
months|9299,9305
.|9305,9306
<EOL>|9307,9308
<EOL>|9308,9309
Medications|9309,9320
:|9320,9321
<EOL>|9321,9322
<EOL>|9322,9323
-|9323,9324
Please|9325,9331
do|9332,9334
NOT|9335,9338
take|9339,9343
any|9344,9347
blood|9348,9353
thinning|9354,9362
medication|9363,9373
(|9374,9375
Aspirin|9375,9382
,|9382,9383
<EOL>|9384,9385
Ibuprofen|9385,9394
,|9394,9395
Plavix|9396,9402
,|9402,9403
Coumadin|9404,9412
)|9412,9413
until|9414,9419
cleared|9420,9427
by|9428,9430
the|9431,9434
neurosurgeon|9435,9447
.|9447,9448
<EOL>|9449,9450
We|9450,9452
held|9453,9457
your|9458,9462
Aspirin|9463,9470
81mg|9471,9475
daily|9476,9481
.|9481,9482
You|9483,9486
are|9487,9490
cleared|9491,9498
to|9499,9501
resume|9502,9508
this|9509,9513
<EOL>|9514,9515
medication|9515,9525
on|9526,9528
POD|9529,9532
14|9533,9535
(|9536,9537
_|9537,9538
_|9538,9539
_|9539,9540
)|9540,9541
.|9541,9542
<EOL>|9543,9544
<EOL>|9544,9545
-|9545,9546
We|9547,9549
held|9550,9554
your|9555,9559
home|9560,9564
Alendronate|9565,9576
during|9577,9583
this|9584,9588
admission|9589,9598
.|9598,9599
You|9600,9603
are|9604,9607
<EOL>|9608,9609
cleared|9609,9616
to|9617,9619
resume|9620,9626
this|9627,9631
medication|9632,9642
on|9643,9645
POD|9646,9649
14|9650,9652
(|9653,9654
_|9654,9655
_|9655,9656
_|9656,9657
)|9657,9658
.|9658,9659
<EOL>|9660,9661
<EOL>|9661,9662
-|9662,9663
You|9664,9667
may|9668,9671
use|9672,9675
Acetaminophen|9676,9689
(|9690,9691
Tylenol|9691,9698
)|9698,9699
for|9700,9703
minor|9704,9709
discomfort|9710,9720
if|9721,9723
<EOL>|9724,9725
you|9725,9728
are|9729,9732
not|9733,9736
otherwise|9737,9746
restricted|9747,9757
from|9758,9762
taking|9763,9769
this|9770,9774
medication|9775,9785
.|9785,9786
<EOL>|9786,9787
<EOL>|9787,9788
-|9788,9789
You|9790,9793
were|9794,9798
started|9799,9806
on|9807,9809
Dexamethasone|9810,9823
,|9823,9824
a|9825,9826
steroid|9827,9834
that|9835,9839
treats|9840,9846
<EOL>|9847,9848
intracranial|9848,9860
swelling|9861,9869
.|9869,9870
This|9871,9875
Dexamethasone|9876,9889
is|9890,9892
being|9893,9898
tapered|9899,9906
down|9907,9911
<EOL>|9912,9913
to|9913,9915
a|9916,9917
maintenance|9918,9929
dose|9930,9934
of|9935,9937
2mg|9938,9941
BID|9942,9945
.|9945,9946
Please|9947,9953
take|9954,9958
this|9959,9963
medication|9964,9974
as|9975,9977
<EOL>|9978,9979
prescribed|9979,9989
.|9989,9990
<EOL>|9990,9991
<EOL>|9991,9992
-|9992,9993
While|9994,9999
admitted|10000,10008
,|10008,10009
you|10010,10013
had|10014,10017
elevated|10018,10026
blood|10027,10032
glucose|10033,10040
levels|10041,10047
that|10048,10052
<EOL>|10053,10054
needed|10054,10060
to|10061,10063
be|10064,10066
treated|10067,10074
by|10075,10077
Insulin|10078,10085
.|10085,10086
You|10087,10090
should|10091,10097
continue|10098,10106
to|10107,10109
check|10110,10115
<EOL>|10116,10117
your|10117,10121
blood|10122,10127
sugars|10128,10134
daily|10135,10140
at|10141,10143
home|10144,10148
with|10149,10153
the|10154,10157
prescribed|10158,10168
glucometer|10169,10179
.|10179,10180
<EOL>|10181,10182
You|10182,10185
visiting|10186,10194
nurse|10195,10200
should|10201,10207
teach|10208,10213
you|10214,10217
how|10218,10221
to|10222,10224
use|10225,10228
this|10229,10233
device|10234,10240
at|10241,10243
<EOL>|10244,10245
home|10245,10249
.|10249,10250
Please|10251,10257
record|10258,10264
your|10265,10269
blood|10270,10275
sugars|10276,10282
and|10283,10286
follow|10287,10293
-|10293,10294
up|10294,10296
with|10297,10301
your|10302,10306
<EOL>|10307,10308
PCP|10308,10311
and|10312,10315
_|10316,10317
_|10317,10318
_|10318,10319
regarding|10320,10329
the|10330,10333
results|10334,10341
.|10341,10342
Your|10343,10347
goal|10348,10352
blood|10353,10358
sugar|10359,10364
<EOL>|10365,10366
is|10366,10368
less|10369,10373
than|10374,10378
200|10379,10382
.|10382,10383
<EOL>|10384,10385
<EOL>|10385,10386
What|10386,10390
You|10391,10394
_|10395,10396
_|10396,10397
_|10397,10398
Experience|10399,10409
:|10409,10410
<EOL>|10410,10411
<EOL>|10411,10412
-|10412,10413
You|10414,10417
may|10418,10421
experience|10422,10432
headaches|10433,10442
and|10443,10446
incisional|10447,10457
pain|10458,10462
.|10462,10463
<EOL>|10464,10465
<EOL>|10465,10466
-|10466,10467
You|10468,10471
may|10472,10475
also|10476,10480
experience|10481,10491
some|10492,10496
post-operative|10497,10511
swelling|10512,10520
around|10521,10527
<EOL>|10528,10529
your|10529,10533
face|10534,10538
and|10539,10542
eyes|10543,10547
.|10547,10548
This|10549,10553
is|10554,10556
normal|10557,10563
after|10564,10569
surgery|10570,10577
and|10578,10581
most|10582,10586
<EOL>|10587,10588
noticeable|10588,10598
on|10599,10601
the|10602,10605
second|10606,10612
and|10613,10616
third|10617,10622
day|10623,10626
of|10627,10629
surgery|10630,10637
.|10637,10638
You|10640,10643
apply|10644,10649
<EOL>|10650,10651
ice|10651,10654
or|10655,10657
a|10658,10659
cool|10660,10664
or|10665,10667
warm|10668,10672
washcloth|10673,10682
to|10683,10685
your|10686,10690
eyes|10691,10695
to|10696,10698
help|10699,10703
with|10704,10708
the|10709,10712
<EOL>|10713,10714
swelling|10714,10722
.|10722,10723
The|10724,10727
swelling|10728,10736
will|10737,10741
be|10742,10744
its|10745,10748
worse|10749,10754
in|10755,10757
the|10758,10761
morning|10762,10769
after|10770,10775
<EOL>|10776,10777
laying|10777,10783
flat|10784,10788
from|10789,10793
sleeping|10794,10802
but|10803,10806
decrease|10807,10815
when|10816,10820
up|10821,10823
.|10823,10824
<EOL>|10825,10826
<EOL>|10826,10827
-|10827,10828
You|10829,10832
may|10833,10836
experience|10837,10847
soreness|10848,10856
with|10857,10861
chewing|10862,10869
.|10869,10870
This|10871,10875
is|10876,10878
normal|10879,10885
from|10886,10890
<EOL>|10891,10892
the|10892,10895
surgery|10896,10903
and|10904,10907
will|10908,10912
improve|10913,10920
with|10921,10925
time|10926,10930
.|10930,10931
Softer|10932,10938
foods|10939,10944
may|10945,10948
be|10949,10951
<EOL>|10952,10953
easier|10953,10959
during|10960,10966
this|10967,10971
time|10972,10976
.|10976,10977
<EOL>|10978,10979
<EOL>|10979,10980
-|10980,10981
Feeling|10982,10989
more|10990,10994
tired|10995,11000
or|11001,11003
restlessness|11004,11016
is|11017,11019
also|11020,11024
common|11025,11031
.|11031,11032
<EOL>|11032,11033
<EOL>|11033,11034
-|11034,11035
Constipation|11036,11048
is|11049,11051
common|11052,11058
.|11058,11059
Be|11060,11062
sure|11063,11067
to|11068,11070
drink|11071,11076
plenty|11077,11083
of|11084,11086
fluids|11087,11093
and|11094,11097
<EOL>|11098,11099
eat|11099,11102
a|11103,11104
high|11105,11109
-|11109,11110
fiber|11110,11115
diet|11116,11120
.|11120,11121
If|11122,11124
you|11125,11128
are|11129,11132
taking|11133,11139
narcotics|11140,11149
(|11150,11151
prescription|11151,11163
<EOL>|11164,11165
pain|11165,11169
medications|11170,11181
)|11181,11182
,|11182,11183
try|11184,11187
an|11188,11190
over-the|11191,11199
-|11199,11200
counter|11200,11207
stool|11208,11213
softener|11214,11222
.|11222,11223
<EOL>|11223,11224
<EOL>|11224,11225
When|11225,11229
to|11230,11232
Call|11233,11237
Your|11238,11242
Doctor|11243,11249
at|11250,11252
_|11253,11254
_|11254,11255
_|11255,11256
for|11257,11260
:|11260,11261
<EOL>|11261,11262
<EOL>|11262,11263
-|11263,11264
Severe|11265,11271
pain|11272,11276
,|11276,11277
swelling|11278,11286
,|11286,11287
redness|11288,11295
or|11296,11298
drainage|11299,11307
from|11308,11312
the|11313,11316
incision|11317,11325
<EOL>|11326,11327
site|11327,11331
.|11331,11332
<EOL>|11333,11334
<EOL>|11334,11335
-|11335,11336
Fever|11337,11342
greater|11343,11350
than|11351,11355
101.5|11356,11361
degrees|11362,11369
Fahrenheit|11370,11380
<EOL>|11380,11381
<EOL>|11381,11382
-|11382,11383
Nausea|11384,11390
and|11391,11394
/|11394,11395
or|11395,11397
vomiting|11398,11406
<EOL>|11406,11407
<EOL>|11407,11408
-|11408,11409
Extreme|11410,11417
sleepiness|11418,11428
and|11429,11432
not|11433,11436
being|11437,11442
able|11443,11447
to|11448,11450
stay|11451,11455
awake|11456,11461
<EOL>|11461,11462
<EOL>|11462,11463
-|11463,11464
Severe|11465,11471
headaches|11472,11481
not|11482,11485
relieved|11486,11494
by|11495,11497
pain|11498,11502
relievers|11503,11512
<EOL>|11512,11513
<EOL>|11513,11514
-|11514,11515
Seizures|11516,11524
<EOL>|11524,11525
<EOL>|11525,11526
-|11526,11527
Any|11528,11531
new|11532,11535
problems|11536,11544
with|11545,11549
your|11550,11554
vision|11555,11561
or|11562,11564
ability|11565,11572
to|11573,11575
speak|11576,11581
<EOL>|11581,11582
<EOL>|11582,11583
-|11583,11584
Weakness|11585,11593
or|11594,11596
changes|11597,11604
in|11605,11607
sensation|11608,11617
in|11618,11620
your|11621,11625
face|11626,11630
,|11630,11631
arms|11632,11636
,|11636,11637
or|11638,11640
leg|11641,11644
<EOL>|11644,11645
<EOL>|11645,11646
Call|11646,11650
_|11651,11652
_|11652,11653
_|11653,11654
and|11655,11658
go|11659,11661
to|11662,11664
the|11665,11668
nearest|11669,11676
Emergency|11677,11686
Room|11687,11691
if|11692,11694
you|11695,11698
experience|11699,11709
<EOL>|11710,11711
any|11711,11714
of|11715,11717
the|11718,11721
following|11722,11731
:|11731,11732
<EOL>|11732,11733
<EOL>|11733,11734
-|11734,11735
Sudden|11736,11742
numbness|11743,11751
or|11752,11754
weakness|11755,11763
in|11764,11766
the|11767,11770
face|11771,11775
,|11775,11776
arm|11777,11780
,|11780,11781
or|11782,11784
leg|11785,11788
<EOL>|11788,11789
<EOL>|11789,11790
-|11790,11791
Sudden|11792,11798
confusion|11799,11808
or|11809,11811
trouble|11812,11819
speaking|11820,11828
or|11829,11831
understanding|11832,11845
<EOL>|11845,11846
<EOL>|11846,11847
-|11847,11848
Sudden|11849,11855
trouble|11856,11863
walking|11864,11871
,|11871,11872
dizziness|11873,11882
,|11882,11883
or|11884,11886
loss|11887,11891
of|11892,11894
balance|11895,11902
or|11903,11905
<EOL>|11906,11907
coordination|11907,11919
<EOL>|11919,11920
<EOL>|11920,11921
-|11921,11922
Sudden|11923,11929
severe|11930,11936
headaches|11937,11946
with|11947,11951
no|11952,11954
known|11955,11960
reason|11961,11967
<EOL>|11967,11968
<EOL>|11968,11969
<EOL>|11970,11971
Followup|11971,11979
Instructions|11980,11992
:|11992,11993
<EOL>|11993,11994
_|11994,11995
_|11995,11996
_|11996,11997
<EOL>|11997,11998

