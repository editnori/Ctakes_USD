 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|164,173|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|185,194|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|210,219|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|222,231|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|246,255|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Event|Event|SIMPLE_SEGMENT|257,263|false|false|false|||Fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|257,263|false|false|false|C0015967|Fever|Fevers
Event|Event|SIMPLE_SEGMENT|268,274|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|268,274|false|false|false|C0085593|Chills|chills
Finding|Classification|SIMPLE_SEGMENT|277,282|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|295,313|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|304,313|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|304,313|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|304,313|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|304,313|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|304,313|false|false|false|C0184661|Interventional procedure|Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|328,336|false|false|false|C4019011|Exchange (clinical)|exchange
Event|Event|SIMPLE_SEGMENT|328,336|false|false|false|||exchange
Finding|Social Behavior|SIMPLE_SEGMENT|328,336|false|false|false|C0678640|degree of relationship - exchange|exchange
Event|Event|SIMPLE_SEGMENT|340,347|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|340,347|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|340,347|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|340,347|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|340,350|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|340,366|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|340,366|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|351,358|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|351,358|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|351,366|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|359,366|false|false|false|C0221423|Illness (finding)|Illness
Finding|Functional Concept|SIMPLE_SEGMENT|406,413|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|406,413|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|406,413|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|406,413|false|false|false|C0199168|Medical service|medical
Finding|Finding|SIMPLE_SEGMENT|406,421|false|false|false|C0262926|Medical History|medical history
Event|Event|SIMPLE_SEGMENT|414,421|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|414,421|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|SIMPLE_SEGMENT|434,441|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|434,441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|434,441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|434,441|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|434,444|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|445,452|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|445,452|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|445,452|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|445,459|true|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|453,459|false|false|false|C0006826|Malignant Neoplasms|cancer
Attribute|Clinical Attribute|SIMPLE_SEGMENT|460,466|false|false|false|C5889824||status
Event|Event|SIMPLE_SEGMENT|460,466|false|false|false|||status
Finding|Idea or Concept|SIMPLE_SEGMENT|460,466|false|false|false|C1546481|What subject filter - Status|status
Finding|Gene or Genome|SIMPLE_SEGMENT|468,472|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Event|Event|SIMPLE_SEGMENT|481,484|false|false|false|||TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|481,484|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|485,488|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|485,488|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|485,488|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Event|Event|SIMPLE_SEGMENT|485,488|false|false|false|||BSO
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|490,493|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|490,493|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|490,493|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|490,493|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|490,493|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|490,493|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|490,493|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|494,501|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|494,512|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|502,512|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|502,512|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|518,523|false|false|false|C0020885|ileum|ileal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|518,528|false|false|false|C1550266|Ileal Loop|ileal loop
Event|Event|SIMPLE_SEGMENT|530,539|false|false|false|||diversion
Finding|Finding|SIMPLE_SEGMENT|530,539|false|false|false|C0439843;C3840275|Diversion|diversion
Finding|Functional Concept|SIMPLE_SEGMENT|530,539|false|false|false|C0439843;C3840275|Diversion|diversion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|530,539|false|false|false|C0185033|Diversion procedure|diversion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|544,552|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|553,564|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|553,564|false|false|false|C0195130|Vaginectomy|vaginectomy
Event|Event|SIMPLE_SEGMENT|572,583|false|false|false|||complicated
Anatomy|Body Location or Region|SIMPLE_SEGMENT|587,596|false|false|false|C0000726|Abdomen|abdominal
Drug|Substance|SIMPLE_SEGMENT|597,602|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|597,602|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|597,602|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|603,612|false|false|false|||requiring
Event|Event|SIMPLE_SEGMENT|613,622|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|613,622|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|613,622|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|626,634|false|false|false|||drainage
Finding|Body Substance|SIMPLE_SEGMENT|626,634|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|SIMPLE_SEGMENT|626,634|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|626,634|false|false|false|C0013103|Drainage procedure|drainage
Event|Event|SIMPLE_SEGMENT|635,644|false|false|false|||catheters
Event|Event|SIMPLE_SEGMENT|654,665|false|false|false|||complicated
Finding|Finding|SIMPLE_SEGMENT|671,677|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|671,677|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|678,702|false|false|false|C0521622|Bilateral hydronephrosis|bilateral hydronephrosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|688,702|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Event|Event|SIMPLE_SEGMENT|688,702|false|false|false|||hydronephrosis
Event|Event|SIMPLE_SEGMENT|703,712|false|false|false|||requiring
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|723,731|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|723,731|false|false|false|C0856443|Urostomy procedure|urostomy
Event|Event|SIMPLE_SEGMENT|732,736|false|false|false|||tube
Finding|Functional Concept|SIMPLE_SEGMENT|732,736|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|SIMPLE_SEGMENT|732,736|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|732,746|false|false|false|C0883304|placement of tube|tube placement
Event|Event|SIMPLE_SEGMENT|737,746|false|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|737,746|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|737,746|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Intellectual Product|SIMPLE_SEGMENT|751,755|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|767,775|false|false|false|C0041951|Ureter|ureteral
Finding|Functional Concept|SIMPLE_SEGMENT|767,775|false|false|false|C1522613|Ureteral Route of Administration|ureteral
Event|Event|SIMPLE_SEGMENT|782,792|false|false|false|||placements
Procedure|Health Care Activity|SIMPLE_SEGMENT|782,792|false|false|false|C0441587|Clinical act of insertion|placements
Event|Event|SIMPLE_SEGMENT|798,809|false|false|false|||improvement
Finding|Conceptual Entity|SIMPLE_SEGMENT|798,809|false|false|false|C2986411|Improvement|improvement
Event|Event|SIMPLE_SEGMENT|814,823|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|831,839|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|844,851|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Finding|Intellectual Product|SIMPLE_SEGMENT|844,851|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|844,851|false|false|false|C1979801|Routine coag|routine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|858,866|false|false|false|C4019011|Exchange (clinical)|exchange
Event|Event|SIMPLE_SEGMENT|858,866|false|false|false|||exchange
Finding|Social Behavior|SIMPLE_SEGMENT|858,866|false|false|false|C0678640|degree of relationship - exchange|exchange
Event|Event|SIMPLE_SEGMENT|871,881|false|false|false|||cystoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|871,881|false|false|false|C0010702|Cystoscopy|cystoscopy
Finding|Body Substance|SIMPLE_SEGMENT|888,895|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|888,895|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|888,895|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|SIMPLE_SEGMENT|924,933|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|924,933|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|924,933|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|924,933|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|924,933|false|false|false|C0184661|Interventional procedure|procedure
Finding|Intellectual Product|SIMPLE_SEGMENT|938,942|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|975,984|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|987,992|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|987,992|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|987,992|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|1010,1021|false|false|false|||tachycardic
Event|Event|SIMPLE_SEGMENT|1042,1046|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|1050,1054|false|false|false|||need
Finding|Functional Concept|SIMPLE_SEGMENT|1050,1054|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Event|Event|SIMPLE_SEGMENT|1055,1064|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1055,1064|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|1055,1078|false|false|false|C0582450|Admission for treatment|admission for treatment
Event|Event|SIMPLE_SEGMENT|1069,1078|false|false|false|||treatment
Finding|Conceptual Entity|SIMPLE_SEGMENT|1069,1078|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|1069,1078|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|1069,1078|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1069,1078|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1082,1088|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|1082,1088|false|false|false|||sepsis
Finding|Finding|SIMPLE_SEGMENT|1100,1104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1100,1104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1100,1104|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Antibiotic|SIMPLE_SEGMENT|1119,1129|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|1119,1129|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|1119,1129|false|false|false|||ampicillin
Drug|Antibiotic|SIMPLE_SEGMENT|1134,1144|false|false|false|C3854019|gentamicin|gentamicin
Drug|Organic Chemical|SIMPLE_SEGMENT|1134,1144|false|false|false|C3854019|gentamicin|gentamicin
Event|Event|SIMPLE_SEGMENT|1134,1144|false|false|false|||gentamicin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1134,1144|false|false|false|C0202391|Gentamicin measurement|gentamicin
Event|Event|SIMPLE_SEGMENT|1155,1162|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1155,1162|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1155,1162|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1155,1162|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1167,1171|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Event|Event|SIMPLE_SEGMENT|1167,1171|false|false|false|||drug
Finding|Finding|SIMPLE_SEGMENT|1167,1171|false|false|false|C0740721|Drug problem|drug
Finding|Functional Concept|SIMPLE_SEGMENT|1172,1181|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Finding|Idea or Concept|SIMPLE_SEGMENT|1172,1181|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1172,1181|false|false|false|C2827757|Antimicrobial Resistance Result|resistant
Event|Event|SIMPLE_SEGMENT|1182,1191|false|false|false|||organisms
Event|Event|SIMPLE_SEGMENT|1198,1206|false|false|false|||reported
Finding|Finding|SIMPLE_SEGMENT|1215,1219|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|1215,1219|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|1215,1219|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|1228,1235|false|false|false|||feeling
Finding|Sign or Symptom|SIMPLE_SEGMENT|1228,1244|false|false|false|C0687681|Feeling feverish|feeling feverish
Event|Event|SIMPLE_SEGMENT|1236,1244|false|false|false|||feverish
Finding|Sign or Symptom|SIMPLE_SEGMENT|1236,1244|false|false|false|C0015967|Fever|feverish
Event|Event|SIMPLE_SEGMENT|1249,1255|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1249,1255|false|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1261,1267|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1261,1267|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1261,1267|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1261,1280|false|false|false|C0027498|Nausea and vomiting|nausea and vomiting
Event|Event|SIMPLE_SEGMENT|1272,1280|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|1272,1280|false|false|false|C0042963|Vomiting|vomiting
Drug|Substance|SIMPLE_SEGMENT|1302,1308|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|1302,1308|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|1302,1308|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1302,1308|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Antibiotic|SIMPLE_SEGMENT|1320,1331|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|1320,1331|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|1340,1348|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|1340,1348|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|1340,1348|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|SIMPLE_SEGMENT|1349,1357|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|1368,1376|false|false|false|||admitted
Finding|Functional Concept|SIMPLE_SEGMENT|1384,1391|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1384,1391|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1384,1391|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1384,1391|false|false|false|C0199168|Medical service|medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1384,1399|false|false|false|C0199168;C0587569|Medical service;Physician service|medical service
Event|Event|SIMPLE_SEGMENT|1392,1399|false|false|false|||service
Event|Occupational Activity|SIMPLE_SEGMENT|1392,1399|false|false|false|C0557854|Services|service
Finding|Idea or Concept|SIMPLE_SEGMENT|1392,1399|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|SIMPLE_SEGMENT|1412,1422|false|false|false|||evaluation
Finding|Idea or Concept|SIMPLE_SEGMENT|1412,1422|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|1412,1422|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Intellectual Product|SIMPLE_SEGMENT|1412,1437|false|false|false|C1317348|Evaluation and management note|evaluation and management
Procedure|Health Care Activity|SIMPLE_SEGMENT|1412,1437|false|false|false|C2945623|Evaluation and Management|evaluation and management
Event|Event|SIMPLE_SEGMENT|1427,1437|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|1427,1437|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|1427,1437|false|false|false|C0376636|Disease Management|management
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1446,1451|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|SIMPLE_SEGMENT|1456,1463|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1456,1463|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1456,1463|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|1464,1471|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1481,1490|false|false|false|||continues
Event|Event|SIMPLE_SEGMENT|1510,1516|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1510,1516|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1523,1528|false|false|false|||feels
Event|Event|SIMPLE_SEGMENT|1538,1546|false|false|false|||nauseous
Finding|Sign or Symptom|SIMPLE_SEGMENT|1538,1546|false|false|false|C0027497|Nausea|nauseous
Event|Event|SIMPLE_SEGMENT|1553,1559|true|false|false|||denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1564,1573|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1564,1578|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1574,1578|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1574,1578|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1574,1578|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1574,1578|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1595,1602|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1615,1622|false|false|false|||feeling
Finding|Mental Process|SIMPLE_SEGMENT|1615,1622|false|false|false|C1527305|Feelings|feeling
Event|Event|SIMPLE_SEGMENT|1624,1630|false|false|false|||better
Finding|Idea or Concept|SIMPLE_SEGMENT|1624,1630|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1678,1683|false|false|false|C1410088|Still|still
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1709,1717|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1709,1717|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1709,1717|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|1724,1731|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|1747,1754|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1747,1754|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1747,1757|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1758,1765|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1758,1771|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|1758,1771|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1758,1782|false|false|false|C0042029;C0262655|Recurrent urinary tract infection;Urinary tract infection|urinary tract infections
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1766,1771|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1772,1782|false|false|false|C0851162|Infection of musculoskeletal system|infections
Event|Event|SIMPLE_SEGMENT|1772,1782|false|false|false|||infections
Finding|Pathologic Function|SIMPLE_SEGMENT|1772,1782|false|false|false|C3714514|Infection|infections
Drug|Organic Chemical|SIMPLE_SEGMENT|1808,1821|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1808,1821|false|false|false|C0008809|ciprofloxacin|ciprofloxacin
Event|Event|SIMPLE_SEGMENT|1808,1821|false|false|false|||ciprofloxacin
Event|Event|SIMPLE_SEGMENT|1836,1843|false|false|false|||reports
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1865,1875|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|1865,1875|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|1865,1875|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Idea or Concept|SIMPLE_SEGMENT|1882,1885|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|1882,1885|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|1886,1892|false|false|false|||course
Finding|Intellectual Product|SIMPLE_SEGMENT|1902,1907|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|1908,1918|true|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|1908,1918|true|false|false|C5441521|Complaint (finding)|complaints
Finding|Finding|SIMPLE_SEGMENT|1923,1943|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1928,1935|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1928,1935|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1928,1935|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1928,1935|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1928,1935|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1928,1943|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1936,1943|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1936,1943|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1936,1943|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1947,1959|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|SIMPLE_SEGMENT|1947,1959|false|false|false|||Hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1969,1972|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1969,1972|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|SIMPLE_SEGMENT|1969,1972|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|SIMPLE_SEGMENT|1969,1972|false|false|false|||lap
Finding|Finding|SIMPLE_SEGMENT|1969,1972|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|SIMPLE_SEGMENT|1969,1972|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1969,1972|false|false|false|C0031150|Laparoscopy|lap
Event|Event|SIMPLE_SEGMENT|1973,1978|false|false|false|||chole
Finding|Functional Concept|SIMPLE_SEGMENT|1988,1992|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1988,1997|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1988,1997|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1993,1997|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1993,1997|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1993,1997|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1993,1997|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1993,2009|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1993,2009|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Event|Event|SIMPLE_SEGMENT|1998,2009|false|false|false|||replacement
Finding|Functional Concept|SIMPLE_SEGMENT|1998,2009|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|SIMPLE_SEGMENT|1998,2009|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1998,2009|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|SIMPLE_SEGMENT|2019,2030|false|false|false|||laminectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2019,2030|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2043,2046|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2043,2046|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|2043,2046|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2056,2063|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2056,2063|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2056,2063|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2056,2070|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder Cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2064,2070|false|false|false|C0006826|Malignant Neoplasms|Cancer
Event|Event|SIMPLE_SEGMENT|2064,2070|false|false|false|||Cancer
Finding|Finding|SIMPLE_SEGMENT|2071,2075|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|2071,2075|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|2071,2075|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|SIMPLE_SEGMENT|2071,2081|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|SIMPLE_SEGMENT|2071,2081|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|SIMPLE_SEGMENT|2076,2081|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|SIMPLE_SEGMENT|2076,2081|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|SIMPLE_SEGMENT|2082,2085|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2082,2085|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2082,2085|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2082,2085|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|SIMPLE_SEGMENT|2082,2085|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2082,2085|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Event|Event|SIMPLE_SEGMENT|2082,2085|false|false|false|||TCC
Event|Event|SIMPLE_SEGMENT|2090,2099|false|false|false|||diagnosed
Finding|Intellectual Product|SIMPLE_SEGMENT|2108,2112|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2118,2124|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2118,2128|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Event|Event|SIMPLE_SEGMENT|2125,2128|false|false|false|||MRI
Finding|Gene or Genome|SIMPLE_SEGMENT|2125,2128|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2125,2128|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|2125,2128|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2131,2139|false|false|false|C1269955|Tumor Cell Invasion|invasion
Event|Event|SIMPLE_SEGMENT|2131,2139|false|false|false|||invasion
Finding|Pathologic Function|SIMPLE_SEGMENT|2131,2139|false|false|false|C2699153|Cell Invasion|invasion
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2145,2152|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2145,2152|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2145,2152|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2145,2157|false|false|false|C0458421|Wall of bladder|bladder wall
Event|Event|SIMPLE_SEGMENT|2159,2170|false|false|false|||perivesical
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2172,2176|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2172,2183|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|2172,2183|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|SIMPLE_SEGMENT|2177,2183|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|SIMPLE_SEGMENT|2177,2183|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2188,2196|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2197,2204|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2197,2204|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|2197,2204|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|2197,2204|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2197,2209|false|false|false|C0447612|Vaginal wall|vaginal wall
Event|Event|SIMPLE_SEGMENT|2211,2212|false|false|false|||/
Event|Event|SIMPLE_SEGMENT|2217,2224|false|false|false|||staging
Finding|Functional Concept|SIMPLE_SEGMENT|2217,2224|false|false|false|C0332305|With staging|staging
Event|Event|SIMPLE_SEGMENT|2234,2246|false|false|false|||hysterectomy
Finding|Finding|SIMPLE_SEGMENT|2234,2246|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2234,2246|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2251,2273|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Event|Event|SIMPLE_SEGMENT|2261,2273|false|false|false|||oophorectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2261,2273|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|SIMPLE_SEGMENT|2278,2283|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|SIMPLE_SEGMENT|2278,2290|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2284,2290|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|SIMPLE_SEGMENT|2284,2290|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2284,2290|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2284,2290|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Event|Event|SIMPLE_SEGMENT|2284,2290|false|false|false|||uterus
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2284,2290|false|false|false|C0869889|examination of uterus|uterus
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2294,2301|false|false|false|C0023267|Fibroid Tumor|fibroid
Event|Event|SIMPLE_SEGMENT|2294,2301|false|false|false|||fibroid
Event|Event|SIMPLE_SEGMENT|2320,2321|false|false|false|||b
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2324,2330|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2324,2341|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|SIMPLE_SEGMENT|2331,2336|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2331,2341|false|false|false|C0024204|lymph nodes|lymph node
Event|Event|SIMPLE_SEGMENT|2342,2351|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2342,2351|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Drug|Chemical Viewed Structurally|SIMPLE_SEGMENT|2359,2366|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2359,2377|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Event|Event|SIMPLE_SEGMENT|2367,2377|false|false|false|||cystectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2367,2377|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2382,2390|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Event|Event|SIMPLE_SEGMENT|2391,2402|false|false|false|||vaginectomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2391,2402|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2408,2415|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|2408,2415|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|SIMPLE_SEGMENT|2408,2415|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|SIMPLE_SEGMENT|2408,2415|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Event|Event|SIMPLE_SEGMENT|2417,2431|false|false|false|||reconstruction
Procedure|Machine Activity|SIMPLE_SEGMENT|2417,2431|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2417,2431|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2437,2442|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2437,2450|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2437,2450|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|SIMPLE_SEGMENT|2451,2459|false|false|false|C1706214|Creation|creation
Event|Event|SIMPLE_SEGMENT|2451,2459|false|false|false|||creation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2451,2459|false|false|false|C0441513|Surgical construction|creation
Event|Event|SIMPLE_SEGMENT|2473,2484|false|false|false|||complicated
Event|Event|SIMPLE_SEGMENT|2488,2498|false|false|false|||bacteremia
Finding|Finding|SIMPLE_SEGMENT|2488,2498|false|false|false|C0004610|Bacteremia|bacteremia
Event|Event|SIMPLE_SEGMENT|2503,2514|true|false|false|||development
Finding|Functional Concept|SIMPLE_SEGMENT|2503,2514|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|SIMPLE_SEGMENT|2503,2514|true|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Event|Event|SIMPLE_SEGMENT|2518,2533|true|false|false|||intra-abdominal
Finding|Functional Concept|SIMPLE_SEGMENT|2518,2533|true|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|SIMPLE_SEGMENT|2535,2540|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|2535,2540|true|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|2541,2551|true|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|2541,2551|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|2541,2551|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|2541,2551|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|2541,2551|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|SIMPLE_SEGMENT|2560,2565|true|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|SIMPLE_SEGMENT|2560,2565|true|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2560,2575|true|false|false|C3495845|Drain placement|drain placement
Event|Event|SIMPLE_SEGMENT|2566,2575|true|false|false|||placement
Procedure|Health Care Activity|SIMPLE_SEGMENT|2566,2575|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2566,2575|true|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Event|Event|SIMPLE_SEGMENT|2593,2594|true|false|false|||/
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2600,2603|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2600,2603|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2600,2603|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|2600,2603|true|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|2624,2639|true|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|2624,2639|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|2624,2639|true|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2624,2639|true|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Functional Concept|SIMPLE_SEGMENT|2644,2650|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2644,2658|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2651,2658|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2651,2658|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2651,2658|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2651,2658|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2664,2670|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2664,2670|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2664,2670|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2664,2670|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2664,2678|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2671,2678|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2671,2678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2671,2678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2671,2678|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|SIMPLE_SEGMENT|2680,2688|false|false|false|||Negative
Finding|Classification|SIMPLE_SEGMENT|2680,2688|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|SIMPLE_SEGMENT|2680,2688|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2680,2688|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|SIMPLE_SEGMENT|2680,2692|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2693,2700|true|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2693,2700|true|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|2693,2700|true|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2693,2700|true|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2693,2703|true|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Event|Event|SIMPLE_SEGMENT|2708,2716|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2708,2716|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2708,2716|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2708,2716|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2708,2721|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2708,2721|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2717,2721|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2717,2721|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2717,2721|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2723,2732|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|2733,2737|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|2733,2737|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2733,2737|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|2740,2746|false|false|false|||VITALS
Event|Event|SIMPLE_SEGMENT|2757,2761|false|false|false|||Temp
Finding|Gene or Genome|SIMPLE_SEGMENT|2757,2761|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2757,2761|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|SIMPLE_SEGMENT|2811,2819|false|false|false|||delivery
Finding|Finding|SIMPLE_SEGMENT|2811,2819|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|SIMPLE_SEGMENT|2811,2819|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|SIMPLE_SEGMENT|2811,2819|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2811,2819|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|SIMPLE_SEGMENT|2824,2831|false|false|false|||Dyspnea
Finding|Finding|SIMPLE_SEGMENT|2824,2831|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2824,2831|false|false|false|C0013404;C2024878|Dyspnea|Dyspnea
Event|Event|SIMPLE_SEGMENT|2835,2839|false|false|false|||RASS
Finding|Intellectual Product|SIMPLE_SEGMENT|2835,2839|false|false|false|C5419117|Richmond Agitation-Sedation Scale Clinical Classification|RASS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2843,2847|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|2843,2847|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2843,2847|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|2843,2853|false|false|false|C0582148|Pain score|Pain Score
Event|Event|SIMPLE_SEGMENT|2848,2853|false|false|false|||Score
Finding|Finding|SIMPLE_SEGMENT|2848,2853|false|false|false|C0449820|Score|Score
Event|Event|SIMPLE_SEGMENT|2860,2867|false|false|false|||GENERAL
Finding|Classification|SIMPLE_SEGMENT|2860,2867|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2860,2867|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2869,2874|true|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|2869,2874|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2869,2874|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|2869,2874|true|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|2869,2874|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|2869,2874|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|2869,2874|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Idea or Concept|SIMPLE_SEGMENT|2885,2893|true|false|false|C0750489|apparent|apparent
Event|Event|SIMPLE_SEGMENT|2894,2902|true|false|false|||distress
Finding|Finding|SIMPLE_SEGMENT|2894,2902|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|SIMPLE_SEGMENT|2894,2902|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2904,2910|true|false|false|C0015450|Face|facial
Event|Event|SIMPLE_SEGMENT|2911,2919|true|false|false|||twitches
Finding|Finding|SIMPLE_SEGMENT|2911,2919|true|false|false|C0231530|Muscle twitch|twitches
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2920,2924|true|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2920,2924|true|false|false|C5848506||EYES
Event|Event|SIMPLE_SEGMENT|2926,2935|false|false|false|||Anicteric
Finding|Finding|SIMPLE_SEGMENT|2926,2935|false|false|false|C0205180|Anicteric|Anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2937,2943|false|false|false|C0034121|Pupil|pupils
Event|Event|SIMPLE_SEGMENT|2952,2957|false|false|false|||round
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2958,2961|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2958,2961|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|SIMPLE_SEGMENT|2958,2961|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|SIMPLE_SEGMENT|2958,2961|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2963,2967|true|false|false|C0013443;C0521421|Ear structure|Ears
Finding|Gene or Genome|SIMPLE_SEGMENT|2963,2967|true|false|false|C1414437|EPRS1 gene|Ears
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2993,3001|true|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|2993,3001|true|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|3003,3009|true|false|false|||masses
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3014,3020|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|3014,3020|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|3014,3020|true|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3023,3033|true|false|false|C0521367|Oropharyngeal|Oropharynx
Finding|Finding|SIMPLE_SEGMENT|3042,3056|true|false|false|C0221198|Lesion|visible lesion
Event|Event|SIMPLE_SEGMENT|3050,3056|true|false|false|||lesion
Finding|Finding|SIMPLE_SEGMENT|3050,3056|true|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|SIMPLE_SEGMENT|3050,3056|true|false|false|C0221198;C1546698|Lesion|lesion
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3058,3066|true|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|3058,3066|true|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|3070,3077|true|false|false|||exudate
Finding|Body Substance|SIMPLE_SEGMENT|3070,3077|true|false|false|C0015388;C1546629|Exudate|exudate
Finding|Intellectual Product|SIMPLE_SEGMENT|3070,3077|true|false|false|C0015388;C1546629|Exudate|exudate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3082,3087|true|false|false|C0018787;C4037974|Chest>Heart;Heart|Heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3082,3087|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|Heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|3082,3087|true|false|false|C0795691|HEART PROBLEM|Heart
Finding|Finding|SIMPLE_SEGMENT|3082,3095|true|false|false|C0425586|Heart regular|Heart regular
Event|Event|SIMPLE_SEGMENT|3088,3095|true|false|false|||regular
Event|Event|SIMPLE_SEGMENT|3100,3106|true|false|false|||murmur
Finding|Finding|SIMPLE_SEGMENT|3100,3106|true|false|false|C0018808|Heart murmur|murmur
Event|Event|SIMPLE_SEGMENT|3126,3129|true|false|false|||JVD
Finding|Finding|SIMPLE_SEGMENT|3126,3129|true|false|false|C0425687|Jugular venous engorgement|JVD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3131,3135|false|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3131,3135|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Event|Event|SIMPLE_SEGMENT|3131,3135|false|false|false|||RESP
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3137,3142|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|3143,3148|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|3143,3148|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|3152,3164|false|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3152,3164|false|false|false|C0004339|Auscultation|auscultation
Finding|Idea or Concept|SIMPLE_SEGMENT|3170,3174|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3175,3178|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3175,3178|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3175,3178|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|3175,3178|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3175,3178|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3175,3178|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3175,3187|false|false|false|C0001868|Air Movements|air movement
Event|Event|SIMPLE_SEGMENT|3179,3187|false|false|false|||movement
Finding|Organism Function|SIMPLE_SEGMENT|3179,3187|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3202,3211|false|false|false|C5885990||Breathing
Event|Event|SIMPLE_SEGMENT|3202,3211|false|false|false|||Breathing
Finding|Finding|SIMPLE_SEGMENT|3202,3211|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|Breathing
Finding|Organism Function|SIMPLE_SEGMENT|3202,3211|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|Breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|3202,3211|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|Breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|3202,3211|false|false|false|C1160636|respiratory system process|Breathing
Event|Event|SIMPLE_SEGMENT|3215,3226|false|false|false|||non-labored
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3231,3238|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3231,3238|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|SIMPLE_SEGMENT|3231,3238|false|false|false|C0941288|Abdomen problem|Abdomen
Finding|Finding|SIMPLE_SEGMENT|3231,3243|false|false|false|C0426663|Abdomen soft|Abdomen soft
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3239,3243|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|3239,3243|false|false|false|||soft
Event|Event|SIMPLE_SEGMENT|3260,3270|false|false|false|||non-tender
Event|Event|SIMPLE_SEGMENT|3274,3283|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3274,3283|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3286,3291|false|false|false|C0021853|Intestines|Bowel
Event|Event|SIMPLE_SEGMENT|3292,3298|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3292,3298|false|false|false|C0037709||sounds
Event|Event|SIMPLE_SEGMENT|3299,3306|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|3299,3306|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|3299,3306|false|false|false|C0150312;C0449450|Present;Presentation|present
Event|Event|SIMPLE_SEGMENT|3312,3315|true|false|false|||HSM
Finding|Gene or Genome|SIMPLE_SEGMENT|3312,3315|true|false|false|C1537594|LRRC4B gene|HSM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3323,3333|true|false|false|C1550314|Suprapubic|suprapubic
Event|Event|SIMPLE_SEGMENT|3334,3342|true|false|false|||fullness
Event|Event|SIMPLE_SEGMENT|3346,3356|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3346,3356|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3346,3356|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|3360,3369|true|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3360,3369|true|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|3371,3376|false|false|false|||foley
Event|Event|SIMPLE_SEGMENT|3377,3385|false|false|false|||catheter
Finding|Intellectual Product|SIMPLE_SEGMENT|3377,3385|false|false|false|C1546572||catheter
Event|Activity|SIMPLE_SEGMENT|3389,3394|false|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3389,3394|false|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3389,3394|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3389,3394|false|false|false|C1533810||place
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3395,3398|false|false|false|C0022681|Medullary sponge kidney|MSK
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3395,3398|false|false|false|C0022681|Medullary sponge kidney|MSK
Event|Event|SIMPLE_SEGMENT|3395,3398|false|false|false|||MSK
Finding|Gene or Genome|SIMPLE_SEGMENT|3395,3398|false|false|false|C1420279|SIK1 gene|MSK
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3400,3404|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3400,3404|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|3400,3404|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Finding|SIMPLE_SEGMENT|3400,3411|false|false|false|C2230237|Supple neck|Neck supple
Event|Event|SIMPLE_SEGMENT|3405,3411|false|false|false|||supple
Finding|Functional Concept|SIMPLE_SEGMENT|3405,3411|false|false|false|C0332254|Supple|supple
Event|Event|SIMPLE_SEGMENT|3413,3418|false|false|false|||moves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3419,3434|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3423,3434|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|3436,3444|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3436,3444|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3453,3457|false|false|false|||full
Event|Event|SIMPLE_SEGMENT|3462,3471|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3462,3471|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3462,3471|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3487,3496|false|false|false|C3687203|All limbs|all limbs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3491,3496|false|false|false|C0015385|Limb structure|limbs
Anatomy|Body System|SIMPLE_SEGMENT|3497,3501|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3497,3501|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3497,3501|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3497,3501|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3497,3501|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3497,3501|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|3506,3512|true|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3506,3512|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|SIMPLE_SEGMENT|3516,3527|true|false|false|||ulcerations
Finding|Pathologic Function|SIMPLE_SEGMENT|3516,3527|true|false|false|C0041582|Ulcer|ulcerations
Event|Event|SIMPLE_SEGMENT|3528,3533|true|false|false|||noted
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3541,3546|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3541,3546|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3541,3546|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|3541,3546|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|3541,3546|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|3541,3546|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3541,3546|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|3548,3556|false|false|false|||oriented
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3558,3562|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3558,3562|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|SIMPLE_SEGMENT|3558,3562|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|SIMPLE_SEGMENT|3563,3572|false|false|false|||symmetric
Finding|Conceptual Entity|SIMPLE_SEGMENT|3563,3572|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3563,3572|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|SIMPLE_SEGMENT|3574,3578|false|false|false|C0553544|Gaze|gaze
Drug|Immunologic Factor|SIMPLE_SEGMENT|3579,3588|false|false|false|C0301869|Immunostimulating conjugate (antigen)|conjugate
Event|Event|SIMPLE_SEGMENT|3579,3588|false|false|false|||conjugate
Event|Event|SIMPLE_SEGMENT|3595,3599|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|3601,3607|false|false|false|||speech
Finding|Organism Function|SIMPLE_SEGMENT|3601,3607|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3601,3607|false|false|false|C0846595|Speech assessment|speech
Event|Event|SIMPLE_SEGMENT|3616,3621|false|false|false|||moves
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3622,3631|false|false|false|C3687203|All limbs|all limbs
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3626,3631|false|false|false|C0015385|Limb structure|limbs
Event|Event|SIMPLE_SEGMENT|3633,3642|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|3633,3642|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3633,3642|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3633,3642|false|false|false|C2229507|sensory exam|sensation
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3646,3651|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3646,3651|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|3646,3651|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|3646,3651|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|3646,3651|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3646,3651|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3646,3651|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|SIMPLE_SEGMENT|3646,3657|false|false|false|C0423553|Light touch|light touch
Event|Event|SIMPLE_SEGMENT|3652,3657|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|3652,3657|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3652,3657|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3652,3657|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|SIMPLE_SEGMENT|3666,3672|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3666,3672|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3684,3689|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|PSYCH
Event|Event|SIMPLE_SEGMENT|3684,3689|false|false|false|||PSYCH
Event|Event|SIMPLE_SEGMENT|3691,3699|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|3691,3699|false|false|false|C2987187|Pleasant|pleasant
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|3701,3719|false|false|false|C0233462|Appropriate affect|appropriate affect
Event|Event|SIMPLE_SEGMENT|3713,3719|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|3713,3719|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|3713,3719|false|false|false|C2237113|assessment of affect|affect
Finding|Body Substance|SIMPLE_SEGMENT|3721,3730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3721,3730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3721,3730|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3721,3730|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|3731,3735|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|3731,3735|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3731,3735|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|3738,3742|false|false|false|||AVSS
Event|Event|SIMPLE_SEGMENT|3744,3754|false|false|false|||ambulating
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3770,3778|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|3770,3778|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|3770,3778|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|3780,3788|true|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3780,3788|true|false|false|C0856443|Urostomy procedure|Urostomy
Event|Event|SIMPLE_SEGMENT|3789,3792|true|false|false|||bag
Finding|Intellectual Product|SIMPLE_SEGMENT|3789,3792|true|false|false|C1552710|Bag Data Type|bag
Event|Activity|SIMPLE_SEGMENT|3796,3801|true|false|false|C1882509|put - instruction imperative|place
Event|Event|SIMPLE_SEGMENT|3796,3801|true|false|false|||place
Finding|Functional Concept|SIMPLE_SEGMENT|3796,3801|true|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|SIMPLE_SEGMENT|3796,3801|true|false|false|C1533810||place
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3820,3828|true|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|3820,3828|true|false|false|||erythema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3832,3836|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3832,3836|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3832,3836|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3832,3836|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3859,3869|false|false|false|C2598148||LABORATORY
Event|Event|SIMPLE_SEGMENT|3859,3869|false|false|false|||LABORATORY
Finding|Functional Concept|SIMPLE_SEGMENT|3859,3869|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|LABORATORY
Finding|Intellectual Product|SIMPLE_SEGMENT|3859,3869|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|LABORATORY
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3859,3869|false|false|false|C4283904|Laboratory observation|LABORATORY
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3859,3877|false|false|false|C1254595|Laboratory Results|LABORATORY RESULTS
Event|Event|SIMPLE_SEGMENT|3870,3877|false|false|false|||RESULTS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3892,3897|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3892,3897|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3892,3897|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3898,3901|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3908,3911|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3908,3911|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3908,3911|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3918,3921|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3918,3921|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3918,3921|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3918,3921|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3927,3930|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3927,3930|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3938,3941|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3938,3941|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3938,3941|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3938,3941|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3938,3941|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3946,3949|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3946,3949|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3946,3949|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3946,3949|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3946,3949|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3946,3949|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3955,3959|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3955,3959|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3987,3990|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4007,4012|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4007,4012|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4007,4012|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4013,4016|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4023,4026|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4023,4026|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4023,4026|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4033,4036|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4033,4036|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4033,4036|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4033,4036|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4043,4046|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4043,4046|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4054,4057|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4054,4057|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4054,4057|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4054,4057|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4054,4057|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4061,4064|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4061,4064|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4061,4064|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4061,4064|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4061,4064|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4061,4064|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4070,4074|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4070,4074|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4102,4105|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4122,4127|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4122,4127|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4122,4127|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4128,4131|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4137,4140|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4137,4140|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4137,4140|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4147,4150|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4147,4150|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4147,4150|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4147,4150|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4157,4160|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4157,4160|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4168,4171|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4168,4171|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4168,4171|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4168,4171|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4168,4171|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4175,4178|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4175,4178|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4175,4178|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4175,4178|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4175,4178|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4175,4178|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4184,4188|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4184,4188|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4216,4219|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4236,4241|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4236,4241|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4236,4241|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4236,4249|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4236,4249|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4236,4249|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4242,4249|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4242,4249|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4242,4249|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4242,4249|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4242,4249|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4242,4249|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4297,4301|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4297,4301|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4297,4301|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4326,4331|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4326,4331|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4326,4331|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4326,4339|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4326,4339|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4326,4339|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4332,4339|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4332,4339|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4332,4339|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4332,4339|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4332,4339|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4332,4339|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4385,4389|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4385,4389|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4385,4389|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4414,4419|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4414,4419|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4414,4419|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4414,4427|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4420,4427|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4420,4427|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4420,4427|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4420,4427|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4420,4427|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|4420,4427|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4420,4427|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4420,4427|false|false|false|C0201925|Calcium measurement|Calcium
Event|Event|SIMPLE_SEGMENT|4450,4462|false|false|false|||MICROBIOLOGY
Finding|Functional Concept|SIMPLE_SEGMENT|4450,4462|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|4450,4462|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4450,4462|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|SIMPLE_SEGMENT|4477,4482|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|4477,4482|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|4477,4482|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4487,4491|false|false|false|C1515974|Anatomic Site|Site
Finding|Intellectual Product|SIMPLE_SEGMENT|4487,4491|false|false|false|C1546778||Site
Event|Event|SIMPLE_SEGMENT|4493,4503|false|false|false|||CYSTOSCOPY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4493,4503|false|false|false|C0010702|Cystoscopy|CYSTOSCOPY
Finding|Functional Concept|SIMPLE_SEGMENT|4509,4514|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4509,4521|false|false|false|C0227613|Right kidney|RIGHT KIDNEY
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4515,4521|false|false|false|C0022646;C0227665|Both kidneys;Kidney|KIDNEY
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4515,4521|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|KIDNEY
Event|Event|SIMPLE_SEGMENT|4515,4521|false|false|false|||KIDNEY
Finding|Sign or Symptom|SIMPLE_SEGMENT|4515,4521|false|false|false|C0812426|Kidney problem|KIDNEY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4515,4521|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4515,4521|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4523,4527|false|false|false|C1883550|Wash Dosage Form|WASH
Event|Activity|SIMPLE_SEGMENT|4523,4527|false|false|false|C0441648|Wash (cleansing action)|WASH
Event|Event|SIMPLE_SEGMENT|4523,4527|false|false|false|||WASH
Finding|Functional Concept|SIMPLE_SEGMENT|4523,4527|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|WASH
Finding|Gene or Genome|SIMPLE_SEGMENT|4523,4527|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|WASH
Finding|Intellectual Product|SIMPLE_SEGMENT|4523,4527|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|WASH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4523,4527|false|false|false|C2699154|Cell Wash|WASH
Finding|Idea or Concept|SIMPLE_SEGMENT|4561,4566|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|SIMPLE_SEGMENT|4561,4573|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4567,4573|false|false|false|C4255046||REPORT
Event|Event|SIMPLE_SEGMENT|4567,4573|false|false|false|||REPORT
Finding|Intellectual Product|SIMPLE_SEGMENT|4567,4573|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|SIMPLE_SEGMENT|4567,4573|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|SIMPLE_SEGMENT|4582,4587|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|SIMPLE_SEGMENT|4582,4587|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|SIMPLE_SEGMENT|4582,4587|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4582,4595|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4588,4595|false|false|false|C1706355|Culture Dose Form|CULTURE
Event|Event|SIMPLE_SEGMENT|4588,4595|false|false|false|||CULTURE
Finding|Functional Concept|SIMPLE_SEGMENT|4588,4595|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|SIMPLE_SEGMENT|4588,4595|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4588,4595|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Event|Event|SIMPLE_SEGMENT|4597,4602|false|false|false|||Final
Finding|Idea or Concept|SIMPLE_SEGMENT|4597,4602|false|false|false|C1546485|Diagnosis Type - Final|Final
Event|Event|SIMPLE_SEGMENT|4628,4635|false|false|false|||FAECIUM
Event|Event|SIMPLE_SEGMENT|4648,4651|false|false|false|||CFU
Event|Activity|SIMPLE_SEGMENT|4676,4684|false|false|false|C1272683||REQUESTS
Event|Event|SIMPLE_SEGMENT|4676,4684|false|false|false|||REQUESTS
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4685,4699|false|false|false|C0012655|Disease susceptibility|SUSCEPTIBILITY
Finding|Functional Concept|SIMPLE_SEGMENT|4685,4699|false|false|false|C1264642|Susceptibility (property) (qualifier value)|SUSCEPTIBILITY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4685,4707|false|false|false|C0806957|Microbial susceptibility tests|SUSCEPTIBILITY TESTING
Event|Event|SIMPLE_SEGMENT|4700,4707|false|false|false|||TESTING
Finding|Functional Concept|SIMPLE_SEGMENT|4700,4707|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TESTING
Finding|Intellectual Product|SIMPLE_SEGMENT|4700,4707|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|TESTING
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4721,4735|false|false|false|C0374989|Unspecified Staphylococcus infection in conditions classified elsewhere and of unspecified site|STAPHYLOCOCCUS
Event|Event|SIMPLE_SEGMENT|4721,4735|false|false|false|||STAPHYLOCOCCUS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4737,4746|false|false|false|C0009118|Coagulase|COAGULASE
Drug|Enzyme|SIMPLE_SEGMENT|4737,4746|false|false|false|C0009118|Coagulase|COAGULASE
Event|Event|SIMPLE_SEGMENT|4747,4755|false|false|false|||NEGATIVE
Finding|Classification|SIMPLE_SEGMENT|4747,4755|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Finding|Finding|SIMPLE_SEGMENT|4747,4755|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|NEGATIVE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4747,4755|false|false|false|C5237010|Expression Negative|NEGATIVE
Event|Event|SIMPLE_SEGMENT|4776,4779|false|false|false|||CFU
Event|Event|SIMPLE_SEGMENT|4807,4814|false|false|false|||SPECIES
Finding|Classification|SIMPLE_SEGMENT|4807,4814|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|SPECIES
Finding|Idea or Concept|SIMPLE_SEGMENT|4807,4814|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|SPECIES
Event|Event|SIMPLE_SEGMENT|4850,4853|false|false|false|||CFU
Event|Event|SIMPLE_SEGMENT|4890,4903|false|false|false|||SENSITIVITIES
Finding|Finding|SIMPLE_SEGMENT|4890,4903|false|false|false|C0427965|Antimicrobial susceptibility|SENSITIVITIES
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4905,4908|false|false|false|C2732473|Ductal Carcinoma In Situ with Microinvasion|MIC
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4905,4908|false|false|false|C0066256|methyl isocyanate|MIC
Drug|Organic Chemical|SIMPLE_SEGMENT|4905,4908|false|false|false|C0066256|methyl isocyanate|MIC
Event|Event|SIMPLE_SEGMENT|4905,4908|false|false|false|||MIC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4905,4908|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4905,4908|false|false|false|C0281162;C0427978|Minimum Inhibitory Concentration Test;cisplatin/ifosfamide/mitomycin protocol|MIC
Event|Event|SIMPLE_SEGMENT|4923,4926|false|false|false|||MCG
Drug|Antibiotic|SIMPLE_SEGMENT|5095,5105|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5095,5105|false|false|false|C0002680;C2095775|ampicillin;ampicillins|AMPICILLIN
Drug|Organic Chemical|SIMPLE_SEGMENT|5126,5140|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5126,5140|false|false|false|C0028156|nitrofurantoin|NITROFURANTOIN
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5157,5169|false|false|false|C0481114|Tetracyclines causing adverse effects in therapeutic use|TETRACYCLINE
Drug|Antibiotic|SIMPLE_SEGMENT|5157,5169|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Drug|Organic Chemical|SIMPLE_SEGMENT|5157,5169|false|false|false|C0039644;C1744619|Tetracycline Antibiotics;tetracycline|TETRACYCLINE
Event|Event|SIMPLE_SEGMENT|5157,5169|false|false|false|||TETRACYCLINE
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5188,5198|false|false|false|C0042313|vancomycin|VANCOMYCIN
Drug|Antibiotic|SIMPLE_SEGMENT|5188,5198|false|false|false|C0042313|vancomycin|VANCOMYCIN
Event|Event|SIMPLE_SEGMENT|5188,5198|false|false|false|||VANCOMYCIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5188,5198|false|false|false|C0489941|Vancomycin measurement|VANCOMYCIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5220,5225|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|5220,5225|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|5220,5225|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5220,5234|false|true|false|C0200949|Blood culture|Blood cultures
Event|Event|SIMPLE_SEGMENT|5226,5234|false|false|false|||cultures
Finding|Idea or Concept|SIMPLE_SEGMENT|5226,5234|false|false|false|C0010453|Culture (Anthropological)|cultures
Event|Event|SIMPLE_SEGMENT|5235,5239|false|false|false|||NGTD
Finding|Intellectual Product|SIMPLE_SEGMENT|5242,5247|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5248,5256|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5248,5263|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5248,5263|false|false|false|C0489547|Hospital course|Hospital Course
Event|Event|SIMPLE_SEGMENT|5277,5285|false|false|false|||admitted
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5291,5297|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|5291,5297|false|false|false|||sepsis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5305,5312|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5305,5318|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|5305,5318|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5313,5318|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5320,5329|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5320,5329|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5320,5329|false|false|false|C3714514|Infection|infection
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5346,5354|false|false|false|C4019011|Exchange (clinical)|exchange
Event|Event|SIMPLE_SEGMENT|5346,5354|false|false|false|||exchange
Finding|Social Behavior|SIMPLE_SEGMENT|5346,5354|false|false|false|C0678640|degree of relationship - exchange|exchange
Event|Event|SIMPLE_SEGMENT|5364,5370|false|false|false|||placed
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5387,5397|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|5387,5397|false|false|false|C0042313|vancomycin|vancomycin
Event|Event|SIMPLE_SEGMENT|5387,5397|false|false|false|||vancomycin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5387,5397|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Antibiotic|SIMPLE_SEGMENT|5402,5410|false|false|false|C0055003|cefepime|cefepime
Drug|Organic Chemical|SIMPLE_SEGMENT|5402,5410|false|false|false|C0055003|cefepime|cefepime
Event|Event|SIMPLE_SEGMENT|5402,5410|false|false|false|||cefepime
Event|Event|SIMPLE_SEGMENT|5412,5420|false|false|false|||narrowed
Drug|Antibiotic|SIMPLE_SEGMENT|5429,5440|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|5429,5440|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|5467,5474|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|5467,5474|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5467,5474|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|5467,5474|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|5467,5477|false|false|false|C0262926|Medical History|history of
Finding|Functional Concept|SIMPLE_SEGMENT|5478,5487|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Finding|Idea or Concept|SIMPLE_SEGMENT|5478,5487|false|false|false|C0332325;C1550464|Resistant (qualifier value);resistant - Observation Interpretation Susceptibility|resistant
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5478,5487|false|false|false|C2827757|Antimicrobial Resistance Result|resistant
Event|Event|SIMPLE_SEGMENT|5488,5497|false|false|false|||organisms
Event|Event|SIMPLE_SEGMENT|5512,5520|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|5526,5531|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|5526,5531|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|5526,5531|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|5526,5531|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|5549,5558|false|false|false|||sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|5549,5558|false|false|false|C0332324|Sensitive|sensitive
Finding|Functional Concept|SIMPLE_SEGMENT|5549,5561|false|false|false|C0332324|Sensitive|sensitive to
Drug|Antibiotic|SIMPLE_SEGMENT|5563,5573|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|5563,5573|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|5563,5573|false|false|false|||ampicillin
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5588,5592|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5593,5597|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5593,5597|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|5593,5597|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|5593,5597|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|5593,5597|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|5602,5608|false|false|false|||placed
Drug|Organic Chemical|SIMPLE_SEGMENT|5624,5632|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5624,5632|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|5624,5632|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|5624,5632|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|5624,5632|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|5624,5632|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Antibiotic|SIMPLE_SEGMENT|5652,5662|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|5652,5662|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|5652,5662|false|false|false|||ampicillin
Finding|Functional Concept|SIMPLE_SEGMENT|5669,5680|false|false|false|C0231242|Complicated|complicated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5681,5688|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5690,5695|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5696,5705|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|5696,5705|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|5696,5705|false|false|false|C3714514|Infection|infection
Finding|Functional Concept|SIMPLE_SEGMENT|5707,5717|false|false|false|C1524062|Additional|additional
Finding|Finding|SIMPLE_SEGMENT|5707,5721|false|false|false|C4534574|Additional day|additional day
Finding|Idea or Concept|SIMPLE_SEGMENT|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5738,5744|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|5768,5778|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|5768,5778|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5768,5778|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|5789,5793|false|false|false|||stop
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5798,5810|false|false|false|C0355642|Drugs used in migraine prophylaxis|prophylactic
Event|Event|SIMPLE_SEGMENT|5798,5810|false|false|false|||prophylactic
Finding|Functional Concept|SIMPLE_SEGMENT|5798,5810|false|false|false|C0445202|Prophylactic behavior|prophylactic
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5811,5814|false|false|false|C0149552|Structure of temporal pole|TMP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5811,5814|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Antibiotic|SIMPLE_SEGMENT|5811,5814|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5811,5814|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5811,5814|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Organic Chemical|SIMPLE_SEGMENT|5811,5814|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Event|Event|SIMPLE_SEGMENT|5811,5814|false|false|false|||TMP
Finding|Gene or Genome|SIMPLE_SEGMENT|5811,5814|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Finding|Intellectual Product|SIMPLE_SEGMENT|5811,5814|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Finding|Receptor|SIMPLE_SEGMENT|5811,5814|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Drug|Antibiotic|SIMPLE_SEGMENT|5825,5835|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|5825,5835|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|5825,5835|false|false|false|||ampicillin
Finding|Intellectual Product|SIMPLE_SEGMENT|5841,5845|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|5846,5852|false|false|false|||resume
Event|Event|SIMPLE_SEGMENT|5859,5868|false|false|false|||finishing
Event|Event|SIMPLE_SEGMENT|5873,5879|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|5883,5893|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|5883,5893|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|5883,5893|false|false|false|||ampicillin
Finding|Functional Concept|SIMPLE_SEGMENT|5909,5919|false|false|false|C1524062|Additional|additional
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5935,5938|false|false|false|C0149552|Structure of temporal pole|TMP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5935,5938|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Antibiotic|SIMPLE_SEGMENT|5935,5938|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5935,5938|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|5935,5938|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Drug|Organic Chemical|SIMPLE_SEGMENT|5935,5938|false|false|false|C0040079;C0041041;C0384479;C1259382|EMP1 protein, human;Thymidine Monophosphate;epithelial membrane protein-1;trimethoprim|TMP
Event|Event|SIMPLE_SEGMENT|5935,5938|false|false|false|||TMP
Finding|Gene or Genome|SIMPLE_SEGMENT|5935,5938|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Finding|Intellectual Product|SIMPLE_SEGMENT|5935,5938|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Finding|Receptor|SIMPLE_SEGMENT|5935,5938|false|false|false|C0384479;C0812384;C1259382;C1706000;C5420102|AML Transfusion Medicine Procedures Table;EMP1 gene;EMP1 protein, human;EMP1 wt Allele, Human;epithelial membrane protein-1|TMP
Event|Event|SIMPLE_SEGMENT|5956,5959|false|false|false|||ppx
Finding|Gene or Genome|SIMPLE_SEGMENT|5956,5959|false|false|false|C1418850|PPP4C gene|ppx
Drug|Antibiotic|SIMPLE_SEGMENT|5966,5976|false|false|false|C0003232|Antibiotics|antibiotic
Event|Event|SIMPLE_SEGMENT|5977,5983|false|false|false|||course
Event|Event|SIMPLE_SEGMENT|5986,5992|false|false|false|||follow
Finding|Functional Concept|SIMPLE_SEGMENT|5986,5992|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5986,5992|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|5986,5995|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|SIMPLE_SEGMENT|5986,5995|false|false|false|C1522577|follow-up|follow up
Event|Event|SIMPLE_SEGMENT|5993,5995|false|false|false|||up
Event|Event|SIMPLE_SEGMENT|6014,6022|false|false|false|||problems
Finding|Idea or Concept|SIMPLE_SEGMENT|6014,6022|false|false|false|C1546466|Problems - What subject filter|problems
Event|Event|SIMPLE_SEGMENT|6023,6032|false|false|false|||addressed
Event|Event|SIMPLE_SEGMENT|6038,6053|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|6038,6053|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Finding|SIMPLE_SEGMENT|6094,6100|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|6094,6100|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6101,6109|false|false|false|C1550297|Prerenal|prerenal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6120,6126|false|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|SIMPLE_SEGMENT|6120,6126|false|false|false|||sepsis
Drug|Substance|SIMPLE_SEGMENT|6144,6150|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|6144,6150|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|6144,6150|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6144,6150|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Antibiotic|SIMPLE_SEGMENT|6155,6166|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|6155,6166|false|false|false|||antibiotics
Finding|Idea or Concept|SIMPLE_SEGMENT|6170,6175|false|false|false|C1552828|Table Frame - above|above
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6186,6196|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|6186,6196|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|6186,6196|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|6186,6196|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6186,6196|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|6202,6209|false|false|false|||trended
Drug|Organic Chemical|SIMPLE_SEGMENT|6211,6219|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6211,6219|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|6211,6219|false|false|false|||Losartan
Event|Event|SIMPLE_SEGMENT|6234,6238|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|6245,6254|false|false|false|||restarted
Event|Event|SIMPLE_SEGMENT|6258,6267|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6258,6267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6258,6267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6258,6267|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6258,6267|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6273,6287|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|6273,6287|false|false|false|||Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|6273,6287|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Event|Event|SIMPLE_SEGMENT|6289,6298|false|false|false|||continued
Drug|Organic Chemical|SIMPLE_SEGMENT|6299,6311|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6299,6311|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|SIMPLE_SEGMENT|6299,6311|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6328,6342|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Event|Event|SIMPLE_SEGMENT|6328,6342|false|false|false|||Hypothyroidism
Event|Event|SIMPLE_SEGMENT|6344,6352|false|false|false|||continue
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6353,6366|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6353,6366|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6353,6366|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6353,6366|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Event|Event|SIMPLE_SEGMENT|6353,6366|false|false|false|||levothyroxine
Event|Event|SIMPLE_SEGMENT|6404,6413|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6404,6413|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6404,6413|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6404,6413|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6404,6413|false|false|false|C0030685|Patient Discharge|discharge
Event|Activity|SIMPLE_SEGMENT|6414,6424|false|false|false|C0441655|Activities|activities
Event|Event|SIMPLE_SEGMENT|6414,6424|false|false|false|||activities
Finding|Finding|SIMPLE_SEGMENT|6414,6424|false|false|false|C2239122|activities (history)|activities
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6429,6440|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6429,6440|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|6429,6440|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6429,6440|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|6429,6453|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|6444,6453|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6444,6453|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6472,6482|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6472,6482|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|6472,6487|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|6483,6487|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|6483,6487|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|6491,6499|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|6504,6512|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6504,6512|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|6504,6512|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|6504,6512|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|6504,6512|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|6504,6512|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|6517,6530|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6517,6530|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|6517,6530|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6517,6530|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|6545,6548|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6549,6553|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|6549,6553|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|6549,6553|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6549,6553|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|SIMPLE_SEGMENT|6556,6560|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|SIMPLE_SEGMENT|6561,6566|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|6561,6566|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|SIMPLE_SEGMENT|6571,6583|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6571,6583|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|6601,6615|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6601,6615|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|6601,6615|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Organic Chemical|SIMPLE_SEGMENT|6638,6646|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6638,6646|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|6638,6646|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|6638,6653|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6638,6653|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6647,6653|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6647,6653|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6647,6653|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|6647,6653|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6647,6653|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6647,6653|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6664,6667|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6664,6667|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6664,6667|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6664,6667|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6664,6667|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6672,6685|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6672,6685|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6672,6685|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6672,6685|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6672,6692|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|6672,6692|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6672,6692|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6686,6692|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6686,6692|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6686,6692|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|6686,6692|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6686,6692|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6686,6692|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|6714,6723|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6714,6723|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|6739,6742|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6743,6750|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|6743,6750|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|6743,6750|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|SIMPLE_SEGMENT|6755,6763|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6755,6763|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|6755,6763|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|6755,6773|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6755,6773|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6764,6773|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6764,6773|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|6764,6773|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6764,6773|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6764,6773|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|6764,6773|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|6764,6773|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6764,6773|false|false|false|C0202194|Potassium measurement|Potassium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6783,6786|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6783,6786|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6783,6786|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|6783,6786|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6783,6786|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6791,6804|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6791,6804|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|6791,6804|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|6791,6804|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6807,6810|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|6807,6810|false|false|false|||TAB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6824,6836|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|6824,6836|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|6824,6836|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|6824,6843|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6824,6843|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6837,6843|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|6837,6843|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|SIMPLE_SEGMENT|6837,6843|false|false|false|||Glycol
Finding|Gene or Genome|SIMPLE_SEGMENT|6858,6861|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|6862,6874|false|false|false|||Constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|6862,6874|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6884,6888|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|6884,6888|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|6884,6888|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|6884,6888|false|false|false|C1546701|line source specimen code|Line
Drug|Antibiotic|SIMPLE_SEGMENT|6894,6906|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|SIMPLE_SEGMENT|6894,6906|false|false|false|C0041041|trimethoprim|Trimethoprim
Event|Event|SIMPLE_SEGMENT|6926,6935|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6926,6935|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6926,6935|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6926,6935|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6926,6935|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6926,6947|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6936,6947|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6936,6947|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|6936,6947|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6936,6947|false|false|false|C4284232|Medications|Medications
Drug|Antibiotic|SIMPLE_SEGMENT|6953,6963|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|6953,6963|false|false|false|C0002680;C2095775|ampicillin;ampicillins|Ampicillin
Drug|Antibiotic|SIMPLE_SEGMENT|6983,6993|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|6983,6993|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Antibiotic|SIMPLE_SEGMENT|6983,7000|false|false|false|C0282052|ampicillin sodium|ampicillin sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|6983,7000|false|false|false|C0282052|ampicillin sodium|ampicillin sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6994,7000|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6994,7000|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6994,7000|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|6994,7000|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6994,7000|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6994,7000|false|false|false|C0337443|Sodium measurement|sodium
Finding|Intellectual Product|SIMPLE_SEGMENT|7018,7023|false|false|false|C1720374|Every - dosing instruction fragment|Every
Event|Activity|SIMPLE_SEGMENT|7036,7040|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|7036,7040|false|false|false|C2828567|PRSS30P gene|Disp
Event|Event|SIMPLE_SEGMENT|7052,7059|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7052,7059|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|SIMPLE_SEGMENT|7067,7077|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|7067,7077|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Antibiotic|SIMPLE_SEGMENT|7067,7084|false|false|false|C0282052|ampicillin sodium|ampicillin sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|7067,7084|false|false|false|C0282052|ampicillin sodium|ampicillin sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7078,7084|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7078,7084|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7078,7084|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|7078,7084|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7078,7084|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7078,7084|false|false|false|C0337443|Sodium measurement|sodium
Finding|Intellectual Product|SIMPLE_SEGMENT|7102,7107|false|false|false|C1720374|Every - dosing instruction fragment|Every
Event|Activity|SIMPLE_SEGMENT|7120,7124|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|7120,7124|false|false|false|C2828567|PRSS30P gene|Disp
Event|Event|SIMPLE_SEGMENT|7136,7143|false|false|false|||Refills
Finding|Idea or Concept|SIMPLE_SEGMENT|7136,7143|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|7152,7165|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7152,7165|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|7152,7165|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7152,7165|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|7180,7183|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7184,7188|false|false|false|C2598155||Pain
Event|Event|SIMPLE_SEGMENT|7184,7188|false|false|false|||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|7184,7188|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7184,7188|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|SIMPLE_SEGMENT|7191,7195|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|SIMPLE_SEGMENT|7196,7201|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|7196,7201|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|SIMPLE_SEGMENT|7208,7220|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7208,7220|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|SIMPLE_SEGMENT|7240,7254|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7240,7254|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|SIMPLE_SEGMENT|7240,7254|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Organic Chemical|SIMPLE_SEGMENT|7279,7287|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7279,7287|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|7279,7287|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|7279,7294|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7279,7294|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7288,7294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7288,7294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7288,7294|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7288,7294|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7288,7294|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7288,7294|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7305,7308|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7305,7308|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7305,7308|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7305,7308|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7305,7308|false|false|false|C1332410|BID gene|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7315,7328|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|7315,7328|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|7315,7328|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7315,7328|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7315,7335|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|SIMPLE_SEGMENT|7315,7335|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7315,7335|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7329,7335|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7329,7335|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7329,7335|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|7329,7335|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|7329,7335|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7329,7335|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|SIMPLE_SEGMENT|7359,7368|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7359,7368|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|SIMPLE_SEGMENT|7384,7387|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7388,7395|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|7388,7395|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|7388,7395|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|SIMPLE_SEGMENT|7402,7410|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7402,7410|false|false|false|C0126174|losartan|Losartan
Event|Event|SIMPLE_SEGMENT|7402,7410|false|false|false|||Losartan
Drug|Organic Chemical|SIMPLE_SEGMENT|7402,7420|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7402,7420|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7411,7420|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7411,7420|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|SIMPLE_SEGMENT|7411,7420|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|7411,7420|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7411,7420|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|SIMPLE_SEGMENT|7411,7420|false|false|false|||Potassium
Finding|Physiologic Function|SIMPLE_SEGMENT|7411,7420|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7411,7420|false|false|false|C0202194|Potassium measurement|Potassium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|7430,7433|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7430,7433|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7430,7433|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|7430,7433|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|7430,7433|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|7440,7453|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7440,7453|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|7440,7453|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|7440,7453|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7456,7459|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|7456,7459|false|false|false|||TAB
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7476,7488|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|7476,7488|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|7476,7488|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|7476,7495|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7476,7495|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7489,7495|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|7489,7495|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|SIMPLE_SEGMENT|7489,7495|false|false|false|||Glycol
Finding|Gene or Genome|SIMPLE_SEGMENT|7510,7513|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|7514,7526|false|false|false|||Constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7514,7526|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7536,7540|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|7536,7540|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|SIMPLE_SEGMENT|7536,7540|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|SIMPLE_SEGMENT|7536,7540|false|false|false|C1546701|line source specimen code|Line
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7547,7551|false|false|false|C0675390|ARID1A protein, human|HELD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7547,7551|false|false|false|C0675390|ARID1A protein, human|HELD
Event|Event|SIMPLE_SEGMENT|7547,7551|false|false|false|||HELD
Finding|Gene or Genome|SIMPLE_SEGMENT|7547,7551|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Finding|Idea or Concept|SIMPLE_SEGMENT|7547,7551|false|false|false|C1948036;C2985160|ARID1A wt Allele;Held - activity status|HELD
Drug|Antibiotic|SIMPLE_SEGMENT|7553,7565|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|SIMPLE_SEGMENT|7553,7565|false|false|false|C0041041|trimethoprim|Trimethoprim
Event|Event|SIMPLE_SEGMENT|7553,7565|false|false|false|||Trimethoprim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7587,7597|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|7587,7597|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7587,7597|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|7602,7606|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|7616,7623|true|false|false|||restart
Drug|Antibiotic|SIMPLE_SEGMENT|7624,7636|true|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|SIMPLE_SEGMENT|7624,7636|true|false|false|C0041041|trimethoprim|Trimethoprim
Event|Event|SIMPLE_SEGMENT|7624,7636|true|false|false|||Trimethoprim
Event|Event|SIMPLE_SEGMENT|7653,7659|true|false|false|||finish
Drug|Antibiotic|SIMPLE_SEGMENT|7666,7676|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|7666,7676|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|7666,7676|false|false|false|||ampicillin
Event|Event|SIMPLE_SEGMENT|7681,7690|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7681,7690|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7681,7690|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7681,7690|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7681,7690|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7681,7702|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|7681,7702|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7691,7702|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|7691,7702|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|7691,7702|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|7704,7712|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|7704,7712|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|7704,7717|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|7713,7717|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|7713,7717|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|7713,7717|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|7713,7717|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|7720,7728|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|7720,7728|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|7736,7745|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7736,7745|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7736,7745|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7736,7745|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7736,7745|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|7736,7755|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7746,7755|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|7746,7755|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7746,7755|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7746,7755|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7746,7755|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7757,7768|false|false|false|C0231242|Complicated|Complicated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7780,7783|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7780,7783|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7780,7783|false|false|false|C0077906|urinastatin|UTI
Event|Event|SIMPLE_SEGMENT|7780,7783|false|false|false|||UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|7780,7783|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Event|Event|SIMPLE_SEGMENT|7787,7796|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7787,7796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7787,7796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7787,7796|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7787,7796|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7797,7806|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7797,7806|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|7797,7806|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|7797,7806|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|7808,7814|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7808,7821|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|7808,7821|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7815,7821|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7815,7821|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|7823,7828|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|7823,7828|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|7833,7841|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|7833,7841|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|7843,7848|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7843,7865|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7843,7865|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|7852,7865|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|7852,7865|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|7852,7865|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7867,7872|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|7867,7872|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7867,7872|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|7867,7872|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|7867,7872|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7867,7872|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|7867,7872|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|7877,7888|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|7877,7888|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|7890,7898|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7890,7898|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|7890,7898|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7899,7905|false|false|false|C5889824||Status
Event|Event|SIMPLE_SEGMENT|7899,7905|false|false|false|||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7899,7905|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|7907,7917|false|false|false|||Ambulatory
Finding|Functional Concept|SIMPLE_SEGMENT|7907,7917|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|7907,7917|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|7907,7917|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|7907,7917|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|SIMPLE_SEGMENT|7920,7931|false|false|false|||Independent
Finding|Finding|SIMPLE_SEGMENT|7920,7931|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|7920,7931|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|SIMPLE_SEGMENT|7935,7944|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|7935,7944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7935,7944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7935,7944|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7935,7944|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7935,7957|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7935,7957|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|7935,7957|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7945,7957|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|7945,7957|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7945,7957|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|7968,7976|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|7984,7992|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|8003,8012|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|8013,8019|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|8013,8019|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|8025,8031|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|8025,8031|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|8042,8051|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|8052,8058|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|8052,8058|false|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|8063,8069|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|8063,8069|false|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|8080,8085|false|false|false|||stent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8087,8095|false|false|false|C4019011|Exchange (clinical)|exchange
Event|Event|SIMPLE_SEGMENT|8087,8095|false|false|false|||exchange
Finding|Social Behavior|SIMPLE_SEGMENT|8087,8095|false|false|false|C0678640|degree of relationship - exchange|exchange
Event|Event|SIMPLE_SEGMENT|8102,8107|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|8102,8107|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|8102,8107|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|8102,8107|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|8108,8112|false|false|false|||grew
Finding|Classification|SIMPLE_SEGMENT|8130,8137|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|species
Finding|Idea or Concept|SIMPLE_SEGMENT|8130,8137|false|false|false|C1548151;C1705920|Species;Species - Nature of Abnormal Testing|species
Event|Event|SIMPLE_SEGMENT|8145,8151|false|false|false|||source
Finding|Finding|SIMPLE_SEGMENT|8145,8151|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|SIMPLE_SEGMENT|8145,8151|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|SIMPLE_SEGMENT|8145,8151|false|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8161,8170|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|8161,8170|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|8161,8170|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|8187,8199|false|false|false|||enterococcus
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8203,8207|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8208,8212|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|8208,8212|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|SIMPLE_SEGMENT|8208,8212|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Event|Event|SIMPLE_SEGMENT|8208,8212|false|false|false|||line
Finding|Intellectual Product|SIMPLE_SEGMENT|8208,8212|false|false|false|C1546701|line source specimen code|line
Event|Event|SIMPLE_SEGMENT|8218,8224|false|false|false|||placed
Event|Event|SIMPLE_SEGMENT|8238,8244|false|false|false|||finish
Finding|Idea or Concept|SIMPLE_SEGMENT|8256,8259|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|8256,8259|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|8260,8266|false|false|false|||course
Drug|Antibiotic|SIMPLE_SEGMENT|8274,8284|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Drug|Organic Chemical|SIMPLE_SEGMENT|8274,8284|false|false|false|C0002680;C2095775|ampicillin;ampicillins|ampicillin
Event|Event|SIMPLE_SEGMENT|8274,8284|false|false|false|||ampicillin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8300,8306|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8300,8306|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|8300,8306|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8300,8306|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8300,8306|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8300,8313|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|8307,8313|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|SIMPLE_SEGMENT|8307,8313|false|false|false|||injury
Event|Event|SIMPLE_SEGMENT|8315,8321|false|false|false|||likely
Finding|Finding|SIMPLE_SEGMENT|8315,8321|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|8315,8321|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8327,8336|false|true|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|8327,8336|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|8327,8336|false|true|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|8343,8351|false|false|false|||resolved
Drug|Antibiotic|SIMPLE_SEGMENT|8358,8369|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|8358,8369|false|false|false|||antibiotics
Drug|Substance|SIMPLE_SEGMENT|8374,8380|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|8374,8380|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|8374,8380|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8374,8380|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|8391,8399|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|8391,8399|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|8391,8399|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|8407,8411|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|8407,8411|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|8407,8411|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8407,8411|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|8407,8414|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|SIMPLE_SEGMENT|8423,8431|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8432,8444|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|8432,8444|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8432,8444|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

