CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Level of Care - Surgery|Finding|false|false||SURGERY
null|Surgical procedure finding|Finding|false|false||SURGERY
null|Surgical aspects|Finding|false|false||SURGERYnull|Operative Surgical Procedures|Procedure|false|false||SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|Corgard|Drug|false|false||Corgard
null|Corgard|Drug|false|false||Corgardnull|Vasotec|Drug|false|false||Vasotec
null|Vasotec|Drug|false|false||Vasotecnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Irreducible inguinal hernia|Disorder|false|false|C0018246|incarcerated inguinal hernianull|In prison (finding)|Finding|false|false|C0018246|incarceratednull|Hernia, Inguinal|Disorder|false|false|C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0019294;C0401074;C0019270;C0392751|inguinalnull|Hernia|Disorder|false|false|C0018246|hernianull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Left inguinal hernia|Disorder|false|false|C0018246|Left inguinal hernianull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Repair of inguinal hernia|Procedure|false|false|C0018246|inguinal hernia repairnull|Hernia, Inguinal|Disorder|false|false|C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0043240;C4319951;C0019270;C0019294;C0262537;C0021446;C0019328;C0374711;C1705181|inguinalnull|Herniorrhaphy|Procedure|false|false|C0018246|hernia repairnull|Hernia|Disorder|false|false|C0018246|hernianull|Repair|Finding|false|false|C0018246|repair
null|Wound Healing|Finding|false|false|C0018246|repairnull|Repair - Remedial Action|Procedure|false|false|C0018246|repair
null|Surgical repair|Procedure|false|false|C0018246|repairnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|Atrial Fibrillation|Disorder|false|false||afibnull|Atrial Fibrillation by ECG Finding|Lab|false|false||afibnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|carotid disease|Disorder|false|false|C0007272|carotid diseasenull|Carotid Arteries|Anatomy|false|false|C0741975|carotidnull|Disease|Disorder|false|false||diseasenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Pulmonary Emphysema|Disorder|false|false||emphysemanull|Pathological accumulation of air in tissues|Finding|false|false||emphysemanull|Recent|Time|false|false||recentnull|Pneumonia|Disorder|false|false||pneumonianull|Visit Priority Code - Elective|Finding|false|false||elective
null|Act Priority - elective|Finding|false|false||elective
null|Admission Type - Elective|Finding|false|false||electivenull|elective|Time|false|false||electivenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Repair of inguinal hernia|Procedure|false|false|C0018246|inguinal hernia repairnull|Hernia, Inguinal|Disorder|false|false|C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0019270;C0019328;C0043240;C4319951;C0019294;C0021446;C0374711;C1705181|inguinalnull|Herniorrhaphy|Procedure|false|false|C0018246|hernia repairnull|Hernia|Disorder|false|false|C0018246|hernianull|Repair|Finding|false|false|C0018246|repair
null|Wound Healing|Finding|false|false|C0018246|repairnull|Repair - Remedial Action|Procedure|false|false|C0018246|repair
null|Surgical repair|Procedure|false|false|C0018246|repairnull|LARGE1 wt Allele|Finding|false|false||large
null|LARGE1 gene|Finding|false|false||largenull|Large|LabModifier|false|false||largenull|In prison (finding)|Finding|false|false||incarceratednull|Malignant neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|sigmoid colon
null|Benign neoplasm of sigmoid colon|Disorder|false|false|C0009368;C4071907;C0227391;C0227391|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0750873;C0009373;C0154061;C0496907;C0496864;C0153436|sigmoid colonnull|Sigmoid colon|Anatomy|false|false|C0496864;C0153436|sigmoidnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false|C0009368;C4071907;C0227391|colon
null|Colonic Diseases|Disorder|false|false|C0009368;C4071907;C0227391|colon
null|Carcinoma in situ of colon|Disorder|false|false|C0009368;C4071907;C0227391|colonnull|COLON PROBLEM|Finding|false|false|C0227391;C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009373;C0154061;C0496907;C0496864;C0153436;C0750873|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009373;C0154061;C0496907;C0496864;C0153436;C0750873|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Bilateral|Modifier|false|false||BILATERALnull|Moderate - Severity of Illness Code|Finding|false|false||MODERATE
null|Moderate|Finding|false|false||MODERATEnull|Moderate (severity modifier)|Modifier|false|false||MODERATE
null|Moderate - Allergy Severity|Modifier|false|false||MODERATE
null|Moderation|Modifier|false|false||MODERATEnull|carotid disease|Disorder|false|false|C0007272|CAROTID DISEASEnull|Carotid Arteries|Anatomy|false|false|C0741975;C0012634|CAROTIDnull|Disease|Disorder|false|false|C0007272|DISEASEnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|CONGESTIVE HEART FAILUREnull|Congestive|Modifier|false|false||CONGESTIVEnull|Congestive heart failure|Disorder|false|false|C4037974;C0018787|HEART FAILURE
null|Heart failure|Disorder|false|false|C4037974;C0018787|HEART FAILUREnull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEART
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|HEARTnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|HEARTnull|Chest>Heart|Anatomy|false|false|C0680095;C0231174;C5200924;C0018801;C0018802;C0018802;C0795691;C0153957;C0153500|HEART
null|Heart|Anatomy|false|false|C0680095;C0231174;C5200924;C0018801;C0018802;C0018802;C0795691;C0153957;C0153500|HEARTnull|Failure (biologic function)|Finding|false|false|C4037974;C0018787|FAILURE
null|Failure|Finding|false|false|C4037974;C0018787|FAILURE
null|Personal failure|Finding|false|false|C4037974;C0018787|FAILUREnull|Coronary Artery Disease|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|CORONARY ARTERY DISEASE
null|Coronary Arteriosclerosis|Disorder|false|false|C0205042;C0018787;C0226004;C0003842|CORONARY ARTERY DISEASEnull|Coronary artery|Anatomy|false|false|C1956346;C0010054;C0012634;C0852949|CORONARY ARTERYnull|Heart|Anatomy|false|false|C0012634;C0852949;C1956346;C0010054|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Arteriopathic disease|Disorder|false|false|C0018787;C0226004;C0003842;C0205042|ARTERY DISEASEnull|Arterial system|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|ARTERY
null|Arteries|Anatomy|false|false|C0852949;C1956346;C0010054;C0012634|ARTERYnull|Disease|Disorder|false|false|C0018787;C0205042;C0226004;C0003842|DISEASEnull|Gastroesophageal reflux disease|Disorder|false|false|C0744316|GASTROESOPHAGEAL REFLUXnull|Infantile Gastroesophageal Reflux|Finding|false|false|C0744316|GASTROESOPHAGEAL REFLUX
null|Acid reflux|Finding|false|false|C0744316|GASTROESOPHAGEAL REFLUXnull|gastroesophageal|Anatomy|false|false|C3813607;C4317146;C0232483;C0017168|GASTROESOPHAGEALnull|Reflux|Finding|false|false|C0744316|REFLUXnull|Hypertensive disease|Disorder|false|false||HYPERTENSIONnull|Severe - Severity of Illness Code|Finding|false|false||SEVERE
null|Intensity and Distress 5|Finding|false|false||SEVERE
null|Severe - Triage Code|Finding|false|false||SEVERE
null|Severe (severity modifier)|Finding|false|false||SEVERE
null|Allergy Severity - Severe|Finding|false|false||SEVEREnull|Pulmonary Emphysema|Disorder|false|false||EMPHYSEMAnull|Pathological accumulation of air in tissues|Finding|false|false||EMPHYSEMAnull|Pulmonary Hypertension|Finding|false|false|C0024109|PULMONARY HYPERTENSIONnull|Pulmonary (intended site)|Finding|false|false|C0024109|PULMONARYnull|Lung|Anatomy|false|false|C0020542;C4522268;C0020538;C2707265|PULMONARYnull|null|Attribute|false|false|C0024109|PULMONARYnull|Pulmonary (qualifier value)|Modifier|false|false||PULMONARYnull|Hypertensive disease|Disorder|false|false|C0024109|HYPERTENSIONnull|Right bundle branch block|Disorder|false|false|C0225916|RIGHT BUNDLE BRANCH BLOCKnull|null|Finding|false|false|C0225916|RIGHT BUNDLE BRANCH BLOCKnull|Structure of right branch of atrioventricular bundle|Anatomy|false|false|C1552823;C1706085;C1881507;C0085615;C1879286;C0006384;C0344421;C0028778;C0332206;C1533157|RIGHT BUNDLE BRANCHnull|Table Cell Horizontal Align - right|Finding|false|false|C0225916|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Bundle-Branch Block|Disorder|false|false|C0225916|BUNDLE BRANCH BLOCK
null|Hereditary bundle branch system defect|Disorder|false|false|C0225916|BUNDLE BRANCH BLOCKnull|Macromolecular Branch|Drug|false|false|C0225916|BRANCHnull|Branch of|Modifier|false|false||BRANCHnull|Block Dosage Form|Drug|false|false|C0225916|BLOCKnull|Fixed Block|Finding|false|false|C0225916|BLOCK
null|Obstruction|Finding|false|false|C0225916|BLOCK
null|Blocking|Finding|false|false|C0225916|BLOCKnull|Geographic Block|Entity|false|false||BLOCKnull|Block (unit of presentation)|LabModifier|false|false||BLOCK
null|Block Dosing Unit|LabModifier|false|false||BLOCK
null|Block (unit of measure)|LabModifier|false|false||BLOCKnull|Benign Prostatic Hyperplasia|Finding|false|false|C0033572|BENIGN PROSTATIC HYPERTROPHYnull|Benign|Modifier|false|false||BENIGNnull|Prostatic Hypertrophy|Disorder|false|false|C0033572|PROSTATIC HYPERTROPHYnull|Benign Prostatic Hyperplasia|Finding|false|false|C0033572|PROSTATIC HYPERTROPHY
null|Prostatic Hyperplasia|Finding|false|false|C0033572|PROSTATIC HYPERTROPHYnull|Prostate|Anatomy|false|false|C2937421;C1704272;C1704272;C0020564;C1739363|PROSTATICnull|Prostatic|Modifier|false|false||PROSTATICnull|Hypertrophy|Finding|false|false|C0033572|HYPERTROPHYnull|Hyperlipidemia|Disorder|false|false||HYPERLIPIDEMIA
null|Hyperlipoproteinemias|Disorder|false|false||HYPERLIPIDEMIAnull|Serum lipids high (finding)|Finding|false|false||HYPERLIPIDEMIAnull|Paroxysmal atrial fibrillation|Disorder|false|false|C0018792|PAROXYSMAL ATRIAL FIBRILLATIONnull|Paroxysmal|Time|false|false||PAROXYSMALnull|Atrial Fibrillation|Disorder|false|false|C0018792|ATRIAL FIBRILLATIONnull|null|Attribute|false|false|C0018792|ATRIAL FIBRILLATIONnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|ATRIAL FIBRILLATIONnull|Heart Atrium|Anatomy|false|false|C0004238;C0235480;C0232197;C2926591;C0344434|ATRIALnull|Fibrillation|Disorder|false|false|C0018792|FIBRILLATIONnull|History of surgery|Finding|false|false||Past Surgical Historynull|history of prior surgery|Finding|false|false||Surgical Historynull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Electric Countershock|Procedure|false|false||CARDIOVERSIONnull|Structure of right lower lobe of lung|Anatomy|false|false|C3539671;C1428707;C1552823;C2003888;C0023928|RIGHT LOWER LOBEnull|Table Cell Horizontal Align - right|Finding|false|false|C1548802;C1261075;C0225758|RIGHTnull|Right sided|Modifier|false|false||RIGHT
null|Right|Modifier|false|false||RIGHTnull|Structure of lower lobe of lung|Anatomy|false|false|C2003888;C0023928;C3539671;C1428707;C1552823|LOWER LOBEnull|Body Site Modifier - Lower|Anatomy|false|false|C0023928;C1552823;C2003888;C3539671;C1428707|LOWERnull|Lower (action)|Event|false|false|C0225758;C1548802;C1261075|LOWERnull|Lower - spatial qualifier|Modifier|false|false||LOWERnull|AKT1S1 wt Allele|Finding|false|false|C1261075;C0225758;C1548802;C0796494|LOBE
null|AKT1S1 gene|Finding|false|false|C1261075;C0225758;C1548802;C0796494|LOBEnull|lobe|Anatomy|false|false|C0023928;C3539671;C1428707|LOBEnull|Lobectomy|Procedure|false|false|C1548802;C0225758;C0796494;C1261075|LOBECTOMYnull|Coronary Artery Bypass Surgery|Procedure|false|false|C0018787|CORONARY BYPASS SURGERYnull|Coronary Artery Bypass Surgery|Procedure|false|false|C0018787|CORONARY BYPASSnull|Heart|Anatomy|false|false|C0010055;C0543467;C0038895;C1457907;C1547138;C0813207;C0010055;C1536078|CORONARYnull|Coronary|Modifier|false|false||CORONARYnull|Bypass surgery|Procedure|false|false|C0018787|BYPASS SURGERYnull|Creation of shunt|Procedure|false|false|C0018787|BYPASSnull|Level of Care - Surgery|Finding|false|false|C0018787|SURGERY
null|Surgical procedure finding|Finding|false|false|C0018787|SURGERY
null|Surgical aspects|Finding|false|false|C0018787|SURGERYnull|Operative Surgical Procedures|Procedure|false|false|C0018787|SURGERYnull|General surgery specialty|Title|false|false||SURGERY
null|Surgery specialty|Title|false|false||SURGERYnull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Irregular|Modifier|false|false||irregularnull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|cetrimonium bromide|Drug|false|false||CTABnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Tender|Modifier|false|false||tendernull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Surgical wound|Disorder|false|false|C2338258|Incisionnull|Surgical incisions|Procedure|false|false|C2338258|Incisionnull|Cranial incision point|Anatomy|false|false|C1947930;C0332803;C0184898|Incisionnull|Cleaning (activity)|Event|false|false|C2338258|cleannull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Erythema|Disorder|false|false||erythemanull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Irreducible inguinal hernia|Disorder|false|false|C0018246|incarcerated inguinal hernianull|In prison (finding)|Finding|false|false|C0018246|incarceratednull|Hernia, Inguinal|Disorder|false|false|C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0019294;C0401074;C0019270;C0392751|inguinalnull|Hernia|Disorder|false|false|C0018246|hernianull|Details|Modifier|false|false||detailsnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Operative report|Finding|false|false||operative reportnull|Operative|Time|false|false||operativenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Postoperative Period|Time|false|false||postoperativenull|Course|Time|false|false||coursenull|Uncomplicated|Modifier|false|false||uncomplicatednull|BRIEF Health Literacy Screening Tool|Finding|false|false||brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||briefnull|Brief|Time|false|false||briefnull|Shortened|Modifier|false|false||briefnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Regular|Modifier|false|false||regularnull|Breast Feeding|Finding|false|false|C3714591|nursingnull|RNAx nursing therapy actions|Procedure|false|false|C3714591|nursingnull|Discipline of Nursing|Title|false|false||nursingnull|Floor (anatomic)|Anatomy|false|false|C0028678;C0006147|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|IV medication|Drug|false|false||IV medicationnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Issue (document)|Finding|true|false||issue
null|Problem|Finding|true|false||issuenull|Issue (action)|Event|true|false||issuenull|Halls|Drug|false|false||halls
null|Halls|Drug|false|false||hallsnull|Bowel Regimen|Procedure|false|false|C0021853|bowel regimennull|Intestines|Anatomy|false|false|C5979615|bowelnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Flatulence|Finding|false|false||flatusnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Oral medication (substance)|Drug|false|false||oral medicationnull|Oral Medication|Procedure|false|false|C0226896|oral medicationnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C0175795;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Ambulate|Finding|false|false||ambulatenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|amiodarone|Drug|false|false||Amiodarone
null|amiodarone|Drug|false|false||Amiodaronenull|Drug assay amiodarone|Procedure|false|false||Amiodaronenull|Daily|Time|false|false||DAILYnull|apixaban|Drug|false|false||Apixaban
null|apixaban|Drug|false|false||Apixabannull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Daily|Time|false|false||DAILYnull|triamterene|Drug|false|false||Triamterene
null|triamterene|Drug|false|false||Triamterenenull|hydrochlorothiazide|Drug|false|false||HCTZ
null|hydrochlorothiazide|Drug|false|false||HCTZnull|capsule (pharmacologic)|Drug|false|false||CAPnull|CATARACT, ANTERIOR POLAR|Disorder|false|false||CAPnull|BRD4 wt Allele|Finding|false|false||CAP
null|HACD1 gene|Finding|false|false||CAP
null|SERPINB6 gene|Finding|false|false||CAP
null|BRD4 gene|Finding|false|false||CAP
null|CAP1 gene|Finding|false|false||CAP
null|SORBS1 gene|Finding|false|false||CAP
null|LNPEP gene|Finding|false|false||CAPnull|CAP Regimen|Procedure|false|false||CAP
null|cisplatin/cyclophosphamide/doxorubicin protocol|Procedure|false|false||CAP
null|cyclophosphamide/doxorubicin/prednisone protocol|Procedure|false|false||CAPnull|Cap (physical object)|Device|false|false||CAP
null|Syringe Caps|Device|false|false||CAP
null|Cap device|Device|false|false||CAPnull|College of American Pathologists|Subject|false|false||CAPnull|Controlled Attenuation Parameter|Modifier|false|false||CAPnull|Capsule Dosing Unit|LabModifier|false|false||CAPnull|Daily|Time|false|false||DAILYnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|g/24h|LabModifier|false|false||grams per daynull|gram|LabModifier|false|false||gramsnull|per day|Time|false|false||per daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|6 Hours|Time|false|false||6 hoursnull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|4 Hours|Time|false|false||4 hoursnull|Hour|Time|false|false||hoursnull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|sennosides, USP|Drug|false|false||sennosides
null|sennosides, USP|Drug|false|false||sennosidesnull|Evac-U-Gen Reformulated Jan 2008|Drug|false|false||Evac-U-Gen
null|Evac-U-Gen|Drug|false|false||Evac-U-Gen
null|Evac-U-Gen|Drug|false|false||Evac-U-Gen
null|Evac-U-Gen Reformulated Jan 2008|Drug|false|false||Evac-U-Gennull|ECHO protocol|Procedure|false|false||Evacnull|sennosides, USP|Drug|false|false||sennosides
null|sennosides, USP|Drug|false|false||sennosidesnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Align|Drug|false|false||Align
null|Align|Drug|false|false||Alignnull|herbal medicines bifidobacterium infantis|Drug|false|false||bifidobacterium infantisnull|Bifidobacterium longum subspecies infantis|Entity|false|false||bifidobacterium infantis
null|Bifidobacterium infantis|Entity|false|false||bifidobacterium infantisnull|Bifidobacterium|Entity|false|false||bifidobacteriumnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10
null|ubidecarenone|Drug|false|false||coenzyme Q10null|Coenzymes|Drug|false|false||coenzyme
null|Coenzymes|Drug|false|false||coenzymenull|AGO2 wt Allele|Finding|false|false||Q10
null|AGO2 gene|Finding|false|false||Q10null|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|rosuvastatin calcium|Drug|false|false||Rosuvastatin Calcium
null|rosuvastatin calcium|Drug|false|false||Rosuvastatin Calciumnull|rosuvastatin|Drug|false|false||Rosuvastatin
null|rosuvastatin|Drug|false|false||Rosuvastatinnull|calcium|Drug|false|false||Calcium 40
null|calcium|Drug|false|false||Calcium 40
null|calcium|Drug|false|false||Calcium 40null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Hernia, Inguinal|Disorder|false|false|C0018246|Inguinal hernianull|Inguinal region|Anatomy|false|false|C0019294;C0019270|Inguinalnull|Hernia|Disorder|false|false|C0018246|hernianull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Repair|Finding|false|false|C0018246|repair
null|Wound Healing|Finding|false|false|C0018246|repairnull|Repair - Remedial Action|Procedure|false|false|C0018246|repair
null|Surgical repair|Procedure|false|false|C0018246|repairnull|Hernia, Inguinal|Disorder|false|false|C0018246|inguinal hernianull|Inguinal region|Anatomy|false|false|C0019294;C0374711;C1705181;C0019270;C0043240;C4319951|inguinalnull|Hernia|Disorder|false|false|C0018246|hernianull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Recommendation|Finding|false|false||recommendationsnull|Uneventful|Finding|false|false||uneventfulnull|Recovery - healing process|Finding|false|false||recoverynull|null|Event|false|false||recoverynull|recovery - adjustment|LabModifier|false|false||recoverynull|Activity (animal life circumstance)|Finding|false|false||ACTIVITY
null|Physical activity|Finding|false|false||ACTIVITYnull|Activities|Event|false|false||ACTIVITYnull|null|Modifier|false|false||ACTIVITYnull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Prior functioning.stairs|Finding|false|false||stairsnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Distance|LabModifier|false|false||distancesnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Visit|Finding|false|false||visitnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|liquid-based cytology (procedure)|Procedure|false|false||lbsnull|Pounds|LabModifier|false|false||lbsnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Bag Data Type|Finding|false|false||bagnull|null|Device|false|false||bagnull|Bag (unit of presentation)|LabModifier|false|false||bag
null|Bag Dosing Unit|LabModifier|false|false||bagnull|applies to - HL7 Value Set and Coded Concept Property Codes|Finding|false|false||applies tonull|Offspring|Subject|false|false||children
null|Child|Subject|false|false||childrennull|ACP2 protein, human|Drug|false|false||lap
null|ACP2 protein, human|Drug|false|false||lapnull|Congenital laryngeal adductor palsy|Disorder|false|false||lapnull|Left atrial pressure|Finding|false|false||lap
null|ACP2 gene|Finding|false|false||lap
null|PICALM wt Allele|Finding|false|false||lap
null|LAP3 wt Allele|Finding|false|false||lap
null|ACP2 wt Allele|Finding|false|false||lap
null|LAP3 gene|Finding|false|false||lap
null|CENPJ gene|Finding|false|false||lap
null|CEBPB wt Allele|Finding|false|false||lap
null|PICALM gene|Finding|false|false||lap
null|CEBPB gene|Finding|false|false||lapnull|Laparoscopy|Procedure|false|false||lapnull|Lap - unit|LabModifier|false|false||lapnull|Light Exercise|Finding|false|false||light exercisenull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|Feeling comfortable|Finding|false|false||comfortablenull|Bathtub|Device|false|false||bathtubsnull|Swimming Pools|Device|false|false||swimming poolsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|Pool (environment)|Entity|false|false||poolsnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false|C2338258|time
null|Time (foundation metadata concept)|Finding|false|false|C2338258|time
null|Value type - Time|Finding|false|false|C2338258|time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false|C2338258|time
null|Data types - Time|Finding|false|false|C2338258|time
null|null|Finding|false|false|C2338258|timenull|Time|Time|false|false||timenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898;C5575590;C2024467;C1548318;C1547403;C3541383;C5400024|incisionnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|TUB gene|Finding|false|false||tubnull|Tub - container|Device|false|false||tubnull|Tub Dosing Unit|LabModifier|false|false||tubnull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|Heavy (weight) (qualifier value)|Modifier|false|false||Heavy
null|Heavy (amount)|Modifier|false|false||Heavynull|Exercise|Finding|false|false||exercisenull|Exercise Pain Management|Procedure|false|false||exercisenull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Sensory perception|Finding|false|false||sensenull|Slow|Modifier|false|false||slowlynull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Sexual Activity|Finding|false|false||sexual activity
null|Sex Behavior|Finding|false|false||sexual activitynull|Sex Behavior|Finding|false|false||sexualnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Feelings|Finding|false|false||FEELnull|Feel Weak (question)|Finding|false|false||feel weak
null|Weakness|Finding|false|false||feel weaknull|Feel Weak (question)|Finding|false|false||weak
null|Weakness|Finding|false|false||weaknull|Weak|Modifier|false|false||weaknull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Neutrophil Activation Probe Imaging Agent|Drug|false|false||napnull|CTNNBL1 gene|Finding|false|false||nap
null|Napping|Finding|false|false||napnull|Neapolitan Language|Entity|false|false||napnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|LITAF gene|Finding|false|false||Simplenull|Simple|Modifier|false|false||Simplenull|exhaust|Drug|false|false||exhaustnull|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of Phenol|Drug|false|false|C0230069;C3665375;C0031354|sore throat
null|Sore Throat brand of benzocaine & menthol|Drug|false|false|C0230069;C3665375;C0031354|sore throatnull|Pharyngitis|Disorder|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore Throat|Finding|false|false|C0230069;C3665375;C0031354|sore throatnull|Sore to touch|Finding|false|false||sore
null|Sore skin|Finding|false|false||sorenull|Sore sensation quality|Modifier|false|false||sorenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Anterior portion of neck|Anatomy|false|false|C3244654;C0723402;C1550663;C1547926;C0242429;C1950455;C0031350|throat
null|Throat|Anatomy|false|false|C3244654;C0723402;C1550663;C1547926;C0242429;C1950455;C0031350|throat
null|Pharyngeal structure|Anatomy|false|false|C3244654;C0723402;C1550663;C1547926;C0242429;C1950455;C0031350|throatnull|Unspecified tube|Finding|false|false||tube
null|TUBE1 gene|Finding|false|false||tubenull|biomedical tube device|Device|false|false||tube
null|Packaging Tube|Device|false|false||tubenull|tube|Modifier|false|false||tubenull|Tube (unit of presentation)|LabModifier|false|false||tube
null|Tube Dosing Unit|LabModifier|false|false||tubenull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354|throatnull|Throat|Anatomy|false|false|C1550663;C1547926;C0038895;C1457907;C1547138;C0543467;C1950455|throat
null|Anterior portion of neck|Anatomy|false|false|C1550663;C1547926;C0038895;C1457907;C1547138;C0543467;C1950455|throat
null|Pharyngeal structure|Anatomy|false|false|C1550663;C1547926;C0038895;C1457907;C1547138;C0543467;C1950455|throatnull|Intraoperative|Time|false|false||during surgerynull|Level of Care - Surgery|Finding|false|false|C0230069;C3665375;C0031354|surgery
null|Surgical procedure finding|Finding|false|false|C0230069;C3665375;C0031354|surgery
null|Surgical aspects|Finding|false|false|C0230069;C3665375;C0031354|surgerynull|Operative Surgical Procedures|Procedure|false|false|C0230069;C3665375;C0031354|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Somewhat|Finding|false|false||somewhatnull|Depressed mood|Disorder|false|false||depressednull|Poor appetite question|Finding|false|false||poor appetite
null|Decrease in appetite|Finding|false|false||poor appetitenull|null|Attribute|false|false||poor appetitenull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Desire for food|Finding|false|false||appetitenull|Food allergenic extracts|Drug|false|false||Food
null|Food|Drug|false|false||Food
null|Food allergenic extracts|Drug|false|false||Foodnull|Subject's Feelings|Finding|false|false||feelings
null|Feelings|Finding|false|false||feelingsnull|Shortened|Modifier|false|false||shortnull|Short Value|LabModifier|false|false||short
null|Short|LabModifier|false|false||shortnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Surgical wound|Disorder|false|false|C2338258|INCISIONnull|Surgical incisions|Procedure|false|false|C2338258|INCISIONnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|INCISIONnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|Along edge (qualifier value)|Modifier|false|false||edgesnull|Steri-Strip|Device|false|false||steri stripsnull|Silene|Entity|false|false||sterinull|strip medical device|Device|false|false||stripsnull|2 Weeks|Time|false|false||2 weeksnull|week|Time|false|false||weeksnull|Thin (qualifier value)|Modifier|false|false||thinnull|Paper Authorization|Finding|false|false||papernull|Paper|Device|false|false||papernull|Paper Dosing Unit|LabModifier|false|false||papernull|strip medical device|Device|false|false||stripsnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Gently|Modifier|false|false||gentlynull|Materials|Drug|false|false|C2338258|materialnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803;C0520510|incisionnull|Firm|Modifier|false|false||firmnull|Ridging|Finding|false|false|C2338258|ridgenull|crest - location|Modifier|false|false||ridgenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332243;C0332803;C0184898|incisionnull|Direct - PostalAddressUse|Finding|false|false||direct
null|direct address|Finding|false|false||directnull|Direct type of relationship|Modifier|false|false||direct
null|Direct (qualifier)|Modifier|false|false||directnull|Sun Exposure|Phenomenon|false|false||sun exposurenull|Sunlight|Phenomenon|false|false||sunnull|The Sun|Entity|false|false||sun
null|Sundanese language|Entity|false|false||sunnull|Exposure to|Modifier|false|false||exposure tonull|Injury due to exposure to external cause|Disorder|false|false|C2338258|exposurenull|exposure history|Finding|false|false||exposurenull|Accident due to exposure to weather conditions|Phenomenon|false|false||exposurenull|Exposure to|Modifier|false|false||exposurenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0274281;C0332803|incisionnull|Academic Research Enhancement Awards|Event|false|false||areanull|Geographic Locations|Entity|false|false||areanull|Area|Modifier|false|false||areanull|Ointments|Drug|false|false||ointmentsnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Red light (physical force)|Phenomenon|false|false||light rednull|Light Red color|Modifier|false|false||light rednull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|DYRK3 gene|Finding|false|false||red
null|Redness|Finding|false|false||red
null|IK gene|Finding|false|false||rednull|Radiological Exposure Device|Device|false|false||rednull|Red color|Modifier|false|false||rednull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing of skin or wound|Procedure|false|false||dressing
null|Dressing patient (procedure)|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Clothing|Device|false|false||clothesnull|Staining (finding)|Finding|false|false||stainingnull|Staining method|Procedure|false|false||stainingnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Table Frame - above|Finding|false|false||abovenull|Upper|Modifier|false|false||abovenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|TUB gene|Finding|false|false||tubnull|Tub - container|Device|false|false||tubnull|Tub Dosing Unit|LabModifier|false|false||tubnull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|month|Time|false|false||monthsnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Prominent|Modifier|false|false||prominentnull|Intestines|Anatomy|false|false||BOWELSnull|Constipation|Finding|false|false||Constipationnull|Common Specifications in HL7 V3 Publishing|Finding|false|false||common
null|shared attribute|Finding|false|false||commonnull|Common (qualifier value)|LabModifier|false|false||commonnull|Adverse effects|Finding|false|false||side effectnull|Side|Modifier|false|false||sidenull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Percocet|Drug|false|false||Percocet
null|Percocet|Drug|false|false||Percocetnull|codeine|Drug|false|false||codeine
null|codeine|Drug|false|false||codeinenull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Gentle Laxative|Drug|false|false||gentle laxative
null|Gentle Laxative|Drug|false|false||gentle laxativenull|Gentle|Drug|false|false||gentle
null|Gentle|Drug|false|false||gentlenull|Laxatives|Drug|false|false||laxativenull|cow milk allergenic extract|Drug|false|false||milk
null|Milk antigen|Drug|false|false||milk
null|Milk Beverage|Drug|false|false||milk
null|Plant-Based Milk|Drug|false|false||milk
null|cow milk allergenic extract|Drug|false|false||milk
null|Milk Specimen|Drug|false|false||milk
null|Cow's milk|Drug|false|false||milk
null|null|Drug|false|false||milknull|Milk (body substance)|Finding|false|false||milk
null|Milk Specimen Code|Finding|false|false||milknull|magnesium oxide|Drug|false|false||magnesia
null|magnesium oxide|Drug|false|false||magnesianull|Townes syndrome|Disorder|false|false||tbsnull|Toxicity Burden Score|Finding|false|false||tbs
null|SALL1 gene|Finding|false|false||tbs
null|SALL1 wt Allele|Finding|false|false||tbsnull|theta-burst stimulation|Procedure|false|false||tbsnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|prescription document|Finding|true|false||prescriptionnull|Prescription (procedure)|Procedure|true|false||prescriptionnull|Prescription (attribute)|Attribute|true|false||prescriptionnull|48 hours|Time|false|false||48 hoursnull|Hour|Time|false|false||hoursnull|Defecation|Finding|true|false|C0021853|bowel movementnull|Intestines|Anatomy|false|false|C0011135|bowelnull|Movement|Finding|true|false||movementnull|Have Pain|Finding|false|false||have painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Intestines|Anatomy|false|false||bowelsnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|ActInformationPrivacyReason - operations|Finding|false|false||operations
null|HL7PublishingSubSection - operations|Finding|false|false||operations
null|Surgical aspects|Finding|false|false||operationsnull|Operation Activity|Event|false|false||operationsnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|Anti-Diarrhea|Drug|false|false||anti-diarrhea
null|Anti-Diarrhea|Drug|false|false||anti-diarrheanull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Feel Ill Question|Finding|false|false||feel ill
null|Malaise|Finding|false|false||feel ill
null|Feeling bad emotionally|Finding|false|false||feel illnull|Malaise|Finding|false|false||illnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Pain management (procedure)|Procedure|false|false||PAIN MANAGEMENTnull|Pain Management (specialty)|Title|false|false||PAIN MANAGEMENTnull|Administration Method - Pain|Finding|false|false||PAIN
null|Pain|Finding|false|false||PAINnull|null|Attribute|false|false||PAINnull|Disease Management|Procedure|false|false||MANAGEMENTnull|Management Occupations|Subject|false|false||MANAGEMENTnull|Management procedure|Event|false|false||MANAGEMENT
null|Administration occupational activities|Event|false|false||MANAGEMENTnull|Discomfort|Finding|false|false||discomfortnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Abdomen|Anatomy|false|false||abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Often - answer to question|Finding|false|false||oftennull|Frequently|Time|false|false||oftennull|Sore to touch|Finding|false|false||sorenessnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|prescription document|Finding|false|false||prescriptionnull|Prescription (procedure)|Procedure|false|false||prescriptionnull|Prescription (attribute)|Attribute|false|false||prescriptionnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false|C0230028;C0226896|medicinenull|Medicine|Title|false|false||medicinenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C0013227;C1527415|mouth
null|Oral region|Anatomy|false|false|C0013227;C1527415|mouthnull|Important|Modifier|false|false||importantnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|More|LabModifier|false|false||morenull|Frequently|Time|false|false||frequentlynull|More|LabModifier|false|false||morenull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|one time|Finding|false|false||one timenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Observation Interpretation - better|Finding|false|false||betternull|Better|Modifier|false|false||betternull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicine
null|Analgesics|Drug|false|false||pain medicinenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Sharp pain|Finding|false|false||sharp painnull|Sharp sensation quality|Finding|false|false||sharp
null|SPEN wt Allele|Finding|false|false||sharp
null|SPEN gene|Finding|false|false||sharpnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Several|LabModifier|false|false||severalnull|Hour|Time|false|false||hoursnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Nature|Finding|false|false||nature
null|Natures|Finding|false|false||naturenull|Quality|Modifier|false|false||qualitynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||MEDICATIONSnull|Medications|Finding|false|false||MEDICATIONSnull|null|Attribute|false|false||MEDICATIONS
null|null|Attribute|false|false||MEDICATIONSnull|Pharmaceutical Preparations|Drug|false|false||medicinesnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Take|Procedure|false|false||takenull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions