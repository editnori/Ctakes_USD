 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|31,35
No|36,38
:|38,39
_|42,43
_|43,44
_|44,45
<EOL>|45,46
<EOL>|47,48
Admission|48,57
Date|58,62
:|62,63
_|65,66
_|66,67
_|67,68
Discharge|82,91
Date|92,96
:|96,97
_|100,101
_|101,102
_|102,103
<EOL>|103,104
<EOL>|105,106
Date|106,110
of|111,113
Birth|114,119
:|119,120
_|122,123
_|123,124
_|124,125
Sex|138,141
:|141,142
M|145,146
<EOL>|146,147
<EOL>|148,149
Service|149,156
:|156,157
ORTHOPAEDICS|158,170
<EOL>|170,171
<EOL>|172,173
Sulfa|185,190
(|191,192
Sulfonamide|192,203
Antibiotics|204,215
)|215,216
/|217,218
Penicillins|219,230
<EOL>|230,231
<EOL>|232,233
Attending|233,242
:|242,243
_|244,245
_|245,246
_|246,247
.|247,248
<EOL>|248,249
<EOL>|250,251
neck|268,272
pain|273,277
s|278,279
/|279,280
p|280,281
fall|282,286
<EOL>|286,287
<EOL>|288,289
Major|289,294
Surgical|295,303
or|304,306
Invasive|307,315
Procedure|316,325
:|325,326
<EOL>|326,327
None|327,331
on|332,334
this|335,339
Admission|340,349
<EOL>|349,350
<EOL>|351,352
_|380,381
_|381,382
_|382,383
male|384,388
transferred|389,400
from|401,405
outside|406,413
hospital|414,422
for|423,426
<EOL>|427,428
evaluation|428,438
of|439,441
cervical|442,450
_|451,452
_|452,453
_|453,454
fracture|455,463
.|463,464
Today|465,470
the|471,474
patient|475,482
was|483,486
<EOL>|487,488
attempting|488,498
to|499,501
use|502,505
the|506,509
bathroom|510,518
and|519,522
bent|523,527
forward|528,535
and|536,539
fell|540,544
hitting|545,552
<EOL>|553,554
the|554,557
back|558,562
of|563,565
his|566,569
head|570,574
.|574,575
There|576,581
was|582,585
no|586,588
loss|589,593
of|594,596
consciousness|597,610
.|610,611
The|612,615
<EOL>|616,617
patient|617,624
complains|625,634
of|635,637
headache|638,646
and|647,650
neck|651,655
pain|656,660
.|660,661
The|662,665
outside|666,673
<EOL>|674,675
hospital|675,683
the|684,687
patient|688,695
had|696,699
the|700,703
head|704,708
laceration|709,719
stapled|720,727
.|727,728
A|729,730
CT|731,733
scan|734,738
<EOL>|739,740
did|740,743
demonstrate|744,755
the|756,759
fracture|760,768
.|768,769
The|770,773
patient|774,781
denies|782,788
any|789,792
numbness|793,801
,|801,802
<EOL>|803,804
tingling|804,812
in|813,815
his|816,819
arms|820,824
or|825,827
legs|828,832
.|832,833
No|834,836
weakness|837,845
in|846,848
his|849,852
arms|853,857
or|858,860
legs|861,865
.|865,866
<EOL>|867,868
Denies|868,874
any|875,878
bowel|879,884
incontinence|885,897
or|898,900
bladder|901,908
retention|909,918
.|918,919
No|920,922
saddle|923,929
<EOL>|930,931
anesthesia|931,941
.|941,942
Denies|943,949
any|950,953
chest|954,959
pain|960,964
,|964,965
shortness|966,975
of|976,978
breath|979,985
or|986,988
<EOL>|989,990
abdominal|990,999
pain|1000,1004
.|1004,1005
<EOL>|1005,1006
<EOL>|1008,1009
<EOL>|1009,1010
<EOL>|1011,1012
PMH|1034,1037
:|1037,1038
a.|1039,1041
fib|1042,1045
,|1045,1046
colon|1047,1052
ca|1053,1055
,|1055,1056
htn|1057,1060
,|1060,1061
copd|1062,1066
<EOL>|1066,1067
<EOL>|1069,1070
MED|1070,1073
:|1073,1074
warfarin|1075,1083
,|1083,1084
allopurinol|1085,1096
,|1096,1097
asacol|1098,1104
<EOL>|1104,1105
<EOL>|1107,1108
ALL|1108,1111
:|1111,1112
pcn|1113,1116
,|1116,1117
sulfa|1118,1123
<EOL>|1123,1124
<EOL>|1124,1125
<EOL>|1126,1127
:|1141,1142
<EOL>|1142,1143
_|1143,1144
_|1144,1145
_|1145,1146
<EOL>|1146,1147
:|1161,1162
<EOL>|1162,1163
NC|1163,1165
<EOL>|1165,1166
<EOL>|1167,1168
C|1183,1184
collar|1185,1191
in|1192,1194
place|1195,1200
<EOL>|1200,1201
<EOL>|1201,1202
UEC5C6C7C8T1|1202,1214
<EOL>|1214,1215
(|1215,1216
lat|1216,1219
arm|1220,1223
)|1223,1224
(|1226,1227
thumb|1227,1232
)|1232,1233
(|1234,1235
mid|1235,1238
fing|1239,1243
)|1243,1244
(|1245,1246
sm|1246,1248
finger|1249,1255
)|1255,1256
(|1257,1258
med|1258,1261
arm|1262,1265
)|1265,1266
<EOL>|1266,1267
Rintact|1267,1274
intact|1280,1286
intact|1294,1300
intact|1308,1314
intact|1322,1328
<EOL>|1328,1329
Lintact|1329,1336
intact|1342,1348
intact|1356,1362
intact|1370,1376
intact|1384,1390
<EOL>|1390,1391
<EOL>|1391,1392
T2|1392,1394
-|1394,1395
L1|1395,1397
(|1398,1399
Trunk|1399,1404
)|1404,1405
intact|1406,1412
<EOL>|1412,1413
<EOL>|1413,1414
_|1414,1415
_|1415,1416
_|1416,1417
L2|1423,1425
L3|1433,1435
L4|1437,1439
L5S1S2|1441,1447
<EOL>|1447,1448
(|1448,1449
Groin|1449,1454
)|1454,1455
(|1455,1456
Knee|1456,1460
)|1460,1461
(|1465,1466
Med|1466,1469
Calf|1470,1474
)|1474,1475
(|1476,1477
Grt|1477,1480
Toe|1481,1484
)|1484,1485
(|1486,1487
Sm|1487,1489
Toe|1490,1493
)|1493,1494
(|1495,1496
Post|1496,1500
Thigh|1501,1506
)|1506,1507
<EOL>|1507,1508
Rintactintactintactintact|1508,1533
intactintact|1540,1552
<EOL>|1552,1553
Lintactintactintactintact|1553,1578
intactintact|1585,1597
<EOL>|1597,1598
<EOL>|1598,1599
Motor|1599,1604
:|1604,1605
<EOL>|1605,1606
UEDlt|1606,1611
(|1611,1612
C5|1612,1614
)|1614,1615
Bic|1615,1618
(|1618,1619
C6|1619,1621
)|1621,1622
WE|1622,1624
(|1624,1625
C6|1625,1627
)|1627,1628
Tri|1628,1631
(|1631,1632
C7|1632,1634
)|1634,1635
WF|1635,1637
(|1637,1638
C7|1638,1640
)|1640,1641
FF|1641,1643
(|1643,1644
C8|1644,1646
)|1646,1647
FinAbd|1647,1653
(|1653,1654
T1|1654,1656
)|1656,1657
<EOL>|1657,1658
R|1658,1659
5|1662,1663
5|1666,1667
5|1671,1672
5|1676,1677
_|1681,1682
_|1682,1683
_|1683,1684
<EOL>|1684,1685
L|1685,1686
5|1689,1690
5|1693,1694
5|1698,1699
5|1703,1704
_|1708,1709
_|1709,1710
_|1710,1711
<EOL>|1711,1712
<EOL>|1712,1713
_|1713,1714
_|1714,1715
_|1715,1716
Flex|1718,1722
(|1722,1723
L1|1723,1725
)|1725,1726
Add|1727,1730
(|1730,1731
L2|1731,1733
)|1733,1734
Quad|1735,1739
(|1739,1740
L3|1740,1742
)|1742,1743
TA|1745,1747
(|1747,1748
L4|1748,1750
)|1750,1751
_|1752,1753
_|1753,1754
_|1754,1755
_|1756,1757
_|1757,1758
_|1758,1759
<EOL>|1759,1760
R|1760,1761
_|1764,1765
_|1765,1766
_|1766,1767
5|1771,1772
5|1776,1777
5|1781,1782
5|1789,1790
<EOL>|1796,1797
L|1797,1798
_|1801,1802
_|1802,1803
_|1803,1804
5|1808,1809
5|1813,1814
5|1818,1819
5|1823,1824
<EOL>|1824,1825
<EOL>|1825,1826
<EOL>|1839,1840
Babinski|1840,1848
:|1848,1849
negative|1851,1859
<EOL>|1860,1861
Clonus|1861,1867
:|1867,1868
not|1869,1872
present|1873,1880
<EOL>|1880,1881
<EOL>|1883,1884
<EOL>|1884,1885
<EOL>|1886,1887
Patient|1910,1917
was|1918,1921
admitted|1922,1930
to|1931,1933
the|1934,1937
_|1938,1939
_|1939,1940
_|1940,1941
_|1942,1943
_|1943,1944
_|1944,1945
Surgery|1946,1953
Service|1954,1961
for|1962,1965
<EOL>|1966,1967
observation|1967,1978
after|1979,1984
a|1985,1986
C2|1987,1989
fracture|1990,1998
.|1998,1999
TEDs|2001,2005
/|2005,2006
pnemoboots|2006,2016
were|2017,2021
used|2022,2026
for|2027,2030
<EOL>|2031,2032
postoperative|2032,2045
DVT|2046,2049
prophylaxis|2050,2061
.|2061,2062
Diet|2064,2068
was|2069,2072
advanced|2073,2081
as|2082,2084
tolerated|2085,2094
.|2094,2095
<EOL>|2097,2098
The|2098,2101
patient|2102,2109
was|2110,2113
tolerated|2114,2123
oral|2124,2128
pain|2129,2133
medication|2134,2144
.|2144,2145
Physical|2146,2154
therapy|2155,2162
<EOL>|2163,2164
was|2164,2167
consulted|2168,2177
for|2178,2181
mobilization|2182,2194
OOB|2195,2198
to|2199,2201
ambulate|2202,2210
.|2210,2211
He|2213,2215
remained|2216,2224
<EOL>|2225,2226
hypertensive|2226,2238
from|2239,2243
160|2244,2247
-|2248,2249
>|2250,2251
180|2251,2254
.|2254,2255
Medicine|2257,2265
consult|2266,2273
appreciated|2274,2285
-|2286,2287
<EOL>|2288,2289
felt|2289,2293
this|2294,2298
was|2299,2302
long|2303,2307
standing|2308,2316
.|2316,2317
recommended|2319,2330
PRN|2331,2334
antihypertensives|2335,2352
<EOL>|2353,2354
but|2354,2357
cautioned|2358,2367
against|2368,2375
bringing|2376,2384
pressure|2385,2393
too|2394,2397
low|2398,2401
too|2402,2405
quickly|2406,2413
.|2413,2414
<EOL>|2416,2417
Hospital|2417,2425
course|2426,2432
was|2433,2436
otherwise|2437,2446
unremarkable|2447,2459
.|2459,2460
On|2462,2464
the|2465,2468
day|2469,2472
of|2473,2475
<EOL>|2476,2477
discharge|2477,2486
the|2487,2490
patient|2491,2498
was|2499,2502
afebrile|2503,2511
with|2512,2516
stable|2517,2523
vital|2524,2529
signs|2530,2535
,|2535,2536
<EOL>|2537,2538
comfortable|2538,2549
on|2550,2552
oral|2553,2557
pain|2558,2562
control|2563,2570
and|2571,2574
tolerating|2575,2585
a|2586,2587
regular|2588,2595
diet|2596,2600
.|2600,2601
<EOL>|2602,2603
<EOL>|2604,2605
Discharge|2605,2614
Medications|2615,2626
:|2626,2627
<EOL>|2627,2628
1.|2628,2630
Acetaminophen|2631,2644
650|2645,2648
mg|2649,2651
PO|2652,2654
Q4H|2655,2658
:|2658,2659
PRN|2659,2662
pain|2663,2667
,|2667,2668
temp|2669,2673
>|2674,2675
100.5|2675,2680
,|2680,2681
headache|2682,2690
<EOL>|2691,2692
2.|2692,2694
Allopurinol|2695,2706
_|2707,2708
_|2708,2709
_|2709,2710
mg|2711,2713
PO|2714,2716
DAILY|2717,2722
<EOL>|2723,2724
3.|2724,2726
Mesalamine|2727,2737
_|2738,2739
_|2739,2740
_|2740,2741
400|2742,2745
mg|2746,2748
PO|2749,2751
TID|2752,2755
<EOL>|2756,2757
4.|2757,2759
Metoprolol|2760,2770
Tartrate|2771,2779
25|2780,2782
mg|2783,2785
PO|2786,2788
BID|2789,2792
<EOL>|2793,2794
5.|2794,2796
Omeprazole|2797,2807
20|2808,2810
mg|2811,2813
PO|2814,2816
DAILY|2817,2822
<EOL>|2823,2824
6.|2824,2826
Warfarin|2827,2835
1|2836,2837
mg|2838,2840
PO|2841,2843
DAILY|2844,2849
<EOL>|2850,2851
7.|2851,2853
OxycoDONE|2854,2863
(|2864,2865
Immediate|2865,2874
Release|2875,2882
)|2882,2883
2|2885,2886
.|2886,2887
5|2887,2888
-|2888,2889
5|2889,2890
mg|2891,2893
PO|2894,2896
Q4H|2897,2900
:|2900,2901
PRN|2901,2904
pain|2905,2909
<EOL>|2910,2911
8.|2911,2913
Diazepam|2914,2922
2|2923,2924
mg|2925,2927
PO|2928,2930
Q12H|2931,2935
:|2935,2936
PRN|2936,2939
spasms|2940,2946
<EOL>|2947,2948
<EOL>|2948,2949
<EOL>|2950,2951
Discharge|2951,2960
Disposition|2961,2972
:|2972,2973
<EOL>|2973,2974
Home|2974,2978
With|2979,2983
Service|2984,2991
<EOL>|2991,2992
<EOL>|2993,2994
Facility|2994,3002
:|3002,3003
<EOL>|3003,3004
_|3004,3005
_|3005,3006
_|3006,3007
<EOL>|3007,3008
<EOL>|3009,3010
Discharge|3010,3019
Diagnosis|3020,3029
:|3029,3030
<EOL>|3030,3031
C2|3031,3033
fracture|3034,3042
<EOL>|3042,3043
<EOL>|3044,3045
Mental|3066,3072
Status|3073,3079
:|3079,3080
Clear|3081,3086
and|3087,3090
coherent|3091,3099
.|3099,3100
<EOL>|3100,3101
Level|3101,3106
of|3107,3109
Consciousness|3110,3123
:|3123,3124
Alert|3125,3130
and|3131,3134
interactive|3135,3146
.|3146,3147
<EOL>|3147,3148
Activity|3148,3156
Status|3157,3163
:|3163,3164
Ambulatory|3165,3175
-|3176,3177
Independent|3178,3189
.|3189,3190
<EOL>|3190,3191
<EOL>|3192,3193
You|3217,3220
have|3221,3225
undergone|3226,3235
the|3236,3239
following|3240,3249
operation|3250,3259
:|3259,3260
Anterior|3261,3269
Cervical|3270,3278
<EOL>|3279,3280
Decompression|3280,3293
and|3294,3297
Fusion|3298,3304
<EOL>|3304,3305
<EOL>|3305,3306
Immediately|3306,3317
after|3318,3323
the|3324,3327
operation|3328,3337
:|3337,3338
<EOL>|3338,3339
-|3339,3340
Activity|3340,3348
:|3348,3349
You|3350,3353
should|3354,3360
not|3361,3364
lift|3365,3369
anything|3370,3378
greater|3379,3386
than|3387,3391
5|3392,3393
lbs|3394,3397
for|3398,3401
<EOL>|3402,3403
2|3403,3404
weeks|3405,3410
.|3410,3411
You|3412,3415
will|3416,3420
be|3421,3423
more|3424,3428
comfortable|3429,3440
if|3441,3443
you|3444,3447
do|3448,3450
not|3451,3454
sit|3455,3458
in|3459,3461
a|3462,3463
car|3464,3467
<EOL>|3468,3469
or|3469,3471
chair|3472,3477
for|3478,3481
more|3482,3486
than|3487,3491
~|3492,3493
45|3493,3495
minutes|3496,3503
without|3504,3511
getting|3512,3519
up|3520,3522
and|3523,3526
<EOL>|3527,3528
walking|3528,3535
around|3536,3542
.|3542,3543
<EOL>|3543,3544
<EOL>|3544,3545
-|3545,3546
Rehabilitation|3546,3560
/|3560,3561
Physical|3562,3570
Therapy|3571,3578
:|3578,3579
<EOL>|3580,3581
o2|3581,3583
-|3583,3584
3|3584,3585
times|3586,3591
a|3592,3593
day|3594,3597
you|3598,3601
should|3602,3608
go|3609,3611
for|3612,3615
a|3616,3617
walk|3618,3622
for|3623,3626
_|3627,3628
_|3628,3629
_|3629,3630
minutes|3631,3638
as|3639,3641
<EOL>|3642,3643
part|3643,3647
of|3648,3650
your|3651,3655
recovery|3656,3664
.|3664,3665
You|3667,3670
can|3671,3674
walk|3675,3679
as|3680,3682
much|3683,3687
as|3688,3690
you|3691,3694
can|3695,3698
<EOL>|3699,3700
tolerate|3700,3708
.|3708,3709
<EOL>|3711,3712
oIsometric|3712,3722
Extension|3723,3732
Exercise|3733,3741
in|3742,3744
the|3745,3748
collar|3749,3755
:|3755,3756
2x|3757,3759
/|3759,3760
day|3760,3763
x|3764,3765
_|3766,3767
_|3767,3768
_|3768,3769
xercises|3769,3777
as|3778,3780
instructed|3781,3791
.|3791,3792
<EOL>|3792,3793
<EOL>|3793,3794
-|3794,3795
Swallowing|3795,3805
:|3805,3806
Difficulty|3807,3817
swallowing|3818,3828
is|3829,3831
not|3832,3835
uncommon|3836,3844
after|3845,3850
this|3851,3855
<EOL>|3856,3857
type|3857,3861
of|3862,3864
surgery|3865,3872
.|3872,3873
This|3874,3878
should|3879,3885
resolve|3886,3893
over|3894,3898
time|3899,3903
.|3903,3904
Please|3906,3912
take|3913,3917
<EOL>|3918,3919
small|3919,3924
bites|3925,3930
and|3931,3934
eat|3935,3938
slowly|3939,3945
.|3945,3946
Removing|3948,3956
the|3957,3960
collar|3961,3967
while|3968,3973
eating|3974,3980
<EOL>|3981,3982
can|3982,3985
be|3986,3988
helpful|3989,3996
|3997,3998
however|3999,4006
,|4006,4007
please|4008,4014
limit|4015,4020
your|4021,4025
movement|4026,4034
of|4035,4037
your|4038,4042
<EOL>|4043,4044
neck|4044,4048
if|4049,4051
you|4052,4055
remove|4056,4062
your|4063,4067
collar|4068,4074
while|4075,4080
eating|4081,4087
.|4087,4088
<EOL>|4088,4089
<EOL>|4089,4090
-|4090,4091
Cervical|4091,4099
Collar|4100,4106
/|4107,4108
Neck|4109,4113
Brace|4114,4119
:|4119,4120
You|4121,4124
need|4125,4129
to|4130,4132
wear|4133,4137
the|4138,4141
brace|4142,4147
at|4148,4150
<EOL>|4151,4152
all|4152,4155
times|4156,4161
until|4162,4167
your|4168,4172
follow|4173,4179
-|4179,4180
up|4180,4182
appointment|4183,4194
which|4195,4200
should|4201,4207
be|4208,4210
in|4211,4213
2|4214,4215
<EOL>|4216,4217
weeks|4217,4222
.|4222,4223
You|4225,4228
may|4229,4232
remove|4233,4239
the|4240,4243
collar|4244,4250
to|4251,4253
take|4254,4258
a|4259,4260
shower|4261,4267
.|4267,4268
Limit|4270,4275
your|4276,4280
<EOL>|4281,4282
motion|4282,4288
of|4289,4291
your|4292,4296
neck|4297,4301
while|4302,4307
the|4308,4311
collar|4312,4318
is|4319,4321
off|4322,4325
.|4325,4326
Place|4327,4332
the|4333,4336
collar|4337,4343
<EOL>|4344,4345
back|4345,4349
on|4350,4352
your|4353,4357
neck|4358,4362
immediately|4363,4374
after|4375,4380
the|4381,4384
shower|4385,4391
.|4391,4392
<EOL>|4392,4393
<EOL>|4393,4394
-|4394,4395
Wound|4395,4400
Care|4401,4405
:|4405,4406
Monitor|4407,4414
laceration|4415,4425
at|4426,4428
scalp|4429,4434
for|4435,4438
drainage|4439,4447
/|4447,4448
redness|4448,4455
.|4455,4456
<EOL>|4458,4459
Your|4459,4463
PCP|4464,4467
may|4468,4471
take|4472,4476
these|4477,4482
staples|4483,4490
out|4491,4494
.|4494,4495
<EOL>|4495,4496
<EOL>|4496,4497
-|4497,4498
You|4498,4501
should|4502,4508
resume|4509,4515
taking|4516,4522
your|4523,4527
normal|4528,4534
home|4535,4539
medications|4540,4551
.|4551,4552
<EOL>|4552,4553
<EOL>|4553,4554
-|4554,4555
You|4555,4558
have|4559,4563
also|4564,4568
been|4569,4573
given|4574,4579
Additional|4580,4590
Medications|4591,4602
to|4603,4605
control|4606,4613
<EOL>|4614,4615
your|4615,4619
pain|4620,4624
.|4624,4625
Please|4627,4633
allow|4634,4639
72|4640,4642
hours|4643,4648
for|4649,4652
refill|4653,4659
of|4660,4662
narcotic|4663,4671
<EOL>|4672,4673
prescriptions|4673,4686
,|4686,4687
so|4688,4690
plan|4691,4695
ahead|4696,4701
.|4701,4702
You|4704,4707
can|4708,4711
either|4712,4718
have|4719,4723
them|4724,4728
mailed|4729,4735
<EOL>|4736,4737
to|4737,4739
your|4740,4744
home|4745,4749
or|4750,4752
pick|4753,4757
them|4758,4762
up|4763,4765
at|4766,4768
the|4769,4772
clinic|4773,4779
located|4780,4787
on|4788,4790
_|4791,4792
_|4792,4793
_|4793,4794
.|4794,4795
<EOL>|4796,4797
We|4798,4800
are|4801,4804
not|4805,4808
allowed|4809,4816
to|4817,4819
call|4820,4824
in|4825,4827
narcotic|4828,4836
(|4837,4838
oxycontin|4838,4847
,|4847,4848
oxycodone|4849,4858
,|4858,4859
<EOL>|4860,4861
percocet|4861,4869
)|4869,4870
prescriptions|4871,4884
to|4885,4887
the|4888,4891
pharmacy|4892,4900
.|4900,4901
In|4904,4906
addition|4907,4915
,|4915,4916
we|4917,4919
are|4920,4923
<EOL>|4924,4925
only|4925,4929
allowed|4930,4937
to|4938,4940
write|4941,4946
for|4947,4950
pain|4951,4955
medications|4956,4967
for|4968,4971
90|4972,4974
days|4975,4979
from|4980,4984
the|4985,4988
<EOL>|4989,4990
date|4990,4994
of|4995,4997
surgery|4998,5005
.|5005,5006
<EOL>|5006,5007
<EOL>|5007,5008
-|5008,5009
Follow|5009,5015
up|5016,5018
:|5018,5019
<EOL>|5019,5020
oPlease|5020,5027
Call|5028,5032
the|5033,5036
office|5037,5043
_|5044,5045
_|5045,5046
_|5046,5047
and|5048,5051
make|5052,5056
an|5057,5059
appointment|5060,5071
<EOL>|5072,5073
with|5073,5077
Dr.|5078,5081
_|5082,5083
_|5083,5084
_|5084,5085
2|5086,5087
weeks|5088,5093
after|5094,5099
the|5100,5103
day|5104,5107
of|5108,5110
your|5111,5115
operation|5116,5125
if|5126,5128
<EOL>|5129,5130
this|5130,5134
has|5135,5138
not|5139,5142
been|5143,5147
done|5148,5152
already|5153,5160
.|5160,5161
<EOL>|5161,5162
oAt|5162,5165
the|5166,5169
2|5170,5171
-|5171,5172
week|5172,5176
visit|5177,5182
we|5183,5185
will|5186,5190
check|5191,5196
your|5197,5201
incision|5202,5210
,|5210,5211
take|5212,5216
baseline|5217,5225
<EOL>|5226,5227
x|5227,5228
rays|5229,5233
and|5234,5237
answer|5238,5244
any|5245,5248
questions|5249,5258
.|5258,5259
<EOL>|5259,5260
oWe|5260,5263
will|5264,5268
then|5269,5273
see|5274,5277
you|5278,5281
at|5282,5284
6|5285,5286
weeks|5287,5292
from|5293,5297
the|5298,5301
day|5302,5305
of|5306,5308
the|5309,5312
operation|5313,5322
.|5322,5323
<EOL>|5324,5325
At|5325,5327
that|5328,5332
time|5333,5337
we|5338,5340
will|5341,5345
most|5346,5350
likely|5351,5357
obtain|5358,5364
Flexion|5365,5372
/|5372,5373
Extension|5373,5382
X-rays|5383,5389
<EOL>|5390,5391
and|5391,5394
often|5395,5400
able|5401,5405
to|5406,5408
place|5409,5414
you|5415,5418
in|5419,5421
a|5422,5423
soft|5424,5428
collar|5429,5435
which|5436,5441
you|5442,5445
will|5446,5450
wean|5451,5455
<EOL>|5456,5457
out|5457,5460
of|5461,5463
over|5464,5468
1|5469,5470
week|5471,5475
.|5475,5476
<EOL>|5478,5479
<EOL>|5479,5480
Please|5480,5486
call|5487,5491
the|5492,5495
office|5496,5502
if|5503,5505
you|5506,5509
have|5510,5514
a|5515,5516
fever|5517,5522
>|5522,5523
101.5|5523,5528
degrees|5529,5536
<EOL>|5537,5538
Fahrenheit|5538,5548
,|5548,5549
drainage|5550,5558
from|5559,5563
your|5564,5568
wound|5569,5574
,|5574,5575
or|5576,5578
have|5579,5583
any|5584,5587
questions|5588,5597
.|5597,5598
<EOL>|5598,5599
<EOL>|5599,5600
Physical|5600,5608
Therapy|5609,5616
:|5616,5617
<EOL>|5617,5618
activity|5618,5626
as|5627,5629
tolerated|5630,5639
<EOL>|5639,5640
C|5640,5641
-|5641,5642
collar|5642,5648
full|5649,5653
time|5654,5658
for|5659,5662
12|5663,5665
weeks|5666,5671
<EOL>|5671,5672
may|5672,5675
use|5676,5679
ambulatory|5680,5690
assistive|5691,5700
devices|5701,5708
for|5709,5712
safety|5713,5719
<EOL>|5719,5720
no|5720,5722
bending|5724,5731
twisting|5732,5740
,|5740,5741
or|5742,5744
lifting|5745,5752
>|5753,5754
5lbs|5754,5758
<EOL>|5758,5759
Treatment|5759,5768
Frequency|5769,5778
:|5778,5779
<EOL>|5779,5780
monitor|5780,5787
skin|5788,5792
at|5793,5795
chin|5796,5800
and|5801,5804
back|5805,5809
of|5810,5812
head|5813,5817
for|5818,5821
breakdown|5822,5831
in|5832,5834
C|5835,5836
-|5836,5837
collar|5837,5843
<EOL>|5843,5844
<EOL>|5845,5846
Followup|5846,5854
Instructions|5855,5867
:|5867,5868
<EOL>|5868,5869
_|5869,5870
_|5870,5871
_|5871,5872
<EOL>|5872,5873

