 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|185,194|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|222,231|false|false|false|C1999232|Attending (action)|Attending
Disorder|Disease or Syndrome|Chief Complaint|257,266|false|false|false|C0018965|Hematuria|Hematuria
Finding|Sign or Symptom|Chief Complaint|268,276|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Classification|Chief Complaint|279,284|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|285,293|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|285,293|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|297,315|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|306,315|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|306,315|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|306,315|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|306,315|false|false|false|C0184661|Interventional procedure|Procedure
Drug|Organic Chemical|History of Present Illness|384,391|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|History of Present Illness|384,391|false|false|false|C0728963|Lovenox|lovenox
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|394,401|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|394,401|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|394,401|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|394,408|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|History of Present Illness|402,408|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|423,426|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|History of Present Illness|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|History of Present Illness|427,430|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Disorder|Disease or Syndrome|History of Present Illness|432,435|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|432,435|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|History of Present Illness|432,435|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|History of Present Illness|432,435|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|History of Present Illness|432,435|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|History of Present Illness|432,435|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|History of Present Illness|436,443|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|436,454|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|444,454|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|460,465|false|false|false|C0020885|ileum|ileal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|460,470|false|false|false|C1550266|Ileal Loop|ileal loop
Finding|Finding|History of Present Illness|472,481|false|false|false|C0439843;C3840275|Diversion|diversion
Finding|Functional Concept|History of Present Illness|472,481|false|false|false|C0439843;C3840275|Diversion|diversion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|472,481|false|false|false|C0185033|Diversion procedure|diversion
Disorder|Disease or Syndrome|History of Present Illness|486,494|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|495,506|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Location or Region|History of Present Illness|518,527|false|false|false|C0000726|Abdomen|abdominal
Drug|Substance|History of Present Illness|529,534|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|529,534|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Health Care Activity|History of Present Illness|545,554|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|545,554|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Body Substance|History of Present Illness|558,566|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|History of Present Illness|558,566|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|558,566|false|false|false|C0013103|Drainage procedure|drainage
Anatomy|Body Location or Region|History of Present Illness|586,595|false|false|false|C0000726|Abdomen|abdominal
Procedure|Diagnostic Procedure|History of Present Illness|586,603|false|false|false|C4481095|abdominal imaging|abdominal imaging
Finding|Finding|History of Present Illness|596,603|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|History of Present Illness|596,603|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Idea or Concept|History of Present Illness|610,619|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Finding|Finding|History of Present Illness|637,643|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|637,643|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|History of Present Illness|645,659|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Finding|Intellectual Product|History of Present Illness|712,723|false|false|false|C1547992|Outside Lab|outside lab
Finding|Gene or Genome|History of Present Illness|720,723|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|History of Present Illness|720,723|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|History of Present Illness|724,729|false|false|false|C1554112|MDF Attribute Type - Value|value
Finding|Body Substance|History of Present Illness|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|732,739|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|History of Present Illness|770,781|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|770,781|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|770,796|false|false|false|C0948143|Nephrostomy tube placement|nephrostomy tube placement
Finding|Functional Concept|History of Present Illness|782,786|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|History of Present Illness|782,786|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|782,796|false|false|false|C0883304|placement of tube|tube placement
Procedure|Health Care Activity|History of Present Illness|787,796|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|787,796|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Sign or Symptom|History of Present Illness|831,843|false|false|false|C3714552|Weakness|feeling weak
Finding|Intellectual Product|History of Present Illness|839,843|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|History of Present Illness|839,843|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Daily or Recreational Activity|History of Present Illness|876,885|false|false|false|C0015259|Exercise|exercises
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|876,885|false|false|false|C0452240|Physical therapy exercises|exercises
Finding|Finding|History of Present Illness|891,903|false|false|false|C0030252|Palpitations|palpitations
Finding|Daily or Recreational Activity|History of Present Illness|909,919|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|History of Present Illness|909,919|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Anatomy|Body Location or Region|History of Present Illness|939,944|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|939,944|false|false|false|C0741025|Chest problem|chest
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|983,988|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|History of Present Illness|983,988|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|History of Present Illness|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|History of Present Illness|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|History of Present Illness|983,988|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|History of Present Illness|983,988|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|983,988|false|false|false|C0031765|Phototherapy|light
Finding|Daily or Recreational Activity|History of Present Illness|1002,1012|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Finding|Functional Concept|History of Present Illness|1002,1012|false|false|false|C0080331;C0945826|Ambulation;Walking (function)|ambulation
Disorder|Disease or Syndrome|History of Present Illness|1036,1045|false|false|false|C0018965|Hematuria|hematuria
Finding|Intellectual Product|History of Present Illness|1053,1056|false|false|false|C1552710|Bag Data Type|bag
Finding|Intellectual Product|History of Present Illness|1072,1075|false|false|false|C1552710|Bag Data Type|bag
Anatomy|Anatomical Structure|History of Present Illness|1097,1105|false|false|false|C0559495|Urological stoma|Urostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1097,1105|false|false|false|C0856443|Urostomy procedure|Urostomy
Disorder|Cell or Molecular Dysfunction|History of Present Illness|1127,1135|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|History of Present Illness|1127,1135|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|History of Present Illness|1127,1135|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|History of Present Illness|1127,1139|false|false|false|C1446409|Positive|positive for
Disorder|Disease or Syndrome|History of Present Illness|1140,1149|false|false|false|C0018965|Hematuria|hematuria
Event|Occupational Activity|History of Present Illness|1194,1204|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|1194,1204|false|false|false|C0376636|Disease Management|management
Finding|Idea or Concept|History of Present Illness|1218,1225|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Gene or Genome|History of Present Illness|1242,1246|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1242,1246|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Lab|Laboratory or Test Result|History of Present Illness|1291,1295|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|History of Present Illness|1311,1314|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|History of Present Illness|1328,1337|false|false|false|C0005821|Blood Platelets|platelets
Drug|Pharmacologic Substance|History of Present Illness|1328,1337|false|false|false|C0443116|Platelets Product|platelets
Procedure|Laboratory Procedure|History of Present Illness|1328,1337|false|false|false|C0032181|Platelet count (procedure)|platelets
Drug|Biologically Active Substance|History of Present Illness|1378,1381|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1378,1381|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|History of Present Illness|1378,1381|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Finding|Finding|History of Present Illness|1412,1423|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1412,1423|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Finding|Intellectual Product|History of Present Illness|1424,1429|false|false|false|C1547937||tubes
Anatomy|Cell|History of Present Illness|1441,1444|false|false|false|C0023516|Leukocytes|WBC
Finding|Finding|History of Present Illness|1446,1454|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|History of Present Illness|1446,1454|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Anatomy|Cell|History of Present Illness|1456,1466|false|false|false|C0023516|Leukocytes|leukocytes
Finding|Body Substance|History of Present Illness|1456,1466|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Finding|Intellectual Product|History of Present Illness|1456,1466|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|leukocytes
Finding|Gene or Genome|History of Present Illness|1472,1477|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Disorder|Disease or Syndrome|History of Present Illness|1478,1483|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|History of Present Illness|1478,1483|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|History of Present Illness|1488,1495|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|1488,1495|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Attribute|Clinical Attribute|History of Present Illness|1514,1520|false|false|false|C1644645||CT abd
Anatomy|Body Location or Region|History of Present Illness|1517,1520|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|History of Present Illness|1517,1520|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1521,1527|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|History of Present Illness|1521,1527|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|History of Present Illness|1521,1527|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|History of Present Illness|1521,1527|false|false|false|C0812455|Pelvis problem|pelvis
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|1532,1540|false|false|false|C0009924|Contrast Media|contrast
Finding|Intellectual Product|History of Present Illness|1542,1550|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Procedure|Health Care Activity|History of Present Illness|1551,1560|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1551,1560|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|History of Present Illness|1574,1586|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Finding|Intellectual Product|History of Present Illness|1607,1612|false|false|false|C1547937||tubes
Finding|Conceptual Entity|History of Present Illness|1618,1626|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|History of Present Illness|1618,1626|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Disorder|Disease or Syndrome|History of Present Illness|1627,1648|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Finding|Pathologic Function|History of Present Illness|1656,1664|true|false|false|C0018944|Hematoma|hematoma
Finding|Body Substance|History of Present Illness|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1670,1677|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Activity|History of Present Illness|1700,1707|false|false|false|C1706079||arrival
Finding|Functional Concept|History of Present Illness|1700,1707|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|1715,1720|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1722,1729|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|History of Present Illness|1756,1775|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1756,1775|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1769,1775|false|false|false|C0225386|Breath|breath
Finding|Idea or Concept|History of Present Illness|1798,1809|false|false|false|C2699427|Conjunction|conjunction
Finding|Finding|History of Present Illness|1816,1822|false|false|false|C4554530|Bloody|bloody
Finding|Conceptual Entity|History of Present Illness|1823,1829|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|History of Present Illness|1823,1829|false|false|false|C3251815|Measurement of fluid output|output
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1839,1845|false|false|false|C0029473|Ostomy|ostomy
Finding|Intellectual Product|History of Present Illness|1846,1851|false|false|false|C1547937||tubes
Finding|Conceptual Entity|History of Present Illness|1872,1878|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|History of Present Illness|1872,1878|false|false|false|C3251815|Measurement of fluid output|output
Finding|Finding|History of Present Illness|1889,1900|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1889,1900|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Finding|Intellectual Product|History of Present Illness|1901,1906|false|false|false|C1547937||tubes
Finding|Idea or Concept|History of Present Illness|1942,1950|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Gene or Genome|History of Present Illness|1958,1961|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Anatomy|Body Location or Region|History of Present Illness|1992,1997|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1992,1997|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|2016,2020|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|2016,2020|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2016,2020|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|2024,2032|true|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|2024,2032|true|false|false|C0033095||pressure
Drug|Organic Chemical|History of Present Illness|2045,2050|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|2045,2050|true|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|2045,2050|true|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|2052,2057|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|2052,2057|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|2060,2066|false|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|History of Present Illness|2068,2077|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|2068,2082|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|2078,2082|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|2078,2082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2078,2082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|2087,2095|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2087,2095|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2124,2130|false|false|false|C0029473|Ostomy|ostomy
Finding|Finding|History of Present Illness|2162,2171|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|2162,2171|true|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|2162,2171|true|false|false|C2229507|sensory exam|sensation
Finding|Sign or Symptom|History of Present Illness|2175,2182|false|false|false|C0013428|Dysuria|dysuria
Finding|Body Substance|History of Present Illness|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|2185,2192|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Sign or Symptom|History of Present Illness|2199,2212|false|false|false|C0849959|feeling dizzy|feeling dizzy
Finding|Sign or Symptom|History of Present Illness|2207,2212|false|false|false|C0012833|Dizziness|dizzy
Finding|Sign or Symptom|History of Present Illness|2217,2228|false|false|false|C0220870|Lightheadedness|lightheaded
Finding|Finding|History of Present Illness|2261,2273|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|Past Medical History|2303,2315|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Past Medical History|2325,2328|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2325,2328|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|Past Medical History|2325,2328|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|Past Medical History|2325,2328|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|Past Medical History|2325,2328|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|Past Medical History|2325,2328|false|false|false|C0031150|Laparoscopy|lap
Finding|Functional Concept|Past Medical History|2344,2348|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Past Medical History|2344,2353|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2344,2353|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|Past Medical History|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Past Medical History|2349,2353|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Past Medical History|2349,2353|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|Past Medical History|2349,2365|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2349,2365|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Finding|Functional Concept|Past Medical History|2354,2365|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|2354,2365|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2354,2365|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2375,2386|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|Past Medical History|2399,2402|false|false|false|C1114365||age
Drug|Biologically Active Substance|Past Medical History|2399,2402|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Past Medical History|2399,2402|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2412,2419|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|Past Medical History|2412,2419|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2412,2419|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|Past Medical History|2412,2426|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder Cancer
Disorder|Neoplastic Process|Past Medical History|2420,2426|false|false|false|C0006826|Malignant Neoplasms|Cancer
Finding|Finding|Past Medical History|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Past Medical History|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Past Medical History|2427,2431|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Past Medical History|2427,2437|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|Past Medical History|2427,2437|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|Past Medical History|2432,2437|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Past Medical History|2432,2437|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|Past Medical History|2438,2441|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|Past Medical History|2438,2441|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|Past Medical History|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|Past Medical History|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|Past Medical History|2438,2441|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Finding|Intellectual Product|Past Medical History|2464,2468|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2474,2480|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|Past Medical History|2474,2484|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Finding|Gene or Genome|Past Medical History|2481,2484|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Past Medical History|2481,2484|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Past Medical History|2481,2484|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Neoplastic Process|Past Medical History|2487,2495|false|false|false|C1269955|Tumor Cell Invasion|invasion
Finding|Pathologic Function|Past Medical History|2487,2495|false|false|false|C2699153|Cell Invasion|invasion
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2501,2508|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Past Medical History|2501,2508|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2501,2508|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2501,2513|false|false|false|C0458421|Wall of bladder|bladder wall
Disorder|Disease or Syndrome|Past Medical History|2528,2532|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Past Medical History|2528,2539|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Past Medical History|2528,2539|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Past Medical History|2533,2539|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Past Medical History|2533,2539|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|Past Medical History|2544,2552|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2553,2560|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|2553,2560|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|2553,2560|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|2553,2560|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2553,2565|false|false|false|C0447612|Vaginal wall|vaginal wall
Finding|Functional Concept|Past Medical History|2573,2580|false|false|false|C0332305|With staging|staging
Finding|Finding|Past Medical History|2590,2602|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2590,2602|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2607,2629|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2617,2629|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|Past Medical History|2634,2639|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|Past Medical History|2634,2646|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2640,2646|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|Past Medical History|2640,2646|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|Past Medical History|2640,2646|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|Past Medical History|2640,2646|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Procedure|Diagnostic Procedure|Past Medical History|2640,2646|false|false|false|C0869889|examination of uterus|uterus
Disorder|Neoplastic Process|Past Medical History|2650,2657|false|false|false|C0023267|Fibroid Tumor|fibroid
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2680,2686|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2680,2697|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|Past Medical History|2687,2692|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2687,2697|false|false|false|C0024204|lymph nodes|lymph node
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2698,2707|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Drug|Chemical Viewed Structurally|Past Medical History|2714,2721|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2714,2732|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2722,2732|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|Past Medical History|2737,2745|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2746,2757|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2763,2770|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|2763,2770|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|2763,2770|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|2763,2770|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Machine Activity|Past Medical History|2772,2786|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2772,2786|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2792,2797|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|Past Medical History|2792,2805|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2792,2805|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|Past Medical History|2806,2814|false|false|false|C1706214|Creation|creation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2806,2814|false|false|false|C0441513|Surgical construction|creation
Finding|Finding|Past Medical History|2843,2853|false|false|false|C0004610|Bacteremia|bacteremia
Finding|Functional Concept|Past Medical History|2858,2869|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|Past Medical History|2858,2869|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Functional Concept|Past Medical History|2873,2888|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|Past Medical History|2890,2895|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Past Medical History|2890,2895|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Past Medical History|2896,2906|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Past Medical History|2896,2906|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Past Medical History|2896,2906|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Past Medical History|2896,2906|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|Past Medical History|2915,2920|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Past Medical History|2915,2920|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2915,2930|false|false|false|C3495845|Drain placement|drain placement
Procedure|Health Care Activity|Past Medical History|2921,2930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2921,2930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Anatomy|Body Location or Region|Past Medical History|2955,2958|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Past Medical History|2955,2958|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Past Medical History|2955,2958|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Organic Chemical|Past Medical History|2969,2976|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Past Medical History|2969,2976|false|false|false|C0728963|Lovenox|lovenox
Finding|Classification|Family Medical History|3018,3026|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Family Medical History|3018,3026|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Family Medical History|3018,3026|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|Family Medical History|3018,3030|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3031,3038|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Family Medical History|3031,3038|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3031,3038|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Family Medical History|3031,3041|false|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Procedure|Health Care Activity|General Exam|3087,3096|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|General Exam|3097,3105|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3097,3105|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3097,3105|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3097,3110|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3097,3110|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|General Exam|3106,3110|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3106,3110|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|General Exam|3140,3145|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|VITAL
Attribute|Clinical Attribute|General Exam|3140,3151|false|false|false|C0488614;C0518766|Vital signs|VITAL SIGNS
Procedure|Health Care Activity|General Exam|3140,3151|false|false|false|C0150404|Taking vital signs|VITAL SIGNS
Finding|Finding|General Exam|3146,3151|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|SIGNS
Finding|Functional Concept|General Exam|3146,3151|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|SIGNS
Finding|Gene or Genome|General Exam|3153,3157|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|3153,3157|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Attribute|Clinical Attribute|General Exam|3191,3195|false|false|false|C2317096|Saturation of Peripheral Oxygen|Spo2
Finding|Classification|General Exam|3203,3210|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3203,3210|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|3212,3216|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|3241,3261|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|3247,3252|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|3253,3261|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3253,3261|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|General Exam|3263,3270|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3263,3270|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|General Exam|3280,3287|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|3288,3293|false|false|false|C0024109|Lung|LUNGS
Finding|Idea or Concept|General Exam|3295,3300|false|false|false|C1550016|Remote control command - Clear|clear
Procedure|Diagnostic Procedure|General Exam|3304,3316|false|false|false|C0004339|Auscultation|auscultation
Anatomy|Body Location or Region|General Exam|3330,3337|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3330,3337|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3330,3337|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3339,3343|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Procedure|Diagnostic Procedure|General Exam|3359,3368|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|General Exam|3377,3382|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3377,3389|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3383,3389|false|false|false|C0037709||sounds
Procedure|Therapeutic or Preventive Procedure|General Exam|3392,3398|false|false|false|C0029473|Ostomy|Ostomy
Disorder|Disease or Syndrome|General Exam|3408,3413|false|false|false|C0155339|Brown Tendon Sheath Syndrome|brown
Finding|Finding|General Exam|3408,3419|false|false|false|C5880922|Brown color of stool|brown stool
Finding|Body Substance|General Exam|3414,3419|false|false|false|C0015733|Feces|stool
Finding|Finding|General Exam|3455,3458|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|General Exam|3455,3458|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Finding|General Exam|3459,3465|false|false|false|C4554530|Bloody|bloody
Finding|Finding|General Exam|3459,3471|false|false|false|C0473237|Frank hematuria|bloody urine
Finding|Body Substance|General Exam|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|General Exam|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|General Exam|3466,3471|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Finding|General Exam|3483,3494|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|General Exam|3483,3494|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Finding|Intellectual Product|General Exam|3495,3500|false|false|false|C1547937||tubes
Disorder|Disease or Syndrome|General Exam|3510,3515|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|3510,3515|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|General Exam|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|General Exam|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|General Exam|3517,3522|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Part, Organ, or Organ Component|General Exam|3525,3536|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|General Exam|3541,3546|true|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3541,3546|true|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|3548,3552|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3548,3552|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|3557,3561|false|false|false|C5575035|Well (answer to question)|well
Finding|Body Substance|General Exam|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3599,3608|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3599,3608|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|General Exam|3609,3617|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3609,3617|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3609,3617|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3609,3622|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3609,3622|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|General Exam|3618,3622|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3618,3622|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|3686,3693|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3686,3693|false|false|false|C3812897|General medical service|GENERAL
Finding|Finding|General Exam|3695,3699|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|3724,3744|false|false|false|C2051415|patient appears in no acute distress (physical finding)|in no acute distress
Finding|Intellectual Product|General Exam|3730,3735|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|3736,3744|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3736,3744|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|General Exam|3746,3753|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3746,3753|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|General Exam|3763,3770|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|3771,3776|false|false|false|C0024109|Lung|LUNGS
Finding|Idea or Concept|General Exam|3778,3783|false|false|false|C1550016|Remote control command - Clear|clear
Procedure|Diagnostic Procedure|General Exam|3787,3799|false|false|false|C0004339|Auscultation|auscultation
Anatomy|Body Location or Region|General Exam|3813,3820|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3813,3820|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|General Exam|3813,3820|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3822,3826|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Procedure|Diagnostic Procedure|General Exam|3842,3851|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|General Exam|3860,3865|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3860,3872|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3866,3872|false|false|false|C0037709||sounds
Finding|Finding|General Exam|3909,3912|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|General Exam|3909,3912|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Finding|General Exam|3913,3919|false|false|false|C4554530|Bloody|bloody
Finding|Finding|General Exam|3913,3925|false|false|false|C0473237|Frank hematuria|bloody urine
Finding|Body Substance|General Exam|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|General Exam|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|General Exam|3920,3925|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Finding|General Exam|3938,3949|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|General Exam|3938,3949|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Finding|Intellectual Product|General Exam|3950,3955|false|false|false|C1547937||tubes
Anatomy|Body Part, Organ, or Organ Component|General Exam|3965,3976|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Attribute|Clinical Attribute|General Exam|3981,3986|true|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3981,3986|true|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|3988,3992|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3988,3992|true|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|3997,4001|false|false|false|C5575035|Well (answer to question)|well
Procedure|Health Care Activity|General Exam|4050,4059|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|4060,4064|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4094,4099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4094,4099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4100,4103|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4108,4111|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4108,4111|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4108,4111|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4118,4121|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4118,4121|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4118,4121|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4118,4121|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4127,4130|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4127,4130|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4138,4141|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4138,4141|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4138,4141|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4145,4148|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4145,4148|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4145,4148|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4145,4148|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4145,4148|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4154,4158|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4186,4189|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4206,4211|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4206,4211|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4212,4215|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4220,4223|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4220,4223|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4220,4223|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4230,4233|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4230,4233|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4230,4233|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4230,4233|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4239,4242|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4239,4242|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4250,4253|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4250,4253|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4250,4253|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4250,4253|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4257,4260|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4257,4260|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4257,4260|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4257,4260|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4257,4260|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4266,4270|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4298,4301|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4318,4323|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4318,4323|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4339,4344|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4350,4353|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|4350,4353|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4453,4458|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4453,4458|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4453,4466|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4453,4466|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4453,4466|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4459,4466|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4459,4466|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4459,4466|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4459,4466|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4459,4466|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4513,4517|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4513,4517|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4513,4517|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Finding|General Exam|4549,4556|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4549,4556|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Procedure|Research Activity|General Exam|4557,4564|false|false|false|C0947630|Scientific Study|STUDIES
Attribute|Clinical Attribute|General Exam|4588,4594|false|false|false|C1644645||CT Abd
Anatomy|Body Location or Region|General Exam|4591,4594|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|General Exam|4591,4594|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Anatomy|Body Location or Region|General Exam|4595,4598|false|false|false|C0449203|PEL (body structure)|Pel
Disorder|Disease or Syndrome|General Exam|4595,4598|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|Pel
Disorder|Neoplastic Process|General Exam|4595,4598|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|Pel
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4603,4611|false|true|false|C0009924|Contrast Media|Contrast
Finding|Intellectual Product|Impression|4632,4640|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Procedure|Health Care Activity|Impression|4641,4650|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Impression|4641,4650|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|Impression|4664,4676|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Finding|Intellectual Product|Impression|4697,4702|false|false|false|C1547937||tubes
Finding|Conceptual Entity|Impression|4708,4716|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Finding|Pathologic Function|Impression|4708,4716|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolved
Disorder|Disease or Syndrome|Impression|4717,4738|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Finding|Pathologic Function|Impression|4748,4756|true|false|false|C0018944|Hematoma|hematoma
Finding|Finding|Impression|4787,4794|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Impression|4787,4794|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Functional Concept|Impression|4802,4807|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Impression|4802,4819|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|Impression|4808,4814|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|Impression|4808,4819|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|Impression|4815,4819|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Impression|4815,4819|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Attribute|Clinical Attribute|Impression|4879,4887|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|Impression|4879,4887|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|Impression|4882,4887|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|4882,4887|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|Impression|4895,4898|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|Impression|4911,4918|false|false|false|C1550127|Special Handling Code - Upright|upright
Phenomenon|Human-caused Phenomenon or Process|Impression|4911,4918|false|false|false|C1550585|Entity Handling - upright|upright
Anatomy|Body Location or Region|Impression|4931,4936|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Impression|4931,4936|false|false|false|C0741025|Chest problem|chest
Finding|Functional Concept|Impression|4940,4945|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Impression|4940,4961|false|false|false|C0230329|Right upper extremity|Right upper extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|4946,4961|false|false|false|C1140618|Upper Extremity|upper extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|4952,4961|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|Impression|4963,4969|false|false|false|C1554204|Role Class - access|access
Procedure|Therapeutic or Preventive Procedure|Impression|4970,4974|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Biologically Active Substance|Impression|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Impression|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Drug|Substance|Impression|4976,4980|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|line
Finding|Intellectual Product|Impression|4976,4980|false|false|false|C1546701|line source specimen code|line
Finding|Gene or Genome|Impression|4998,5001|false|false|false|C1705504;C1823282;C1825626;C1825978|ITFG1 gene;KAT5 wt Allele;METTL8 gene;TIPRL gene|tip
Procedure|Therapeutic or Preventive Procedure|Impression|4998,5001|false|false|false|C0673828|TIP regimen|tip
Finding|Finding|Impression|5015,5018|false|false|false|C0231957|Slow vital capacity|SVC
Finding|Intellectual Product|Impression|5031,5034|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Impression|5031,5034|false|false|false|C1623258|Electrocardiography|EKG
Finding|Finding|Impression|5046,5053|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|Impression|5046,5053|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|Impression|5056,5061|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|Impression|5066,5071|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Intellectual Product|Impression|5107,5113|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|Impression|5116,5120|false|false|false|C0443157|Bony|Bony
Finding|Finding|Impression|5136,5142|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|Impression|5161,5173|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|Impression|5161,5173|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|Impression|5161,5173|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Finding|Body Substance|Impression|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|Impression|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|Impression|5201,5206|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|Impression|5212,5216|false|false|false|C1552822|Table Cell Horizontal Align - left|LEFT
Finding|Finding|Impression|5217,5228|false|false|false|C0481713|Has nephrostomy|NEPHROSTOMY
Procedure|Therapeutic or Preventive Procedure|Impression|5217,5228|false|false|false|C0278314|Nephrostomy (procedure)|NEPHROSTOMY
Finding|Functional Concept|Impression|5229,5233|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Finding|Gene or Genome|Impression|5229,5233|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|TUBE
Finding|Idea or Concept|Impression|5266,5271|false|false|false|C1546485|Diagnosis Type - Final|FINAL
Finding|Intellectual Product|Impression|5266,5278|false|false|false|C0460114|Final report|FINAL REPORT
Attribute|Clinical Attribute|Impression|5272,5278|false|false|false|C4255046||REPORT
Finding|Intellectual Product|Impression|5272,5278|false|false|false|C0684224|Report (document)|REPORT
Procedure|Health Care Activity|Impression|5272,5278|false|false|false|C0700287|Reporting|REPORT
Finding|Body Substance|Impression|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|Impression|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|Impression|5286,5291|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Procedure|Laboratory Procedure|Impression|5286,5299|false|false|false|C0430404|Urine culture|URINE CULTURE
Drug|Biomedical or Dental Material|Impression|5292,5299|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|Impression|5292,5299|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|Impression|5292,5299|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|Impression|5292,5299|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|Impression|5301,5306|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|Impression|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|Impression|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|Impression|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|Impression|5318,5324|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|Impression|5318,5324|true|false|false|C2911660|Growth action|GROWTH
Finding|Body Substance|Impression|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Impression|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Impression|5345,5354|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Impression|5345,5354|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|Impression|5355,5359|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Impression|5389,5394|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5389,5394|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|5395,5398|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|5403,5406|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|5403,5406|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|5403,5406|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|5413,5416|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|5413,5416|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|5413,5416|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|5413,5416|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|5422,5425|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|5422,5425|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|5433,5436|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Impression|5433,5436|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|5433,5436|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|5433,5436|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|5440,5443|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|5440,5443|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Impression|5440,5443|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|5440,5443|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|5440,5443|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Impression|5449,5453|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|5481,5484|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|5501,5506|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5501,5506|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|5501,5514|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|5501,5514|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|5501,5514|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|5507,5514|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|5507,5514|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|5507,5514|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Impression|5507,5514|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|5507,5514|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|5559,5563|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|5559,5563|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|5559,5563|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|5588,5593|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5588,5593|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|5588,5601|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|5594,5601|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Impression|5594,5601|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|5594,5601|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Idea or Concept|Hospital Course|5666,5670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|5666,5670|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Conceptual Entity|Hospital Course|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5686,5693|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5686,5696|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|Hospital Course|5707,5710|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|5707,5710|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|5707,5710|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Organic Chemical|Hospital Course|5718,5725|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|5718,5725|false|false|false|C0728963|Lovenox|lovenox
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5728,5735|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|5728,5735|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5728,5735|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Hospital Course|5728,5742|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|Hospital Course|5736,5742|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5755,5758|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|Hospital Course|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|Hospital Course|5759,5762|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Disorder|Disease or Syndrome|Hospital Course|5764,5767|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5764,5767|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|Hospital Course|5764,5767|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|Hospital Course|5764,5767|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|Hospital Course|5764,5767|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|Hospital Course|5764,5767|false|false|false|C0031150|Laparoscopy|lap
Drug|Chemical Viewed Structurally|Hospital Course|5769,5776|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5769,5787|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5777,5787|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5793,5798|false|false|false|C0020885|ileum|ileal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5793,5803|false|false|false|C1550266|Ileal Loop|ileal loop
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5799,5813|false|false|false|C4489477|Loop diversion|loop diversion
Finding|Finding|Hospital Course|5804,5813|false|false|false|C0439843;C3840275|Diversion|diversion
Finding|Functional Concept|Hospital Course|5804,5813|false|false|false|C0439843;C3840275|Diversion|diversion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5804,5813|false|false|false|C0185033|Diversion procedure|diversion
Disorder|Disease or Syndrome|Hospital Course|5818,5826|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5828,5839|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Location or Region|Hospital Course|5851,5860|false|false|false|C0000726|Abdomen|abdominal
Finding|Body Substance|Hospital Course|5851,5866|false|false|false|C2699330|Abdominal Fluid|abdominal fluid
Drug|Substance|Hospital Course|5861,5866|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|5861,5866|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Health Care Activity|Hospital Course|5878,5887|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5878,5887|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Body Substance|Hospital Course|5891,5899|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Hospital Course|5891,5899|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5891,5899|false|false|false|C0013103|Drainage procedure|drainage
Disorder|Disease or Syndrome|Hospital Course|5922,5936|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Procedure|Health Care Activity|Hospital Course|5948,5957|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5948,5957|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Drug|Organic Chemical|Hospital Course|5971,5974|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|Hospital Course|5971,5974|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|Hospital Course|5971,5974|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Finding|Intellectual Product|Hospital Course|5975,5980|false|false|false|C1547937||tubes
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6006,6011|false|false|false|C0034991|Rehabilitation therapy|rehab
Disorder|Disease or Syndrome|Hospital Course|6017,6026|false|false|false|C0018965|Hematuria|hematuria
Finding|Sign or Symptom|Hospital Course|6031,6039|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Activity|Hospital Course|6045,6052|false|false|false|C1706079||arrival
Finding|Functional Concept|Hospital Course|6045,6052|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Finding|Idea or Concept|Hospital Course|6061,6069|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|6061,6072|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Hospital Course|6073,6078|false|false|false|C0398650|Immune thrombocytopenic purpura|frank
Finding|Finding|Hospital Course|6073,6088|false|false|false|C0473237|Frank hematuria|frank hematuria
Disorder|Disease or Syndrome|Hospital Course|6079,6088|false|false|false|C0018965|Hematuria|hematuria
Anatomy|Anatomical Structure|Hospital Course|6096,6104|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6096,6104|false|false|false|C0856443|Urostomy procedure|urostomy
Finding|Intellectual Product|Hospital Course|6106,6109|false|false|false|C1552710|Bag Data Type|bag
Drug|Organic Chemical|Hospital Course|6114,6117|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|Hospital Course|6114,6117|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|Hospital Course|6114,6117|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Finding|Intellectual Product|Hospital Course|6118,6123|false|false|false|C1547937||tubes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|6129,6139|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Finding|Finding|Hospital Course|6129,6139|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|6129,6139|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Drug|Organic Chemical|Hospital Course|6198,6205|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|6198,6205|false|false|false|C0728963|Lovenox|lovenox
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|6274,6284|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Finding|Finding|Hospital Course|6274,6284|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|6274,6284|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Disorder|Disease or Syndrome|Hospital Course|6299,6308|false|false|false|C0018965|Hematuria|Hematuria
Finding|Finding|Hospital Course|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6313,6319|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Mental Process|Hospital Course|6361,6368|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|6372,6387|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|6372,6387|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6372,6387|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Disorder|Disease or Syndrome|Hospital Course|6393,6402|false|false|false|C0018965|Hematuria|hematuria
Finding|Sign or Symptom|Hospital Course|6425,6434|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Finding|Sign or Symptom|Hospital Course|6435,6443|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Drug|Organic Chemical|Hospital Course|6493,6496|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|Hospital Course|6493,6496|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|Hospital Course|6493,6496|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Finding|Intellectual Product|Hospital Course|6497,6502|false|false|false|C1547937||tubes
Finding|Social Behavior|Hospital Course|6510,6520|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6510,6520|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Body Substance|Hospital Course|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6530,6537|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|6582,6589|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|6582,6589|false|false|false|C0728963|Lovenox|lovenox
Finding|Conceptual Entity|Hospital Course|6590,6599|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6590,6599|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6590,6599|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6590,6599|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Anatomy|Body Location or Region|Hospital Course|6616,6619|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|6616,6619|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|6616,6619|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Mental Process|Hospital Course|6644,6651|false|false|false|C0542559|contextual factors|setting
Event|Activity|Hospital Course|6659,6667|false|false|false|C0237820||recovery
Finding|Organism Function|Hospital Course|6659,6667|false|false|false|C2004454|Recovery - healing process|recovery
Finding|Finding|Hospital Course|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|6674,6681|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6674,6681|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Conceptual Entity|Hospital Course|6729,6738|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6729,6738|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6729,6738|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6729,6738|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Neoplastic Process|Hospital Course|6741,6750|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|6741,6750|false|false|false|C1522484|metastatic qualifier|Secondary
Finding|Finding|Hospital Course|6762,6774|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|Asymptomatic
Finding|Body Substance|Hospital Course|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6787,6794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|Hospital Course|6800,6812|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Mental Process|Hospital Course|6828,6835|false|false|false|C0542559|contextual factors|setting
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6857,6869|false|false|false|C0185111;C0947647|Manipulation procedure;Surgical Manipulation|manipulation
Finding|Finding|Hospital Course|6879,6887|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|Hospital Course|6901,6913|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|6901,6913|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Conceptual Entity|Hospital Course|6918,6927|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|6918,6927|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|6918,6927|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6918,6927|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Antibiotic|Hospital Course|6933,6944|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Disorder|Disease or Syndrome|Hospital Course|6963,6977|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|Hospital Course|6963,6977|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Organic Chemical|Hospital Course|6989,7001|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6989,7001|false|false|false|C0286651|atorvastatin|atorvastatin
Disorder|Disease or Syndrome|Hospital Course|7017,7031|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|7042,7055|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Finding|Idea or Concept|Hospital Course|7091,7103|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Drug|Pharmacologic Substance|Hospital Course|7131,7141|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|7131,7141|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Functional Concept|Hospital Course|7142,7149|false|false|false|C0392747|Changing|Changes
Drug|Organic Chemical|Hospital Course|7151,7158|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Hospital Course|7151,7158|false|false|false|C0728963|Lovenox|Lovenox
Attribute|Clinical Attribute|Hospital Course|7172,7182|false|false|false|C1644645||CT Abdomen
Procedure|Diagnostic Procedure|Hospital Course|7172,7182|false|false|false|C0412620|CT of abdomen|CT Abdomen
Anatomy|Body Location or Region|Hospital Course|7175,7182|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|Hospital Course|7175,7182|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|Hospital Course|7175,7182|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7183,7189|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Anatomy|Body Space or Junction|Hospital Course|7183,7189|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|Pelvis
Disorder|Neoplastic Process|Hospital Course|7183,7189|false|false|false|C0153663|Malignant neoplasm of pelvis|Pelvis
Finding|Finding|Hospital Course|7183,7189|false|false|false|C0812455|Pelvis problem|Pelvis
Finding|Finding|Hospital Course|7222,7229|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Pathologic Function|Hospital Course|7222,7229|false|false|false|C0029053;C1265876|Abnormally opaque structure (morphologic abnormality);Decreased translucency|opacity
Finding|Functional Concept|Hospital Course|7238,7243|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7238,7255|false|false|false|C4281590|Structure of middle lobe of right lung|right middle lobe
Finding|Intellectual Product|Hospital Course|7244,7250|false|false|false|C1552826|Table Cell Vertical Align - middle|middle
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7244,7255|false|false|false|C4281590|Structure of middle lobe of right lung|middle lobe
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7251,7255|false|false|false|C0796494|lobe|lobe
Finding|Gene or Genome|Hospital Course|7251,7255|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|lobe
Attribute|Clinical Attribute|Hospital Course|7314,7322|false|false|false|C0881858||CT chest
Procedure|Diagnostic Procedure|Hospital Course|7314,7322|false|false|false|C0202823|Chest CT|CT chest
Anatomy|Body Location or Region|Hospital Course|7317,7322|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|7317,7322|false|false|false|C0741025|Chest problem|chest
Drug|Organic Chemical|Hospital Course|7334,7337|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Drug|Pharmacologic Substance|Hospital Course|7334,7337|false|false|false|C0033017|Pregnenolone Carbonitrile|PCN
Finding|Gene or Genome|Hospital Course|7334,7337|false|false|false|C1418643;C1826553;C4050150|PCNT gene;PLEC gene;PLEC wt Allele|PCN
Finding|Intellectual Product|Hospital Course|7338,7343|false|false|false|C1547937||tubes
Finding|Idea or Concept|Hospital Course|7364,7378|false|false|false|C0034866|Recommendation|recommendation
Procedure|Health Care Activity|Hospital Course|7391,7406|false|false|false|C0019993|Hospitalization|hospitalization
Procedure|Health Care Activity|Hospital Course|7442,7450|false|false|false|C1522577|follow-up|followup
Finding|Idea or Concept|Hospital Course|7470,7474|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|Hospital Course|7470,7474|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Event|Occupational Activity|Hospital Course|7475,7485|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|7475,7485|false|false|false|C0376636|Disease Management|management
Disorder|Disease or Syndrome|Hospital Course|7505,7514|false|false|false|C0018965|Hematuria|hematuria
Finding|Sign or Symptom|Hospital Course|7522,7537|false|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Functional Concept|Hospital Course|7548,7556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|7548,7556|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|Hospital Course|7560,7566|false|false|false|C0002871|Anemia|anemia
Anatomy|Cell Component|Hospital Course|7570,7573|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|7570,7573|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Pathologic Function|Hospital Course|7609,7617|false|false|false|C0019080|Hemorrhage|bleeding
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Biologically Active Substance|Hospital Course|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Organic Chemical|Hospital Course|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Drug|Pharmacologic Substance|Hospital Course|7622,7632|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|Hemoglobin
Finding|Finding|Hospital Course|7622,7632|false|false|false|C1561562|Hemoglobin finding|Hemoglobin
Procedure|Laboratory Procedure|Hospital Course|7622,7632|false|false|false|C0518015|Hemoglobin measurement|Hemoglobin
Attribute|Clinical Attribute|Hospital Course|7633,7643|false|false|false|C1542366|hematocrit attribute|Hematocrit
Finding|Finding|Hospital Course|7633,7643|false|false|false|C0518014|Hematocrit level|Hematocrit
Procedure|Laboratory Procedure|Hospital Course|7633,7643|false|false|false|C0018935|Hematocrit Measurement|Hematocrit
Finding|Body Substance|Hospital Course|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7647,7656|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7647,7656|false|false|false|C0030685|Patient Discharge|discharge
Event|Occupational Activity|Hospital Course|7670,7674|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|7670,7674|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Event|Activity|Hospital Course|7692,7699|false|false|false|C3812666|Personal Contact|CONTACT
Finding|Functional Concept|Hospital Course|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|7692,7699|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|7692,7699|false|false|false|C0392367|Physical contact|CONTACT
Anatomy|Cell|Hospital Course|7715,7719|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|Hospital Course|7715,7719|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Finding|Idea or Concept|Hospital Course|7727,7731|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7727,7731|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7727,7731|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|7737,7748|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|7737,7748|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|7737,7748|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|7737,7761|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|7752,7761|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|7780,7790|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|7780,7790|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|7780,7795|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|7791,7795|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|7812,7820|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|7812,7820|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|7812,7820|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|7825,7837|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7825,7837|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|7855,7865|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|7855,7865|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|Hospital Course|7855,7872|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|7855,7872|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7866,7872|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|7866,7872|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7866,7872|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Idea or Concept|Hospital Course|7912,7916|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|Hospital Course|7917,7924|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|7917,7924|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|7917,7924|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|7925,7939|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7925,7939|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|7940,7944|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|7949,7962|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|7949,7969|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|7963,7969|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|7963,7969|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|7963,7969|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|7991,8004|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|8007,8010|false|false|false|C0039225|Tablet Dosage Form|TAB
Anatomy|Body System|Hospital Course|8034,8043|false|false|false|C0012240|Gastrointestinal system|Digestive
Finding|Organism Function|Hospital Course|8034,8043|false|false|false|C0012238|Digestion|Digestive
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Enzyme|Hospital Course|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Pharmacologic Substance|Hospital Course|8034,8051|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Procedure|Laboratory Procedure|Hospital Course|8034,8051|false|false|false|C0863186|Digestive enzyme test|Digestive Enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Enzyme|Hospital Course|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Pharmacologic Substance|Hospital Course|8044,8051|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Finding|Functional Concept|Hospital Course|8044,8051|false|false|false|C0014445|enzymology|Enzymes
Disorder|Neoplastic Process|Hospital Course|8068,8071|false|false|false|C1321878|Desmoplastic infantile ganglioglioma|dig
Anatomy|Body Space or Junction|Hospital Course|8087,8091|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8087,8091|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8087,8091|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8087,8091|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Body Substance|Hospital Course|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8102,8111|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8102,8111|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8102,8123|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8112,8123|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8112,8123|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8112,8123|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8129,8141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8129,8141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|8161,8174|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|8161,8181|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8175,8181|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|8175,8181|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8175,8181|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|8205,8218|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|8221,8224|false|false|false|C0039225|Tablet Dosage Form|TAB
Anatomy|Body System|Hospital Course|8250,8259|false|false|false|C0012240|Gastrointestinal system|Digestive
Finding|Organism Function|Hospital Course|8250,8259|false|false|false|C0012238|Digestion|Digestive
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Enzyme|Hospital Course|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Drug|Pharmacologic Substance|Hospital Course|8250,8267|false|false|false|C0544420|Digestive Enzymes|Digestive Enzymes
Procedure|Laboratory Procedure|Hospital Course|8250,8267|false|false|false|C0863186|Digestive enzyme test|Digestive Enzymes
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Enzyme|Hospital Course|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Drug|Pharmacologic Substance|Hospital Course|8260,8267|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|Enzymes
Finding|Functional Concept|Hospital Course|8260,8267|false|false|false|C0014445|enzymology|Enzymes
Disorder|Neoplastic Process|Hospital Course|8284,8287|false|false|false|C1321878|Desmoplastic infantile ganglioglioma|dig
Anatomy|Body Space or Junction|Hospital Course|8303,8307|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|8303,8307|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|8303,8307|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|8303,8307|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Body Substance|Hospital Course|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8319,8328|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8319,8328|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|8319,8340|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|8319,8340|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|8329,8340|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|8329,8340|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|8342,8350|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8342,8350|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|8342,8355|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|8351,8355|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|8351,8355|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|8351,8355|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|8358,8366|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8374,8383|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8374,8383|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8374,8393|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|8384,8393|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|8384,8393|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|8384,8393|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8384,8393|false|false|false|C0011900|Diagnosis|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|8403,8412|false|false|false|C0011900|Diagnosis|Diagnoses
Disorder|Disease or Syndrome|Hospital Course|8414,8423|false|false|false|C0018965|Hematuria|Hematuria
Disorder|Disease or Syndrome|Hospital Course|8425,8431|false|false|false|C0002871|Anemia|anemia
Disorder|Neoplastic Process|Hospital Course|8433,8442|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|8433,8442|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|Hospital Course|8443,8452|false|false|false|C0011900|Diagnosis|Diagnoses
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8454,8461|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|Hospital Course|8454,8461|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8454,8461|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|Hospital Course|8454,8468|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder cancer
Disorder|Neoplastic Process|Hospital Course|8462,8468|false|false|false|C0006826|Malignant Neoplasms|cancer
Disorder|Disease or Syndrome|Hospital Course|8470,8484|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Disorder|Disease or Syndrome|Hospital Course|8487,8501|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Anatomy|Body Location or Region|Hospital Course|8503,8506|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|8503,8506|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|8503,8506|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Mental Process|Discharge Condition|8534,8540|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8534,8547|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8534,8547|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8541,8547|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8541,8547|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|8549,8554|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|8559,8567|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|8569,8591|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8569,8591|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|8578,8591|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8578,8591|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8593,8598|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8593,8598|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8593,8598|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8593,8598|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8603,8614|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8616,8624|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8616,8624|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8616,8624|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8625,8631|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8625,8631|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8633,8643|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8633,8643|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|8646,8657|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8646,8657|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|8686,8690|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|Discharge Instructions|8711,8719|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|8711,8719|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|8727,8731|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|8727,8731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|8727,8731|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|8727,8734|false|false|false|C1555558|care of - AddressPartType|care of
Finding|Idea or Concept|Discharge Instructions|8773,8781|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Disorder|Disease or Syndrome|Discharge Instructions|8795,8800|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|8795,8800|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Discharge Instructions|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Discharge Instructions|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Discharge Instructions|8809,8814|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Mental Process|Discharge Instructions|8829,8836|false|false|false|C1527305|Feelings|feeling
Finding|Intellectual Product|Discharge Instructions|8838,8842|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|8838,8842|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|8843,8854|false|false|false|C0220870|Lightheadedness|lightheaded
Event|Activity|Discharge Instructions|8862,8870|false|false|false|C1709305|Occur (action)|HAPPENED
Disorder|Disease or Syndrome|Discharge Instructions|8917,8922|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|8917,8922|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Pharmacologic Substance|Discharge Instructions|8931,8941|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|8931,8941|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|8943,8950|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Discharge Instructions|8943,8950|false|false|false|C0728963|Lovenox|Lovenox
Disorder|Disease or Syndrome|Discharge Instructions|8980,8985|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|8980,8985|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Disorder|Disease or Syndrome|Discharge Instructions|8991,8996|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|8991,8996|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Body Substance|Discharge Instructions|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Discharge Instructions|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Discharge Instructions|9005,9010|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Idea or Concept|Discharge Instructions|9064,9072|false|false|false|C1547192|Organization unit type - Hospital|HOSPITAL
Drug|Organic Chemical|Discharge Instructions|9159,9166|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Discharge Instructions|9159,9166|false|false|false|C0728963|Lovenox|Lovenox
Attribute|Clinical Attribute|Discharge Instructions|9242,9253|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9242,9253|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|9242,9253|false|false|false|C4284232|Medications|medications
Procedure|Health Care Activity|Discharge Instructions|9275,9283|false|false|false|C1522577|follow-up|followup
Event|Activity|Discharge Instructions|9284,9296|false|false|false|C0003629|Appointments|appointments
Finding|Intellectual Product|Discharge Instructions|9332,9340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9332,9340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|9348,9352|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|9348,9352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9348,9352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9348,9355|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|Discharge Instructions|9391,9399|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9400,9412|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|9400,9412|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

