 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
.|12,13
Unit|23,27
No|28,30
:|30,31
_|34,35
_|35,36
_|36,37
<EOL>|37,38
<EOL>|39,40
Admission|40,49
Date|50,54
:|54,55
_|57,58
_|58,59
_|59,60
Discharge|74,83
Date|84,88
:|88,89
_|92,93
_|93,94
_|94,95
<EOL>|95,96
<EOL>|97,98
Date|98,102
of|103,105
Birth|106,111
:|111,112
_|114,115
_|115,116
_|116,117
Sex|130,133
:|133,134
F|137,138
<EOL>|138,139
<EOL>|140,141
Service|141,148
:|148,149
MEDICINE|150,158
<EOL>|158,159
<EOL>|160,161
Tramadol|173,181
<EOL>|181,182
<EOL>|183,184
Attending|184,193
:|193,194
_|195,196
_|196,197
_|197,198
.|198,199
<EOL>|199,200
<EOL>|201,202
Abdominal|219,228
distention|229,239
,|239,240
back|241,245
pain|246,250
,|250,251
fever|252,257
;|257,258
leukocytosis|259,271
.|271,272
<EOL>|272,273
<EOL>|274,275
Major|275,280
Surgical|281,289
or|290,292
Invasive|293,301
Procedure|302,311
:|311,312
<EOL>|312,313
Paracentesis|313,325
x|326,327
3|328,329
.|329,330
<EOL>|330,331
<EOL>|331,332
<EOL>|333,334
This|362,366
is|367,369
a|370,371
_|372,373
_|373,374
_|374,375
woman|376,381
with|382,386
a|387,388
history|389,396
of|397,399
ETOH|400,404
abuse|405,410
who|411,414
<EOL>|415,416
presents|416,424
with|425,429
abdominal|430,439
distention|440,450
,|450,451
back|452,456
pain|457,461
,|461,462
fever|463,468
,|468,469
and|470,473
<EOL>|474,475
elevated|475,483
white|484,489
count|490,495
from|496,500
Liver|501,506
Clinic|507,513
.|513,514
Ms.|516,519
_|520,521
_|521,522
_|522,523
was|524,527
<EOL>|528,529
recently|529,537
admitted|538,546
to|547,549
this|550,554
hospital|555,563
about|564,569
1|570,571
week|572,576
ago|577,580
for|581,584
<EOL>|585,586
treatment|586,595
of|596,598
ascites|599,606
and|607,610
work|611,615
-|615,616
up|616,618
of|619,621
alcoholic|622,631
hepatitis|632,641
.|641,642
At|644,646
<EOL>|647,648
that|648,652
time|653,657
she|658,661
had|662,665
a|666,667
diagnostic|668,678
and|679,682
therapeutic|683,694
paracentesis|695,707
and|708,711
<EOL>|712,713
was|713,716
treated|717,724
for|725,728
a|729,730
UTI|731,734
.|734,735
She|737,740
was|741,744
discharged|745,755
home|756,760
and|761,764
instructed|765,775
<EOL>|776,777
to|777,779
follow|780,786
-|786,787
up|787,789
in|790,792
Liver|793,798
Clinic|799,805
in|806,808
1|809,810
week|811,815
.|815,816
On|818,820
day|821,824
of|825,827
presentation|828,840
<EOL>|841,842
to|842,844
liver|845,850
clinic|851,857
,|857,858
patient|859,866
complained|867,877
of|878,880
worsening|881,890
abdominal|891,900
pain|901,905
<EOL>|906,907
and|907,910
low|911,914
-|914,915
grade|915,920
fevers|921,927
at|928,930
home|931,935
.|935,936
Her|938,941
labwork|942,949
was|950,953
also|954,958
significant|959,970
<EOL>|971,972
for|972,975
an|976,978
elevated|979,987
white|988,993
count|994,999
.|999,1000
As|1002,1004
such|1005,1009
,|1009,1010
Ms.|1011,1014
_|1015,1016
_|1016,1017
_|1017,1018
was|1019,1022
<EOL>|1023,1024
admitted|1024,1032
for|1033,1036
work|1037,1041
-|1041,1042
up|1042,1044
of|1045,1047
fever|1048,1053
and|1054,1057
white|1058,1063
count|1064,1069
,|1069,1070
and|1071,1074
for|1075,1078
treatment|1079,1088
<EOL>|1089,1090
of|1090,1092
recurrent|1093,1102
ascites|1103,1110
.|1110,1111
<EOL>|1111,1112
<EOL>|1113,1114
-|1136,1137
-|1137,1138
Alcohol|1138,1145
abuse|1146,1151
<EOL>|1151,1152
-|1152,1153
-|1153,1154
Chronic|1154,1161
back|1162,1166
pain|1167,1171
<EOL>|1171,1172
<EOL>|1173,1174
:|1188,1189
<EOL>|1189,1190
_|1190,1191
_|1191,1192
_|1192,1193
<EOL>|1193,1194
:|1208,1209
<EOL>|1209,1210
Breast|1210,1216
cancer|1217,1223
in|1224,1226
mother|1227,1233
age|1234,1237
_|1238,1239
_|1239,1240
_|1240,1241
,|1241,1242
No|1243,1245
IBD|1246,1249
,|1249,1250
liver|1251,1256
failure|1257,1264
.|1264,1265
Multiple|1267,1275
<EOL>|1276,1277
relatives|1277,1286
with|1287,1291
alcoholism|1292,1302
.|1302,1303
<EOL>|1303,1304
<EOL>|1305,1306
VS|1321,1323
:|1323,1324
97.9|1325,1329
,|1329,1330
103|1331,1334
/|1334,1335
73|1335,1337
,|1337,1338
86|1339,1341
,|1341,1342
18|1343,1345
,|1345,1346
96|1347,1349
%|1349,1350
RA|1351,1353
<EOL>|1355,1356
GEN|1356,1359
:|1359,1360
A|1361,1362
/|1362,1363
Ox3|1363,1366
,|1366,1367
pleasant|1368,1376
,|1376,1377
appropriate|1378,1389
,|1389,1390
well|1391,1395
appearing|1396,1405
<EOL>|1407,1408
HEENT|1408,1413
:|1413,1414
No|1415,1417
temporal|1418,1426
wasting|1427,1434
,|1434,1435
JVD|1436,1439
not|1440,1443
elevated|1444,1452
,|1452,1453
neck|1454,1458
veins|1459,1464
fill|1465,1469
<EOL>|1470,1471
from|1471,1475
above|1476,1481
.|1481,1482
<EOL>|1484,1485
CV|1485,1487
:|1487,1488
RRR|1489,1492
,|1492,1493
No|1494,1496
MRG|1497,1500
<EOL>|1502,1503
PULM|1503,1507
:|1507,1508
CTAB|1509,1513
but|1514,1517
decreased|1518,1527
BS|1528,1530
in|1531,1533
R|1534,1535
base|1536,1540
.|1540,1541
<EOL>|1543,1544
ABD|1544,1547
:|1547,1548
Distended|1549,1558
and|1559,1562
tight|1563,1568
,|1568,1569
diffusely|1570,1579
tender|1580,1586
to|1587,1589
palpation|1590,1599
,|1599,1600
BS|1601,1603
+|1603,1604
,|1604,1605
+|1606,1607
<EOL>|1608,1609
passing|1609,1616
flatulence|1617,1627
.|1627,1628
<EOL>|1630,1631
LIMBS|1631,1636
:|1636,1637
2|1638,1639
+|1639,1640
edema|1641,1646
of|1647,1649
the|1650,1653
LEs|1654,1657
to|1658,1660
knee|1661,1665
bilaterally|1666,1677
_|1678,1679
_|1679,1680
_|1680,1681
pulses|1682,1688
2|1689,1690
+|1690,1691
<EOL>|1692,1693
bilaterally|1693,1704
<EOL>|1706,1707
NEURO|1707,1712
:|1712,1713
No|1714,1716
asterixis|1717,1726
,|1726,1727
very|1728,1732
mild|1733,1737
general|1738,1745
tremor|1746,1752
.|1752,1753
<EOL>|1753,1754
<EOL>|1755,1756
Pertinent|1756,1765
Results|1766,1773
:|1773,1774
<EOL>|1774,1775
Labs|1775,1779
at|1780,1782
Admission|1783,1792
:|1792,1793
<EOL>|1793,1794
<EOL>|1794,1795
_|1795,1796
_|1796,1797
_|1797,1798
09|1799,1801
:|1801,1802
47AM|1802,1806
BLOOD|1807,1812
WBC|1813,1816
-|1816,1817
26|1817,1819
.|1819,1820
2|1820,1821
*|1821,1822
#|1822,1823
RBC|1824,1827
-|1827,1828
3|1828,1829
.|1829,1830
86|1830,1832
*|1832,1833
Hgb|1834,1837
-|1837,1838
13.0|1838,1842
Hct|1843,1846
-|1846,1847
43.3|1847,1851
<EOL>|1852,1853
MCV|1853,1856
-|1856,1857
112|1857,1860
*|1860,1861
MCH|1862,1865
-|1865,1866
33|1866,1868
.|1868,1869
7|1869,1870
*|1870,1871
MCHC|1872,1876
-|1876,1877
30|1877,1879
.|1879,1880
0|1880,1881
*|1881,1882
RDW|1883,1886
-|1886,1887
12.7|1887,1891
Plt|1892,1895
_|1896,1897
_|1897,1898
_|1898,1899
<EOL>|1899,1900
_|1900,1901
_|1901,1902
_|1902,1903
09|1904,1906
:|1906,1907
47AM|1907,1911
BLOOD|1912,1917
Neuts|1918,1923
-|1923,1924
88|1924,1926
*|1926,1927
Bands|1928,1933
-|1933,1934
1|1934,1935
Lymphs|1936,1942
-|1942,1943
2|1943,1944
*|1944,1945
Monos|1946,1951
-|1951,1952
7|1952,1953
Eos|1954,1957
-|1957,1958
1|1958,1959
<EOL>|1960,1961
Baso|1961,1965
-|1965,1966
1|1966,1967
_|1968,1969
_|1969,1970
_|1970,1971
Myelos|1972,1978
-|1978,1979
0|1979,1980
<EOL>|1980,1981
_|1981,1982
_|1982,1983
_|1983,1984
09|1985,1987
:|1987,1988
20PM|1988,1992
BLOOD|1993,1998
_|1999,2000
_|2000,2001
_|2001,2002
<EOL>|2002,2003
_|2003,2004
_|2004,2005
_|2005,2006
09|2007,2009
:|2009,2010
47AM|2010,2014
BLOOD|2015,2020
UreaN|2021,2026
-|2026,2027
8|2027,2028
Creat|2029,2034
-|2034,2035
0.5|2035,2038
Na|2039,2041
-|2041,2042
133|2042,2045
K|2046,2047
-|2047,2048
5.1|2048,2051
Cl|2052,2054
-|2054,2055
92|2055,2057
*|2057,2058
<EOL>|2059,2060
HCO3|2060,2064
-|2064,2065
26|2065,2067
AnGap|2068,2073
-|2073,2074
20|2074,2076
<EOL>|2076,2077
_|2077,2078
_|2078,2079
_|2079,2080
09|2081,2083
:|2083,2084
47AM|2084,2088
BLOOD|2089,2094
ALT|2095,2098
-|2098,2099
45|2099,2101
*|2101,2102
AST|2103,2106
-|2106,2107
165|2107,2110
*|2110,2111
LD|2112,2114
(|2114,2115
LDH|2115,2118
)|2118,2119
-|2119,2120
345|2120,2123
*|2123,2124
<EOL>|2125,2126
AlkPhos|2126,2133
-|2133,2134
200|2134,2137
*|2137,2138
TotBili|2139,2146
-|2146,2147
2|2147,2148
.|2148,2149
0|2149,2150
*|2150,2151
<EOL>|2151,2152
_|2152,2153
_|2153,2154
_|2154,2155
09|2156,2158
:|2158,2159
47AM|2159,2163
BLOOD|2164,2169
Albumin|2170,2177
-|2177,2178
2|2178,2179
.|2179,2180
9|2180,2181
*|2181,2182
Calcium|2183,2190
-|2190,2191
8|2191,2192
.|2192,2193
1|2193,2194
*|2194,2195
Phos|2196,2200
-|2200,2201
4.0|2201,2204
Mg|2205,2207
-|2207,2208
2.2|2208,2211
<EOL>|2211,2212
_|2212,2213
_|2213,2214
_|2214,2215
09|2216,2218
:|2218,2219
20PM|2219,2223
BLOOD|2224,2229
Ethanol|2230,2237
-|2237,2238
NEG|2238,2241
Bnzodzp|2242,2249
-|2249,2250
NEG|2250,2253
<EOL>|2253,2254
<EOL>|2254,2255
Labs|2255,2259
at|2260,2262
Discharge|2263,2272
:|2272,2273
<EOL>|2273,2274
<EOL>|2274,2275
_|2275,2276
_|2276,2277
_|2277,2278
07|2279,2281
:|2281,2282
20AM|2282,2286
BLOOD|2287,2292
WBC|2293,2296
-|2296,2297
20|2297,2299
.|2299,2300
7|2300,2301
*|2301,2302
RBC|2303,2306
-|2306,2307
3|2307,2308
.|2308,2309
03|2309,2311
*|2311,2312
Hgb|2313,2316
-|2316,2317
10|2317,2319
.|2319,2320
3|2320,2321
*|2321,2322
Hct|2323,2326
-|2326,2327
32|2327,2329
.|2329,2330
0|2330,2331
*|2331,2332
<EOL>|2333,2334
MCV|2334,2337
-|2337,2338
106|2338,2341
*|2341,2342
MCH|2343,2346
-|2346,2347
33|2347,2349
.|2349,2350
9|2350,2351
*|2351,2352
MCHC|2353,2357
-|2357,2358
32.1|2358,2362
RDW|2363,2366
-|2366,2367
13.7|2367,2371
Plt|2372,2375
_|2376,2377
_|2377,2378
_|2378,2379
<EOL>|2379,2380
_|2380,2381
_|2381,2382
_|2382,2383
07|2384,2386
:|2386,2387
20AM|2387,2391
BLOOD|2392,2397
_|2398,2399
_|2399,2400
_|2400,2401
PTT|2402,2405
-|2405,2406
42|2406,2408
.|2408,2409
0|2409,2410
*|2410,2411
_|2412,2413
_|2413,2414
_|2414,2415
<EOL>|2415,2416
_|2416,2417
_|2417,2418
_|2418,2419
07|2420,2422
:|2422,2423
20AM|2423,2427
BLOOD|2428,2433
Glucose|2434,2441
-|2441,2442
96|2442,2444
UreaN|2445,2450
-|2450,2451
7|2451,2452
Creat|2453,2458
-|2458,2459
0.4|2459,2462
Na|2463,2465
-|2465,2466
125|2466,2469
*|2469,2470
<EOL>|2471,2472
K|2472,2473
-|2473,2474
4.4|2474,2477
Cl|2478,2480
-|2480,2481
90|2481,2483
*|2483,2484
HCO3|2485,2489
-|2489,2490
30|2490,2492
AnGap|2493,2498
-|2498,2499
9|2499,2500
<EOL>|2500,2501
_|2501,2502
_|2502,2503
_|2503,2504
07|2505,2507
:|2507,2508
20AM|2508,2512
BLOOD|2513,2518
ALT|2519,2522
-|2522,2523
35|2523,2525
AST|2526,2529
-|2529,2530
131|2530,2533
*|2533,2534
LD|2535,2537
(|2537,2538
_|2538,2539
_|2539,2540
_|2540,2541
)|2541,2542
-|2542,2543
265|2543,2546
*|2546,2547
AlkPhos|2548,2555
-|2555,2556
184|2556,2559
*|2559,2560
<EOL>|2561,2562
TotBili|2562,2569
-|2569,2570
1|2570,2571
.|2571,2572
9|2572,2573
*|2573,2574
<EOL>|2574,2575
_|2575,2576
_|2576,2577
_|2577,2578
07|2579,2581
:|2581,2582
20AM|2582,2586
BLOOD|2587,2592
Albumin|2593,2600
-|2600,2601
2|2601,2602
.|2602,2603
5|2603,2604
*|2604,2605
Calcium|2606,2613
-|2613,2614
7|2614,2615
.|2615,2616
2|2616,2617
*|2617,2618
Phos|2619,2623
-|2623,2624
2|2624,2625
.|2625,2626
6|2626,2627
*|2627,2628
<EOL>|2629,2630
Mg|2630,2632
-|2632,2633
2.0|2633,2636
<EOL>|2636,2637
<EOL>|2637,2638
Micro|2638,2643
Data|2644,2648
:|2648,2649
<EOL>|2649,2650
<EOL>|2650,2651
_|2651,2652
_|2652,2653
_|2653,2654
PERITONEAL|2655,2665
FLUID|2666,2671
GRAM|2672,2676
STAIN|2677,2682
-|2682,2683
negative|2684,2692
;|2692,2693
FLUID|2694,2699
<EOL>|2700,2701
CULTURE|2701,2708
-|2708,2709
PENDING|2709,2716
;|2716,2717
ANAEROBIC|2718,2727
CULTURE|2728,2735
-|2735,2736
negative|2737,2745
<EOL>|2745,2746
_|2746,2747
_|2747,2748
_|2748,2749
STOOL|2750,2755
CLOSTRIDIUM|2756,2767
DIFFICILE|2768,2777
TOXIN|2778,2783
A|2784,2785
&|2786,2787
B|2788,2789
<EOL>|2790,2791
TEST|2791,2795
-|2795,2796
negative|2797,2805
<EOL>|2805,2806
_|2806,2807
_|2807,2808
_|2808,2809
URINE|2810,2815
URINE|2816,2821
CULTURE|2822,2829
-|2829,2830
negative|2831,2839
<EOL>|2839,2840
_|2840,2841
_|2841,2842
_|2842,2843
SWAB|2844,2848
R|2849,2850
/|2850,2851
O|2851,2852
VANCOMYCIN|2853,2863
RESISTANT|2864,2873
ENTEROCOCCUS|2874,2886
-|2886,2887
<EOL>|2888,2889
negative|2889,2897
<EOL>|2897,2898
_|2898,2899
_|2899,2900
_|2900,2901
STOOL|2902,2907
CLOSTRIDIUM|2908,2919
DIFFICILE|2920,2929
TOXIN|2930,2935
A|2936,2937
&|2938,2939
B|2940,2941
<EOL>|2942,2943
TEST|2943,2947
-|2947,2948
negative|2949,2957
<EOL>|2957,2958
_|2958,2959
_|2959,2960
_|2960,2961
FLUID|2962,2967
RECEIVED|2968,2976
IN|2977,2979
BLOOD|2980,2985
CULTURE|2986,2993
BOTTLES|2994,3001
<EOL>|3002,3003
Fluid|3003,3008
Culture|3009,3016
in|3017,3019
Bottles|3020,3027
-|3027,3028
negative|3029,3037
<EOL>|3037,3038
_|3038,3039
_|3039,3040
_|3040,3041
PERITONEAL|3042,3052
FLUID|3053,3058
GRAM|3059,3063
STAIN|3064,3069
-|3069,3070
FINAL|3070,3075
;|3075,3076
FLUID|3077,3082
<EOL>|3083,3084
CULTURE|3084,3091
-|3091,3092
FINAL|3092,3097
;|3097,3098
ANAEROBIC|3099,3108
CULTURE|3109,3116
-|3116,3117
negative|3118,3126
<EOL>|3126,3127
_|3127,3128
_|3128,3129
_|3129,3130
BLOOD|3131,3136
CULTURE|3137,3144
Blood|3145,3150
Culture|3151,3158
,|3158,3159
Routine|3160,3167
-|3167,3168
<EOL>|3169,3170
negative|3170,3178
<EOL>|3179,3180
_|3180,3181
_|3181,3182
_|3182,3183
BLOOD|3184,3189
CULTURE|3190,3197
Blood|3198,3203
Culture|3204,3211
,|3211,3212
<EOL>|3213,3214
Routine|3214,3221
-|3221,3222
negative|3222,3230
<EOL>|3231,3232
_|3232,3233
_|3233,3234
_|3234,3235
URINE|3236,3241
URINE|3242,3247
CULTURE|3248,3255
-|3255,3256
FINAL|3256,3261
{|3262,3263
GRAM|3263,3267
POSITIVE|3268,3276
<EOL>|3277,3278
BACTERIA|3278,3286
}|3286,3287
INPATIENT|3288,3297
<EOL>|3298,3299
_|3299,3300
_|3300,3301
_|3301,3302
FLUID|3303,3308
RECEIVED|3309,3317
IN|3318,3320
BLOOD|3321,3326
CULTURE|3327,3334
BOTTLES|3335,3342
<EOL>|3343,3344
negative|3344,3352
<EOL>|3352,3353
<EOL>|3353,3354
Imaging|3354,3361
Results|3362,3369
:|3369,3370
<EOL>|3370,3371
<EOL>|3371,3372
CTA|3372,3375
(|3376,3377
_|3377,3378
_|3378,3379
_|3379,3380
)|3380,3381
:|3381,3382
<EOL>|3382,3383
1|3383,3384
.|3384,3385
No|3386,3388
evidence|3389,3397
of|3398,3400
pulmonary|3401,3410
embolism|3411,3419
.|3419,3420
<EOL>|3421,3422
2.|3422,3424
Stable|3425,3431
atelectasis|3432,3443
at|3444,3446
the|3447,3450
right|3451,3456
lung|3457,3461
base|3462,3466
.|3466,3467
<EOL>|3468,3469
3.|3469,3471
Moderate|3472,3480
right|3481,3486
and|3487,3490
small|3491,3496
left|3497,3501
pleural|3502,3509
effusions|3510,3519
,|3519,3520
unchanged|3521,3530
.|3530,3531
<EOL>|3532,3533
<EOL>|3533,3534
CTAP|3534,3538
(|3539,3540
_|3540,3541
_|3541,3542
_|3542,3543
)|3543,3544
:|3544,3545
<EOL>|3545,3546
1.|3546,3548
Hepatomegaly|3549,3561
and|3562,3565
large|3566,3571
ascites|3572,3579
consistent|3580,3590
with|3591,3595
stated|3596,3602
history|3603,3610
<EOL>|3611,3612
of|3612,3614
liver|3615,3620
<EOL>|3621,3622
disease|3622,3629
.|3629,3630
No|3631,3633
evidence|3634,3642
of|3643,3645
portal|3646,3652
venous|3653,3659
thrombosis|3660,3670
suggesting|3671,3681
that|3682,3686
<EOL>|3687,3688
the|3688,3691
findings|3692,3700
on|3701,3703
the|3704,3707
prior|3708,3713
ultrasound|3714,3724
may|3725,3728
have|3729,3733
resulted|3734,3742
from|3743,3747
<EOL>|3748,3749
extremely|3749,3758
slow|3759,3763
/|3764,3765
undetectable|3766,3778
flow|3779,3783
.|3783,3784
<EOL>|3786,3787
2.|3787,3789
Moderate|3790,3798
right|3799,3804
and|3805,3808
small|3809,3814
left|3815,3819
pleural|3820,3827
effusions|3828,3837
,|3837,3838
increased|3839,3848
on|3849,3851
<EOL>|3852,3853
the|3853,3856
right|3857,3862
<EOL>|3863,3864
with|3864,3868
right|3869,3874
basilar|3875,3882
atelectasis|3883,3894
.|3894,3895
<EOL>|3896,3897
3.|3897,3899
Replaced|3900,3908
right|3909,3914
hepatic|3915,3922
artery|3923,3929
arising|3930,3937
from|3938,3942
the|3943,3946
SMA|3947,3950
,|3950,3951
otherwise|3952,3961
<EOL>|3962,3963
conventional|3963,3975
arterial|3976,3984
and|3985,3988
venous|3989,3995
anatomy|3996,4003
.|4003,4004
<EOL>|4004,4005
<EOL>|4006,4007
This|4030,4034
is|4035,4037
a|4038,4039
_|4040,4041
_|4041,4042
_|4042,4043
woman|4044,4049
with|4050,4054
likely|4055,4061
alcoholic|4062,4071
hepatitis|4072,4081
and|4082,4085
<EOL>|4086,4087
recurrent|4087,4096
ascites|4097,4104
who|4105,4108
is|4109,4111
admitted|4112,4120
with|4121,4125
low|4126,4129
-|4129,4130
grade|4130,4135
fevers|4136,4142
,|4142,4143
high|4144,4148
<EOL>|4149,4150
white|4150,4155
count|4156,4161
,|4161,4162
and|4163,4166
abdominal|4167,4176
pain|4177,4181
.|4181,4182
<EOL>|4182,4183
<EOL>|4184,4185
#|4185,4186
ASCITES|4187,4194
/|4194,4195
ALC|4195,4198
HEPATITIS|4199,4208
/|4208,4209
LEUKOCYTOSIS|4209,4221
:|4221,4222
Patient|4223,4230
with|4231,4235
fatty|4236,4241
liver|4242,4247
<EOL>|4248,4249
and|4249,4252
ascites|4253,4260
in|4261,4263
setting|4264,4271
of|4272,4274
extensive|4275,4284
drinking|4285,4293
history|4294,4301
and|4302,4305
AST|4306,4309
/|4309,4310
ALT|4310,4313
<EOL>|4314,4315
elevation|4315,4324
>|4325,4326
2|4326,4327
.|4327,4328
Discriminant|4329,4341
function|4342,4350
on|4351,4353
admission|4354,4363
was|4364,4367
~|4368,4369
30|4369,4371
.|4371,4372
<EOL>|4374,4375
Patient|4375,4382
had|4383,4386
a|4387,4388
paracentesis|4389,4401
on|4402,4404
_|4405,4406
_|4406,4407
_|4407,4408
and|4409,4412
4L|4413,4415
was|4416,4419
removed|4420,4427
;|4427,4428
<EOL>|4429,4430
peritoneal|4430,4440
fluid|4441,4446
was|4447,4450
negative|4451,4459
for|4460,4463
SBP|4464,4467
.|4467,4468
Diuretics|4469,4478
were|4479,4483
initially|4484,4493
<EOL>|4494,4495
held|4495,4499
in|4500,4502
the|4503,4506
setting|4507,4514
of|4515,4517
hyponatremia|4518,4530
.|4530,4531
She|4532,4535
was|4536,4539
treated|4540,4547
<EOL>|4548,4549
supportively|4549,4561
with|4562,4566
nutrition|4567,4576
,|4576,4577
brief|4578,4583
antibiotics|4584,4595
for|4596,4599
urinary|4600,4607
tract|4608,4613
<EOL>|4614,4615
infection|4615,4624
(|4625,4626
3|4626,4627
-|4627,4628
days|4628,4632
of|4633,4635
ceftriaxone|4636,4647
)|4647,4648
,|4648,4649
and|4650,4653
therapeutic|4654,4665
paracenteses|4666,4678
<EOL>|4679,4680
x3|4680,4682
.|4682,4683
Her|4684,4687
symptoms|4688,4696
,|4696,4697
white|4698,4703
cell|4704,4708
count|4709,4714
,|4714,4715
and|4716,4719
total|4720,4725
bilirubin|4726,4735
were|4736,4740
<EOL>|4741,4742
improving|4742,4751
at|4752,4754
time|4755,4759
of|4760,4762
discharge|4763,4772
.|4772,4773
She|4774,4777
will|4778,4782
follow|4783,4789
-|4789,4790
up|4790,4792
with|4793,4797
Dr|4798,4800
.|4800,4801
<EOL>|4802,4803
_|4803,4804
_|4804,4805
_|4805,4806
in|4807,4809
liver|4810,4815
clinic|4816,4822
and|4823,4826
with|4827,4831
her|4832,4835
primary|4836,4843
care|4844,4848
provider|4849,4857
,|4857,4858
Dr|4859,4861
.|4861,4862
<EOL>|4863,4864
_|4864,4865
_|4865,4866
_|4866,4867
,|4867,4868
in|4869,4871
two|4872,4875
weeks|4876,4881
.|4881,4882
<EOL>|4883,4884
<EOL>|4884,4885
#|4885,4886
HYPONATREMIA|4887,4899
:|4899,4900
Likely|4901,4907
hypovolemic|4908,4919
hyponatremia|4920,4932
with|4933,4937
some|4938,4942
<EOL>|4943,4944
component|4944,4953
of|4954,4956
euvolemic|4957,4966
hyponatremia|4967,4979
from|4980,4984
liver|4985,4990
disease|4991,4998
.|4998,4999
Her|5000,5003
<EOL>|5004,5005
spironlactone|5005,5018
was|5019,5022
held|5023,5027
and|5028,5031
can|5032,5035
be|5036,5038
restarted|5039,5048
at|5049,5051
the|5052,5055
discretion|5056,5066
of|5067,5069
<EOL>|5070,5071
her|5071,5074
outpatient|5075,5085
liver|5086,5091
team|5092,5096
,|5096,5097
if|5098,5100
necessary|5101,5110
.|5110,5111
Sodium|5112,5118
at|5119,5121
time|5122,5126
of|5127,5129
<EOL>|5130,5131
discharge|5131,5140
was|5141,5144
125|5145,5148
.|5148,5149
She|5150,5153
has|5154,5157
been|5158,5162
advised|5163,5170
to|5171,5173
continue|5174,5182
a|5183,5184
low|5185,5188
sodium|5189,5195
<EOL>|5196,5197
diet|5197,5201
and|5202,5205
free|5206,5210
water|5211,5216
restriction|5217,5228
to|5229,5231
_|5232,5233
_|5233,5234
_|5234,5235
liters|5236,5242
daily|5243,5248
.|5248,5249
<EOL>|5249,5250
<EOL>|5251,5252
#|5252,5253
ALCOHOLISM|5254,5264
:|5264,5265
Patient|5266,5273
has|5274,5277
been|5278,5282
trying|5283,5289
to|5290,5292
cut|5293,5296
back|5297,5301
recently|5302,5310
,|5310,5311
but|5312,5315
<EOL>|5316,5317
reports|5317,5324
daily|5325,5330
heavy|5331,5336
alcohol|5337,5344
intake|5345,5351
for|5352,5355
the|5356,5359
past|5360,5364
_|5365,5366
_|5366,5367
_|5367,5368
years|5369,5374
;|5374,5375
she|5376,5379
has|5380,5383
<EOL>|5384,5385
had|5385,5388
withdrawal|5389,5399
symptoms|5400,5408
before|5409,5415
but|5416,5419
no|5420,5422
seizures|5423,5431
.|5431,5432
Shakes|5433,5439
and|5440,5443
<EOL>|5444,5445
hallucinations|5445,5459
.|5459,5460
Reports|5462,5469
sobriety|5470,5478
since|5479,5484
prior|5485,5490
admission|5491,5500
.|5500,5501
She|5502,5505
<EOL>|5506,5507
will|5507,5511
continue|5512,5520
outpatient|5521,5531
rehab|5532,5537
.|5537,5538
<EOL>|5538,5539
<EOL>|5541,5542
#|5542,5543
URINARY|5544,5551
TRACT|5552,5557
INFECTION|5558,5567
:|5567,5568
she|5569,5572
was|5573,5576
treated|5577,5584
with|5585,5589
a|5590,5591
three|5592,5597
-|5597,5598
day|5598,5601
<EOL>|5602,5603
course|5603,5609
of|5610,5612
empiric|5613,5620
ceftriaxone|5621,5632
for|5633,5636
concern|5637,5644
of|5645,5647
UTI|5648,5651
.|5651,5652
<EOL>|5652,5653
<EOL>|5653,5654
#|5654,5655
BACK|5656,5660
PAIN|5661,5665
/|5665,5666
ABDOMINAL|5666,5675
PAIN|5676,5680
:|5680,5681
this|5682,5686
was|5687,5690
treated|5691,5698
in|5699,5701
house|5702,5707
with|5708,5712
<EOL>|5713,5714
lidocaine|5714,5723
patches|5724,5731
as|5732,5734
needed|5735,5741
and|5742,5745
oxycodone|5746,5755
as|5756,5758
needed|5759,5765
.|5765,5766
She|5767,5770
has|5771,5774
<EOL>|5775,5776
been|5776,5780
provided|5781,5789
with|5790,5794
a|5795,5796
short|5797,5802
course|5803,5809
of|5810,5812
Tramadol|5813,5821
to|5822,5824
take|5825,5829
as|5830,5832
needed|5833,5839
<EOL>|5840,5841
until|5841,5846
follow|5847,5853
-|5853,5854
up|5854,5856
with|5857,5861
her|5862,5865
primary|5866,5873
care|5874,5878
provider|5879,5887
.|5887,5888
She|5889,5892
understands|5893,5904
<EOL>|5905,5906
that|5906,5910
this|5911,5915
is|5916,5918
only|5919,5923
a|5924,5925
temporary|5926,5935
medication|5936,5946
and|5947,5950
will|5951,5955
be|5956,5958
<EOL>|5959,5960
discontinued|5960,5972
when|5973,5977
her|5978,5981
acute|5982,5987
hepatitis|5988,5997
resolves|5998,6006
.|6006,6007
<EOL>|6007,6008
<EOL>|6008,6009
#|6009,6010
Prophylaxis|6011,6022
:|6022,6023
<EOL>|6025,6026
-|6026,6027
DVT|6027,6030
ppx|6031,6034
with|6035,6039
SC|6040,6042
heparin|6043,6050
<EOL>|6052,6053
-|6053,6054
Bowel|6054,6059
regimen|6060,6067
with|6068,6072
lactulose|6073,6082
,|6082,6083
no|6084,6086
PPI|6087,6090
<EOL>|6092,6093
-|6093,6094
Pain|6094,6098
management|6099,6109
with|6110,6114
oxycodone|6115,6124
and|6125,6128
lidocaine|6129,6138
patch|6139,6144
<EOL>|6146,6147
#|6147,6148
Communication|6149,6162
:|6162,6163
Patient|6164,6171
<EOL>|6173,6174
#|6174,6175
Code|6176,6180
:|6180,6181
presumed|6182,6190
full|6191,6195
<EOL>|6195,6196
<EOL>|6197,6198
Medications|6198,6209
on|6210,6212
Admission|6213,6222
:|6222,6223
<EOL>|6223,6224
Multivitamin|6224,6236
,|6236,6237
thiamine|6238,6246
,|6246,6247
folate|6248,6254
,|6254,6255
spironolactone|6256,6270
25mg|6271,6275
daily|6276,6281
,|6281,6282
<EOL>|6283,6284
lidocaine|6284,6293
patch|6294,6299
prn|6300,6303
,|6303,6304
nicotine|6305,6313
patch|6314,6319
.|6319,6320
<EOL>|6320,6321
<EOL>|6322,6323
Discharge|6323,6332
Medications|6333,6344
:|6344,6345
<EOL>|6345,6346
1.|6346,6348
Multivitamin|6349,6361
Tablet|6366,6372
Sig|6373,6376
:|6376,6377
One|6378,6381
(|6382,6383
1|6383,6384
)|6384,6385
Tablet|6386,6392
PO|6393,6395
DAILY|6396,6401
(|6402,6403
Daily|6403,6408
)|6408,6409
.|6409,6410
<EOL>|6411,6412
<EOL>|6413,6414
2.|6414,6416
Thiamine|6417,6425
HCl|6426,6429
100|6430,6433
mg|6434,6436
Tablet|6437,6443
Sig|6444,6447
:|6447,6448
One|6449,6452
(|6453,6454
1|6454,6455
)|6455,6456
Tablet|6457,6463
PO|6464,6466
DAILY|6467,6472
<EOL>|6473,6474
(|6474,6475
Daily|6475,6480
)|6480,6481
.|6481,6482
<EOL>|6484,6485
3.|6485,6487
Folic|6488,6493
Acid|6494,6498
1|6499,6500
mg|6501,6503
Tablet|6504,6510
Sig|6511,6514
:|6514,6515
One|6516,6519
(|6520,6521
1|6521,6522
)|6522,6523
Tablet|6524,6530
PO|6531,6533
DAILY|6534,6539
(|6540,6541
Daily|6541,6546
)|6546,6547
.|6547,6548
<EOL>|6550,6551
<EOL>|6551,6552
4.|6552,6554
Nicotine|6555,6563
14|6564,6566
mg|6567,6569
/|6569,6570
24|6570,6572
hr|6573,6575
Patch|6576,6581
24|6582,6584
hr|6585,6587
Sig|6588,6591
:|6591,6592
One|6593,6596
(|6597,6598
1|6598,6599
)|6599,6600
Patch|6601,6606
24|6607,6609
hr|6610,6612
<EOL>|6613,6614
Transdermal|6614,6625
DAILY|6626,6631
(|6632,6633
Daily|6633,6638
)|6638,6639
.|6639,6640
<EOL>|6642,6643
5.|6643,6645
Lidocaine|6646,6655
5|6656,6657
%|6658,6659
(|6659,6660
700|6660,6663
mg|6664,6666
/|6666,6667
patch|6667,6672
)|6672,6673
Adhesive|6674,6682
Patch|6683,6688
,|6688,6689
Medicated|6690,6699
Sig|6700,6703
:|6703,6704
<EOL>|6705,6706
One|6706,6709
(|6710,6711
1|6711,6712
)|6712,6713
Adhesive|6714,6722
Patch|6723,6728
,|6728,6729
Medicated|6730,6739
Topical|6740,6747
DAILY|6748,6753
(|6754,6755
Daily|6755,6760
)|6760,6761
.|6761,6762
<EOL>|6764,6765
6.|6765,6767
Tramadol|6768,6776
50|6777,6779
mg|6780,6782
Tablet|6783,6789
Sig|6790,6793
:|6793,6794
One|6795,6798
(|6799,6800
1|6800,6801
)|6801,6802
Tablet|6803,6809
PO|6810,6812
every|6813,6818
eight|6819,6824
(|6825,6826
8|6826,6827
)|6827,6828
<EOL>|6829,6830
hours|6830,6835
as|6836,6838
needed|6839,6845
for|6846,6849
pain|6850,6854
.|6854,6855
<EOL>|6855,6856
Disp|6856,6860
:|6860,6861
*|6861,6862
30|6862,6864
Tablet|6865,6871
(|6871,6872
s|6872,6873
)|6873,6874
*|6874,6875
Refills|6876,6883
:|6883,6884
*|6884,6885
0|6885,6886
*|6886,6887
<EOL>|6887,6888
<EOL>|6888,6889
<EOL>|6890,6891
Discharge|6891,6900
Disposition|6901,6912
:|6912,6913
<EOL>|6913,6914
Home|6914,6918
<EOL>|6918,6919
<EOL>|6920,6921
Discharge|6921,6930
Diagnosis|6931,6940
:|6940,6941
<EOL>|6941,6942
Primary|6942,6949
diagnosis|6950,6959
:|6959,6960
Alcoholic|6961,6970
hepatitis|6971,6980
.|6980,6981
<EOL>|6981,6982
<EOL>|6983,6984
Mental|7005,7011
Status|7012,7018
:|7018,7019
Clear|7020,7025
and|7026,7029
coherent|7030,7038
.|7038,7039
<EOL>|7039,7040
Level|7040,7045
of|7046,7048
Consciousness|7049,7062
:|7062,7063
Alert|7064,7069
and|7070,7073
interactive|7074,7085
.|7085,7086
<EOL>|7086,7087
Activity|7087,7095
Status|7096,7102
:|7102,7103
Ambulatory|7104,7114
-|7115,7116
Independent|7117,7128
.|7128,7129
<EOL>|7129,7130
<EOL>|7131,7132
You|7156,7159
were|7160,7164
admitted|7165,7173
to|7174,7176
the|7177,7180
hospital|7181,7189
for|7190,7193
alcoholic|7194,7203
hepatitis|7204,7213
.|7213,7214
This|7215,7219
<EOL>|7220,7221
is|7221,7223
a|7224,7225
condition|7226,7235
in|7236,7238
which|7239,7244
your|7245,7249
liver|7250,7255
becomes|7256,7263
inflamed|7264,7272
due|7273,7276
to|7277,7279
<EOL>|7280,7281
excessive|7281,7290
alcohol|7291,7298
intake|7299,7305
.|7305,7306
You|7307,7310
were|7311,7315
also|7316,7320
noted|7321,7326
to|7327,7329
have|7330,7334
an|7335,7337
<EOL>|7338,7339
elevated|7339,7347
white|7348,7353
cell|7354,7358
count|7359,7364
which|7365,7370
can|7371,7374
sometimes|7375,7384
indicate|7385,7393
<EOL>|7394,7395
infection|7395,7404
.|7404,7405
You|7406,7409
were|7410,7414
treated|7415,7422
with|7423,7427
a|7428,7429
brief|7430,7435
course|7436,7442
of|7443,7445
antibiotics|7446,7457
<EOL>|7458,7459
for|7459,7462
a|7463,7464
urinary|7465,7472
tract|7473,7478
infection|7479,7488
.|7488,7489
Otherwise|7490,7499
your|7500,7504
blood|7505,7510
and|7511,7514
<EOL>|7515,7516
peritoneal|7516,7526
fluid|7527,7532
cultures|7533,7541
remain|7542,7548
negative|7549,7557
.|7557,7558
<EOL>|7558,7559
<EOL>|7559,7560
We|7560,7562
made|7563,7567
the|7568,7571
following|7572,7581
changes|7582,7589
to|7590,7592
your|7593,7597
medications|7598,7609
:|7609,7610
<EOL>|7611,7612
We|7612,7614
stopped|7615,7622
your|7623,7627
spironolactone|7628,7642
because|7643,7650
your|7651,7655
blood|7656,7661
sodium|7662,7668
levels|7669,7675
<EOL>|7676,7677
were|7677,7681
too|7682,7685
low|7686,7689
.|7689,7690
<EOL>|7690,7691
We|7691,7693
added|7694,7699
Tramadol|7700,7708
to|7709,7711
take|7712,7716
as|7717,7719
needed|7720,7726
for|7727,7730
back|7731,7735
pain|7736,7740
.|7740,7741
<EOL>|7742,7743
<EOL>|7744,7745
Followup|7745,7753
Instructions|7754,7766
:|7766,7767
<EOL>|7767,7768
_|7768,7769
_|7769,7770
_|7770,7771
<EOL>|7771,7772

