 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
SURGERY|156,163
<EOL>|163,164
<EOL>|165,166
Allergies|166,175
:|175,176
<EOL>|177,178
_|178,179
_|179,180
_|180,181
<EOL>|181,182
<EOL>|183,184
Attending|184,193
:|193,194
_|195,196
_|196,197
_|197,198
.|198,199
<EOL>|199,200
<EOL>|201,202
Chief|202,207
Complaint|208,217
:|217,218
<EOL>|218,219
Morbid|219,225
obesity|226,233
<EOL>|233,234
<EOL>|235,236
Major|236,241
Surgical|242,250
or|251,253
Invasive|254,262
Procedure|263,272
:|272,273
<EOL>|273,274
_|274,275
_|275,276
_|276,277
:|277,278
<EOL>|279,280
1.|280,282
Laparoscopic|283,295
repair|296,302
of|303,305
paraesophageal|306,320
hernia|321,327
.|327,328
<EOL>|328,329
2.|329,331
Laparoscopic|332,344
adjustable|345,355
gastric|356,363
band|364,368
.|368,369
<EOL>|369,370
<EOL>|370,371
<EOL>|372,373
History|373,380
of|381,383
Present|384,391
Illness|392,399
:|399,400
<EOL>|400,401
Per|401,404
Dr.|405,408
_|409,410
_|410,411
_|411,412
has|413,416
class|417,422
III|423,426
morbid|427,433
obesity|434,441
with|442,446
<EOL>|447,448
_|448,449
_|449,450
_|450,451
of|452,454
238.4|455,460
pounds|461,467
as|468,470
of|471,473
_|474,475
_|475,476
_|476,477
with|478,482
initial|483,490
screen|491,497
_|498,499
_|499,500
_|500,501
<EOL>|502,503
of|503,505
241.4|506,511
pounds|512,518
on|519,521
_|522,523
_|523,524
_|524,525
,|525,526
height|527,533
is|534,536
64|537,539
inches|540,546
and|547,550
BMI|551,554
of|555,557
40.9|558,562
.|562,563
<EOL>|564,565
Her|566,569
previous|570,578
_|579,580
_|580,581
_|581,582
loss|583,587
efforts|588,595
have|596,600
included|601,609
_|610,611
_|611,612
_|612,613
Watchers|614,622
,|622,623
<EOL>|624,625
_|625,626
_|626,627
_|627,628
Loss|629,633
,|633,634
Slim|635,639
-|639,640
Fast|640,644
,|644,645
over-the|646,654
-|654,655
counter|655,662
pancreatic|663,673
lipase|674,680
<EOL>|681,682
inhibitor|682,691
_|692,693
_|693,694
_|694,695
visits|696,702
.|702,703
She|705,708
has|709,712
lost|713,717
up|718,720
to|721,723
20|724,726
pounds|727,733
but|734,737
<EOL>|738,739
unable|739,745
to|746,748
maintain|749,757
the|758,761
_|762,763
_|763,764
_|764,765
.|765,766
Her|768,771
lowest|772,778
_|779,780
_|780,781
_|781,782
as|783,785
an|786,788
adult|789,794
<EOL>|795,796
was|796,799
180|800,803
pounds|804,810
and|811,814
her|815,818
highest|819,826
_|827,828
_|828,829
_|829,830
was|831,834
her|835,838
initial|839,846
screen|847,853
<EOL>|854,855
_|855,856
_|856,857
_|857,858
of|859,861
241.4|862,867
pounds|868,874
.|874,875
She|877,880
weighed|881,888
225.4|889,894
pounds|895,901
_|902,903
_|903,904
_|904,905
years|906,911
ago|912,915
<EOL>|916,917
and|917,920
235|921,924
pounds|925,931
one|932,935
year|936,940
ago|941,944
.|944,945
She|947,950
stated|951,957
that|958,962
she|963,966
has|967,970
been|971,975
<EOL>|976,977
struggling|977,987
with|988,992
_|993,994
_|994,995
_|995,996
since|997,1002
_|1003,1004
_|1004,1005
_|1005,1006
years|1007,1012
of|1013,1015
age|1016,1019
and|1020,1023
cites|1024,1029
as|1030,1032
<EOL>|1033,1034
factors|1034,1041
contributing|1042,1054
to|1055,1057
her|1058,1061
excess|1062,1068
_|1069,1070
_|1070,1071
_|1071,1072
genetics|1073,1081
,|1081,1082
inconsistent|1083,1095
<EOL>|1096,1097
meal|1097,1101
pattern|1102,1109
,|1109,1110
late|1111,1115
night|1116,1121
eating|1122,1128
,|1128,1129
large|1130,1135
portions|1136,1144
,|1144,1145
too|1146,1149
many|1150,1154
<EOL>|1155,1156
carbohydrates|1156,1169
,|1169,1170
grazing|1171,1178
and|1179,1182
emotional|1183,1192
eating|1193,1199
at|1200,1202
times|1203,1208
.|1208,1209
For|1211,1214
<EOL>|1215,1216
exercise|1216,1224
she|1225,1228
does|1229,1233
_|1234,1235
_|1235,1236
_|1236,1237
one|1238,1241
hour|1242,1246
_|1247,1248
_|1248,1249
_|1249,1250
times|1251,1256
per|1257,1260
week|1261,1265
,|1265,1266
elliptical|1267,1277
<EOL>|1278,1279
_|1279,1280
_|1280,1281
_|1281,1282
minutes|1283,1290
_|1291,1292
_|1292,1293
_|1293,1294
times|1295,1300
per|1301,1304
week|1305,1309
and|1310,1313
some|1314,1318
kettle|1319,1325
bell|1326,1330
training|1331,1339
.|1339,1340
<EOL>|1341,1342
She|1342,1345
denied|1346,1352
history|1353,1360
of|1361,1363
eating|1364,1370
disorders|1371,1380
and|1381,1384
does|1385,1389
have|1390,1394
depression|1395,1405
,|1405,1406
<EOL>|1406,1407
has|1407,1410
not|1411,1414
been|1415,1419
seen|1420,1424
by|1425,1427
a|1428,1429
therapist|1430,1439
nor|1440,1443
has|1444,1447
she|1448,1451
been|1452,1456
hospitalized|1457,1469
<EOL>|1470,1471
for|1471,1474
any|1475,1478
mental|1479,1485
health|1486,1492
issues|1493,1499
and|1500,1503
she|1504,1507
is|1508,1510
not|1511,1514
on|1515,1517
any|1518,1521
psychotropic|1522,1534
<EOL>|1535,1536
medications|1536,1547
at|1548,1550
this|1551,1555
time|1556,1560
.|1560,1561
<EOL>|1561,1562
<EOL>|1562,1563
<EOL>|1564,1565
Past|1565,1569
Medical|1570,1577
History|1578,1585
:|1585,1586
<EOL>|1586,1587
PMHx|1587,1591
:|1591,1592
Hyperlipidemia|1593,1607
and|1608,1611
with|1612,1616
elevated|1617,1625
triglyceride|1626,1638
,|1638,1639
iron|1640,1644
<EOL>|1644,1645
deficiency|1645,1655
anemia|1656,1662
,|1662,1663
irritable|1664,1673
bowel|1674,1679
syndrome|1680,1688
,|1688,1689
allergic|1690,1698
rhinitis|1699,1707
,|1707,1708
<EOL>|1708,1709
dysmenorrhea|1709,1721
,|1721,1722
vitamin|1723,1730
D|1731,1732
deficiency|1733,1743
,|1743,1744
question|1745,1753
of|1754,1756
hypothyroidism|1757,1771
<EOL>|1771,1772
with|1772,1776
elevated|1777,1785
TSH|1786,1789
level|1790,1795
,|1795,1796
thalassemia|1797,1808
trait|1809,1814
,|1814,1815
fatty|1816,1821
liver|1822,1827
and|1828,1831
<EOL>|1831,1832
cholelithiasis|1832,1846
by|1847,1849
ultrasound|1850,1860
study|1861,1866
.|1866,1867
A|1868,1869
history|1870,1877
of|1878,1880
kissing|1881,1888
tonsils|1889,1896
<EOL>|1896,1897
that|1897,1901
was|1902,1905
associated|1906,1916
with|1917,1921
obstructive|1922,1933
sleep|1934,1939
apnea|1940,1945
and|1946,1949
<EOL>|1949,1950
gastroesophageal|1950,1966
reflux|1967,1973
,|1973,1974
these|1975,1980
have|1981,1985
resolved|1986,1994
completely|1995,2005
after|2006,2011
<EOL>|2012,2013
the|2013,2016
<EOL>|2016,2017
tonsillectomy|2017,2030
in|2031,2033
_|2034,2035
_|2035,2036
_|2036,2037
.|2037,2038
History|2039,2046
of|2047,2049
polycystic|2050,2060
ovary|2061,2066
<EOL>|2066,2067
syndrome|2067,2075
<EOL>|2075,2076
<EOL>|2077,2078
Family|2078,2084
History|2085,2092
:|2092,2093
<EOL>|2093,2094
bladder|2094,2101
CA|2102,2104
;|2104,2105
with|2106,2110
diabetes|2111,2119
,|2119,2120
breast|2121,2127
neoplasia|2128,2137
,|2137,2138
colon|2139,2144
CA|2145,2147
,|2147,2148
ovarian|2149,2156
<EOL>|2157,2158
CA|2158,2160
and|2161,2164
sarcoma|2165,2172
<EOL>|2172,2173
<EOL>|2174,2175
Physical|2175,2183
Exam|2184,2188
:|2188,2189
<EOL>|2189,2190
VSS|2190,2193
<EOL>|2193,2194
Constitutional|2194,2208
:|2208,2209
NAD|2210,2213
<EOL>|2213,2214
Neuro|2214,2219
:|2219,2220
Alert|2221,2226
and|2227,2230
oriented|2231,2239
x|2240,2241
3|2242,2243
<EOL>|2243,2244
Cardiac|2244,2251
:|2251,2252
RRR|2253,2256
,|2256,2257
NL|2258,2260
S1|2261,2263
,|2263,2264
S2|2264,2266
<EOL>|2266,2267
Lungs|2267,2272
:|2272,2273
CTA|2274,2277
B|2278,2279
<EOL>|2279,2280
Abd|2280,2283
:|2283,2284
Obese|2285,2290
,|2290,2291
soft|2292,2296
,|2296,2297
non-distened|2298,2310
,|2310,2311
appropriate|2312,2323
_|2324,2325
_|2325,2326
_|2326,2327
<EOL>|2328,2329
tenderness|2329,2339
,|2339,2340
no|2341,2343
rebound|2344,2351
tenderness|2352,2362
/|2362,2363
guarding|2363,2371
<EOL>|2371,2372
Wounds|2372,2378
:|2378,2379
Abd|2380,2383
lap|2384,2387
sites|2388,2393
with|2394,2398
primary|2399,2406
dsg|2407,2410
,|2410,2411
slight|2412,2418
serosanguinous|2419,2433
<EOL>|2434,2435
staining|2435,2443
x|2444,2445
1|2446,2447
,|2447,2448
no|2449,2451
periwound|2452,2461
erythema|2462,2470
<EOL>|2470,2471
Ext|2471,2474
:|2474,2475
No|2476,2478
edema|2479,2484
<EOL>|2484,2485
<EOL>|2486,2487
Pertinent|2487,2496
Results|2497,2504
:|2504,2505
<EOL>|2505,2506
LABS|2506,2510
:|2510,2511
<EOL>|2511,2512
_|2512,2513
_|2513,2514
_|2514,2515
09|2516,2518
:|2518,2519
20AM|2519,2523
BLOOD|2524,2529
WBC|2530,2533
-|2533,2534
9.8|2534,2537
RBC|2538,2541
-|2541,2542
5|2542,2543
.|2543,2544
19|2544,2546
Hgb|2547,2550
-|2550,2551
14.0|2551,2555
Hct|2556,2559
-|2559,2560
41.9|2560,2564
<EOL>|2565,2566
MCV|2566,2569
-|2569,2570
81|2570,2572
*|2572,2573
MCH|2574,2577
-|2577,2578
27.0|2578,2582
MCHC|2583,2587
-|2587,2588
33.5|2588,2592
RDW|2593,2596
-|2596,2597
13.5|2597,2601
Plt|2602,2605
_|2606,2607
_|2607,2608
_|2608,2609
<EOL>|2609,2610
_|2610,2611
_|2611,2612
_|2612,2613
09|2614,2616
:|2616,2617
20AM|2617,2621
BLOOD|2622,2627
Plt|2628,2631
_|2632,2633
_|2633,2634
_|2634,2635
<EOL>|2635,2636
<EOL>|2636,2637
_|2637,2638
_|2638,2639
_|2639,2640
UGI|2641,2644
SGL|2645,2648
CONTRAST|2649,2657
W|2658,2659
/|2659,2660
KUB|2661,2664
:|2664,2665
<EOL>|2665,2666
IMPRESSION|2666,2676
:|2676,2677
Slightly|2678,2686
horizontally|2687,2699
positioned|2700,2710
lap|2711,2714
band|2715,2719
with|2720,2724
a|2725,2726
<EOL>|2727,2728
patent|2728,2734
stoma|2735,2740
and|2741,2744
no|2745,2747
evidence|2748,2756
of|2757,2759
leak|2760,2764
.|2764,2765
<EOL>|2766,2767
<EOL>|2767,2768
<EOL>|2769,2770
Brief|2770,2775
Hospital|2776,2784
Course|2785,2791
:|2791,2792
<EOL>|2792,2793
Ms.|2793,2796
_|2797,2798
_|2798,2799
_|2799,2800
presented|2801,2810
to|2811,2813
_|2814,2815
_|2815,2816
_|2816,2817
on|2818,2820
_|2821,2822
_|2822,2823
_|2823,2824
.|2824,2825
Pt|2826,2828
was|2829,2832
<EOL>|2833,2834
evaluated|2834,2843
by|2844,2846
anaesthesia|2847,2858
and|2859,2862
taken|2863,2868
to|2869,2871
the|2872,2875
operating|2876,2885
room|2886,2890
where|2891,2896
<EOL>|2897,2898
she|2898,2901
underwent|2902,2911
a|2912,2913
laparoscopic|2914,2926
adjustable|2927,2937
gastric|2938,2945
band|2946,2950
placement|2951,2960
<EOL>|2961,2962
and|2962,2965
repair|2966,2972
of|2973,2975
paraesophageal|2976,2990
hernia|2991,2997
.|2997,2998
There|2999,3004
were|3005,3009
no|3010,3012
adverse|3013,3020
<EOL>|3021,3022
events|3022,3028
in|3029,3031
the|3032,3035
operating|3036,3045
room|3046,3050
;|3050,3051
please|3052,3058
see|3059,3062
the|3063,3066
operative|3067,3076
note|3077,3081
for|3082,3085
<EOL>|3086,3087
details|3087,3094
.|3094,3095
Pt|3096,3098
was|3099,3102
extubated|3103,3112
,|3112,3113
taken|3114,3119
to|3120,3122
the|3123,3126
PACU|3127,3131
until|3132,3137
stable|3138,3144
,|3144,3145
then|3146,3150
<EOL>|3151,3152
transferred|3152,3163
to|3164,3166
the|3167,3170
ward|3171,3175
for|3176,3179
observation|3180,3191
.|3191,3192
<EOL>|3193,3194
<EOL>|3194,3195
Post-operatively|3195,3211
,|3211,3212
the|3213,3216
patient|3217,3224
remained|3225,3233
afebrile|3234,3242
with|3243,3247
stable|3248,3254
<EOL>|3255,3256
vital|3256,3261
signs|3262,3267
.|3267,3268
The|3270,3273
patient|3274,3281
|3281,3282
s|3282,3283
pain|3284,3288
was|3289,3292
well|3293,3297
controlled|3298,3308
with|3309,3313
oral|3314,3318
<EOL>|3319,3320
Roxicet|3320,3327
prn|3328,3331
.|3331,3332
The|3334,3337
patient|3338,3345
remained|3346,3354
stable|3355,3361
from|3362,3366
both|3367,3371
a|3372,3373
<EOL>|3374,3375
cardiovascular|3375,3389
and|3390,3393
pulmonary|3394,3403
standpoint|3404,3414
;|3414,3415
she|3416,3419
was|3420,3423
maintained|3424,3434
on|3435,3437
<EOL>|3438,3439
CPAP|3439,3443
overnight|3444,3453
for|3454,3457
known|3458,3463
sleep|3464,3469
apnea|3470,3475
.|3475,3476
The|3478,3481
patient|3482,3489
was|3490,3493
initially|3494,3503
<EOL>|3504,3505
on|3505,3507
a|3508,3509
bariatric|3510,3519
stage|3520,3525
1|3526,3527
diet|3528,3532
,|3532,3533
but|3534,3537
was|3538,3541
made|3542,3546
NPO|3547,3550
at|3551,3553
_|3554,3555
_|3555,3556
_|3556,3557
POD1|3558,3562
for|3563,3566
an|3567,3569
<EOL>|3570,3571
UGI|3571,3574
series|3575,3581
.|3581,3582
The|3584,3587
UGI|3588,3591
was|3592,3595
negative|3596,3604
for|3605,3608
leak|3609,3613
or|3614,3616
obstruction|3617,3628
,|3628,3629
<EOL>|3630,3631
therefore|3631,3640
,|3640,3641
the|3642,3645
patient|3646,3653
's|3653,3655
diet|3656,3660
advanced|3661,3669
sequentially|3670,3682
to|3683,3685
bariatric|3686,3695
<EOL>|3696,3697
stage|3697,3702
3|3703,3704
and|3705,3708
well|3709,3713
tolerated|3714,3723
;|3723,3724
pt|3725,3727
|3727,3728
s|3728,3729
intake|3730,3736
and|3737,3740
output|3741,3747
were|3748,3752
closely|3753,3760
<EOL>|3761,3762
monitored|3762,3771
.|3771,3772
Urine|3774,3779
output|3780,3786
remained|3787,3795
adequate|3796,3804
throughout|3805,3815
the|3816,3819
<EOL>|3820,3821
hospitalization|3821,3836
.|3836,3837
The|3839,3842
received|3843,3851
subcutaneous|3852,3864
heparin|3865,3872
and|3873,3876
venodyne|3877,3885
<EOL>|3886,3887
boots|3887,3892
were|3893,3897
used|3898,3902
during|3903,3909
admission|3910,3919
;|3919,3920
early|3921,3926
and|3927,3930
frequent|3931,3939
ambulation|3940,3950
<EOL>|3951,3952
were|3952,3956
strongly|3957,3965
encouraged|3966,3976
.|3976,3977
<EOL>|3977,3978
<EOL>|3978,3979
The|3979,3982
patient|3983,3990
was|3991,3994
subsequently|3995,4007
discharged|4008,4018
to|4019,4021
home|4022,4026
on|4027,4029
POD1|4030,4034
.|4034,4035
The|4037,4040
<EOL>|4041,4042
patient|4042,4049
received|4050,4058
discharge|4059,4068
teaching|4069,4077
and|4078,4081
follow|4082,4088
-|4088,4089
up|4089,4091
instructions|4092,4104
<EOL>|4105,4106
with|4106,4110
understanding|4111,4124
verbalized|4125,4135
and|4136,4139
agreement|4140,4149
with|4150,4154
the|4155,4158
discharge|4159,4168
<EOL>|4169,4170
plan|4170,4174
.|4174,4175
She|4176,4179
will|4180,4184
follow|4185,4191
-|4191,4192
up|4192,4194
with|4195,4199
Dr.|4200,4203
_|4204,4205
_|4205,4206
_|4206,4207
the|4208,4211
bariatric|4212,4221
<EOL>|4222,4223
dietitian|4223,4232
in|4233,4235
clinic|4236,4242
in|4243,4245
2|4246,4247
weeks|4248,4253
.|4253,4254
<EOL>|4254,4255
<EOL>|4255,4256
<EOL>|4257,4258
Medications|4258,4269
on|4270,4272
Admission|4273,4282
:|4282,4283
<EOL>|4283,4284
The|4284,4287
Preadmission|4288,4300
Medication|4301,4311
list|4312,4316
may|4317,4320
be|4321,4323
inaccurate|4324,4334
and|4335,4338
requires|4339,4347
<EOL>|4348,4349
futher|4349,4355
investigation|4356,4369
.|4369,4370
<EOL>|4370,4371
1.|4371,4373
Multivitamins|4374,4387
W|4388,4389
/|4389,4390
minerals|4390,4398
1|4399,4400
TAB|4401,4404
PO|4405,4407
DAILY|4408,4413
<EOL>|4414,4415
2.|4415,4417
Ascorbic|4418,4426
Acid|4427,4431
_|4432,4433
_|4433,4434
_|4434,4435
mg|4436,4438
PO|4439,4441
DAILY|4442,4447
<EOL>|4448,4449
3.|4449,4451
cholecalciferol|4452,4467
(|4468,4469
vitamin|4469,4476
D3|4477,4479
)|4479,4480
*|4481,4482
NF|4482,4484
*|4484,4485
3,000|4486,4491
unit|4492,4496
Oral|4497,4501
daily|4502,4507
<EOL>|4508,4509
4.|4509,4511
Cyclobenzaprine|4512,4527
_|4528,4529
_|4529,4530
_|4530,4531
mg|4532,4534
PO|4535,4537
TID|4538,4541
:|4541,4542
PRN|4542,4545
muscle|4546,4552
spasms|4553,4559
<EOL>|4560,4561
<EOL>|4561,4562
<EOL>|4563,4564
Discharge|4564,4573
Medications|4574,4585
:|4585,4586
<EOL>|4586,4587
1.|4587,4589
OxycoDONE|4590,4599
-|4599,4600
Acetaminophen|4600,4613
Elixir|4614,4620
_|4621,4622
_|4622,4623
_|4623,4624
mL|4625,4627
PO|4628,4630
Q4H|4631,4634
:|4634,4635
PRN|4635,4638
Pain|4639,4643
<EOL>|4644,4645
RX|4645,4647
*|4648,4649
oxycodone|4649,4658
-|4658,4659
acetaminophen|4659,4672
[|4673,4674
Roxicet|4674,4681
]|4681,4682
5|4683,4684
mg|4685,4687
-|4687,4688
325|4688,4691
mg|4692,4694
/|4694,4695
5|4695,4696
mL|4697,4699
_|4700,4701
_|4701,4702
_|4702,4703
ml|4704,4706
<EOL>|4707,4708
by|4708,4710
mouth|4711,4716
every|4717,4722
four|4723,4727
(|4728,4729
4|4729,4730
)|4730,4731
hours|4732,4737
Disp|4738,4742
#|4743,4744
*|4744,4745
250|4745,4748
Milliliter|4749,4759
Refills|4760,4767
:|4767,4768
*|4768,4769
0|4769,4770
<EOL>|4770,4771
2.|4771,4773
Docusate|4774,4782
Sodium|4783,4789
(|4790,4791
Liquid|4791,4797
)|4797,4798
100|4799,4802
mg|4803,4805
PO|4806,4808
BID|4809,4812
:|4812,4813
PRN|4813,4816
Constipation|4817,4829
<EOL>|4830,4831
RX|4831,4833
*|4834,4835
docusate|4835,4843
sodium|4844,4850
50|4851,4853
mg|4854,4856
/|4856,4857
5|4857,4858
mL|4859,4861
_|4862,4863
_|4863,4864
_|4864,4865
ml|4866,4868
by|4869,4871
mouth|4872,4877
twice|4878,4883
a|4884,4885
day|4886,4889
Disp|4890,4894
<EOL>|4895,4896
#|4896,4897
*|4897,4898
250|4898,4901
Milliliter|4902,4912
Refills|4913,4920
:|4920,4921
*|4921,4922
0|4922,4923
<EOL>|4923,4924
3.|4924,4926
Ascorbic|4927,4935
Acid|4936,4940
_|4941,4942
_|4942,4943
_|4943,4944
mg|4945,4947
PO|4948,4950
DAILY|4951,4956
<EOL>|4957,4958
4.|4958,4960
cholecalciferol|4961,4976
(|4977,4978
vitamin|4978,4985
D3|4986,4988
)|4988,4989
*|4990,4991
NF|4991,4993
*|4993,4994
3,000|4995,5000
unit|5001,5005
Oral|5006,5010
daily|5011,5016
<EOL>|5017,5018
5.|5018,5020
Multivitamins|5021,5034
W|5035,5036
/|5036,5037
minerals|5037,5045
1|5046,5047
TAB|5048,5051
PO|5052,5054
DAILY|5055,5060
<EOL>|5061,5062
<EOL>|5062,5063
<EOL>|5064,5065
Discharge|5065,5074
Disposition|5075,5086
:|5086,5087
<EOL>|5087,5088
Home|5088,5092
<EOL>|5092,5093
<EOL>|5094,5095
Discharge|5095,5104
Diagnosis|5105,5114
:|5114,5115
<EOL>|5115,5116
Morbid|5116,5122
obesity|5123,5130
<EOL>|5130,5131
Obstructive|5131,5142
sleep|5143,5148
apnea|5149,5154
<EOL>|5154,5155
<EOL>|5155,5156
<EOL>|5157,5158
Discharge|5158,5167
Condition|5168,5177
:|5177,5178
<EOL>|5178,5179
Mental|5179,5185
Status|5186,5192
:|5192,5193
Clear|5194,5199
and|5200,5203
coherent|5204,5212
.|5212,5213
<EOL>|5213,5214
Level|5214,5219
of|5220,5222
Consciousness|5223,5236
:|5236,5237
Alert|5238,5243
and|5244,5247
interactive|5248,5259
.|5259,5260
<EOL>|5260,5261
Activity|5261,5269
Status|5270,5276
:|5276,5277
Ambulatory|5278,5288
-|5289,5290
Independent|5291,5302
.|5302,5303
<EOL>|5303,5304
<EOL>|5304,5305
<EOL>|5306,5307
Discharge|5307,5316
Instructions|5317,5329
:|5329,5330
<EOL>|5330,5331
Discharge|5331,5340
Instructions|5341,5353
:|5353,5354
Please|5355,5361
call|5362,5366
your|5367,5371
surgeon|5372,5379
or|5380,5382
return|5383,5389
to|5390,5392
<EOL>|5393,5394
the|5394,5397
emergency|5398,5407
department|5408,5418
if|5419,5421
you|5422,5425
develop|5426,5433
a|5434,5435
fever|5436,5441
greater|5442,5449
than|5450,5454
<EOL>|5455,5456
101.5|5456,5461
,|5461,5462
chest|5463,5468
pain|5469,5473
,|5473,5474
shortness|5475,5484
of|5485,5487
breath|5488,5494
,|5494,5495
severe|5496,5502
abdominal|5503,5512
pain|5513,5517
,|5517,5518
<EOL>|5519,5520
pain|5520,5524
unrelieved|5525,5535
by|5536,5538
your|5539,5543
pain|5544,5548
medication|5549,5559
,|5559,5560
severe|5561,5567
nausea|5568,5574
or|5575,5577
<EOL>|5578,5579
vomiting|5579,5587
,|5587,5588
severe|5589,5595
abdominal|5596,5605
bloating|5606,5614
,|5614,5615
inability|5616,5625
to|5626,5628
eat|5629,5632
or|5633,5635
drink|5636,5641
,|5641,5642
<EOL>|5643,5644
foul|5644,5648
smelling|5649,5657
or|5658,5660
colorful|5661,5669
drainage|5670,5678
from|5679,5683
your|5684,5688
incisions|5689,5698
,|5698,5699
redness|5700,5707
<EOL>|5708,5709
or|5709,5711
swelling|5712,5720
around|5721,5727
your|5728,5732
incisions|5733,5742
,|5742,5743
or|5744,5746
any|5747,5750
other|5751,5756
symptoms|5757,5765
which|5766,5771
<EOL>|5772,5773
are|5773,5776
concerning|5777,5787
to|5788,5790
you|5791,5794
.|5794,5795
<EOL>|5795,5796
<EOL>|5796,5797
Diet|5797,5801
:|5801,5802
Stay|5803,5807
on|5808,5810
Stage|5811,5816
III|5817,5820
diet|5821,5825
until|5826,5831
your|5832,5836
follow|5837,5843
up|5844,5846
appointment|5847,5858
.|5858,5859
<EOL>|5860,5861
Do|5861,5863
not|5864,5867
self|5868,5872
advance|5873,5880
diet|5881,5885
,|5885,5886
do|5887,5889
not|5890,5893
drink|5894,5899
out|5900,5903
of|5904,5906
a|5907,5908
straw|5909,5914
or|5915,5917
chew|5918,5922
<EOL>|5923,5924
gum|5924,5927
.|5927,5928
<EOL>|5928,5929
<EOL>|5929,5930
Medication|5930,5940
Instructions|5941,5953
:|5953,5954
<EOL>|5954,5955
Resume|5955,5961
your|5962,5966
home|5967,5971
medications|5972,5983
except|5984,5990
please|5991,5997
do|5998,6000
not|6001,6004
take|6005,6009
your|6010,6014
<EOL>|6015,6016
cyclobenzaprine|6016,6031
while|6032,6037
taking|6038,6044
pain|6045,6049
medicaiton|6050,6060
.|6060,6061
<EOL>|6061,6062
<EOL>|6062,6063
CRUSH|6063,6068
ALL|6069,6072
PILLS|6073,6078
.|6078,6079
<EOL>|6079,6080
You|6080,6083
will|6084,6088
be|6089,6091
starting|6092,6100
some|6101,6105
new|6106,6109
medications|6110,6121
:|6121,6122
<EOL>|6122,6123
1|6123,6124
.|6124,6125
You|6127,6130
are|6131,6134
being|6135,6140
discharged|6141,6151
on|6152,6154
medications|6155,6166
to|6167,6169
treat|6170,6175
the|6176,6179
pain|6180,6184
<EOL>|6185,6186
from|6186,6190
your|6191,6195
operation|6196,6205
.|6205,6206
These|6207,6212
medications|6213,6224
will|6225,6229
make|6230,6234
you|6235,6238
drowsy|6239,6245
and|6246,6249
<EOL>|6250,6251
impair|6251,6257
your|6258,6262
ability|6263,6270
to|6271,6273
drive|6274,6279
a|6280,6281
motor|6282,6287
vehicle|6288,6295
or|6296,6298
operate|6299,6306
<EOL>|6307,6308
machinery|6308,6317
safely|6318,6324
.|6324,6325
You|6326,6329
MUST|6330,6334
refrain|6335,6342
from|6343,6347
such|6348,6352
activities|6353,6363
while|6364,6369
<EOL>|6370,6371
taking|6371,6377
these|6378,6383
medications|6384,6395
.|6395,6396
<EOL>|6396,6397
2|6397,6398
.|6398,6399
You|6400,6403
should|6404,6410
begin|6411,6416
taking|6417,6423
a|6424,6425
chewable|6426,6434
complete|6435,6443
multivitamin|6444,6456
with|6457,6461
<EOL>|6462,6463
minerals|6463,6471
.|6471,6472
No|6473,6475
gummy|6476,6481
vitamins|6482,6490
.|6490,6491
<EOL>|6491,6492
3|6492,6493
.|6493,6494
You|6495,6498
should|6499,6505
take|6506,6510
a|6511,6512
stool|6513,6518
softener|6519,6527
,|6527,6528
Colace|6529,6535
,|6535,6536
twice|6537,6542
daily|6543,6548
for|6549,6552
<EOL>|6553,6554
constipation|6554,6566
as|6567,6569
needed|6570,6576
,|6576,6577
or|6578,6580
until|6581,6586
you|6587,6590
resume|6591,6597
a|6598,6599
normal|6600,6606
bowel|6607,6612
<EOL>|6613,6614
pattern|6614,6621
.|6621,6622
<EOL>|6622,6623
4|6623,6624
.|6624,6625
You|6626,6629
must|6630,6634
not|6635,6638
use|6639,6642
NSAIDS|6643,6649
(|6650,6651
non-steroidal|6651,6664
anti-inflammatory|6665,6682
<EOL>|6683,6684
drugs|6684,6689
)|6689,6690
Examples|6691,6699
are|6700,6703
Ibuprofen|6704,6713
,|6713,6714
Motrin|6715,6721
,|6721,6722
Aleve|6723,6728
,|6728,6729
Nuprin|6730,6736
and|6737,6740
<EOL>|6741,6742
Naproxen|6742,6750
.|6750,6751
These|6752,6757
agents|6758,6764
will|6765,6769
cause|6770,6775
bleeding|6776,6784
and|6785,6788
ulcers|6789,6795
in|6796,6798
your|6799,6803
<EOL>|6804,6805
digestive|6805,6814
system|6815,6821
.|6821,6822
<EOL>|6822,6823
<EOL>|6823,6824
Activity|6824,6832
:|6832,6833
<EOL>|6833,6834
No|6834,6836
heavy|6837,6842
lifting|6843,6850
of|6851,6853
items|6854,6859
_|6860,6861
_|6861,6862
_|6862,6863
pounds|6864,6870
for|6871,6874
6|6875,6876
weeks|6877,6882
.|6882,6883
You|6884,6887
may|6888,6891
<EOL>|6892,6893
resume|6893,6899
moderate|6900,6908
exercise|6909,6917
at|6918,6920
your|6921,6925
discretion|6926,6936
,|6936,6937
no|6938,6940
abdominal|6941,6950
<EOL>|6951,6952
exercises|6952,6961
.|6961,6962
<EOL>|6962,6963
<EOL>|6963,6964
Wound|6964,6969
Care|6970,6974
:|6974,6975
<EOL>|6975,6976
You|6976,6979
may|6980,6983
shower|6984,6990
,|6990,6991
no|6992,6994
tub|6995,6998
baths|6999,7004
or|7005,7007
swimming|7008,7016
.|7016,7017
<EOL>|7018,7019
If|7019,7021
there|7022,7027
is|7028,7030
clear|7031,7036
drainage|7037,7045
from|7046,7050
your|7051,7055
incisions|7056,7065
,|7065,7066
cover|7067,7072
with|7073,7077
<EOL>|7078,7079
clean|7079,7084
,|7084,7085
dry|7086,7089
gauze|7090,7095
.|7095,7096
<EOL>|7097,7098
Your|7098,7102
steri|7103,7108
-|7108,7109
strips|7109,7115
will|7116,7120
fall|7121,7125
off|7126,7129
on|7130,7132
their|7133,7138
own|7139,7142
.|7142,7143
Please|7144,7150
remove|7151,7157
any|7158,7161
<EOL>|7162,7163
remaining|7163,7172
strips|7173,7179
_|7180,7181
_|7181,7182
_|7182,7183
days|7184,7188
after|7189,7194
surgery|7195,7202
.|7202,7203
<EOL>|7203,7204
Please|7204,7210
call|7211,7215
the|7216,7219
doctor|7220,7226
if|7227,7229
you|7230,7233
have|7234,7238
increased|7239,7248
pain|7249,7253
,|7253,7254
swelling|7255,7263
,|7263,7264
<EOL>|7265,7266
redness|7266,7273
,|7273,7274
or|7275,7277
drainage|7278,7286
from|7287,7291
the|7292,7295
incision|7296,7304
sites|7305,7310
.|7310,7311
<EOL>|7312,7313
<EOL>|7313,7314
<EOL>|7315,7316
Followup|7316,7324
Instructions|7325,7337
:|7337,7338
<EOL>|7338,7339
_|7339,7340
_|7340,7341
_|7341,7342
<EOL>|7342,7343

