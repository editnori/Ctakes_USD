 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
OBSTETRICS|152,162
/|162,163
GYNECOLOGY|163,173
<EOL>|173,174
<EOL>|175,176
Codeine|188,195
/|196,197
gabapentin|198,208
/|209,210
morphine|211,219
/|220,221
Amoxicillin|222,233
/|234,235
metronidazole|236,249
/|250,251
<EOL>|252,253
propoxyphene|253,265
/|266,267
rofecoxib|268,277
/|278,279
Macrobid|280,288
/|289,290
furosemide|291,301
/|302,303
Amitiza|304,311
/|312,313
<EOL>|314,315
Sulfa|315,320
(|321,322
Sulfonamide|322,333
Antibiotics|334,345
)|345,346
/|347,348
Tylenol|349,356
/|357,358
Hydromorphone|359,372
/|373,374
<EOL>|375,376
Toradol|376,383
<EOL>|383,384
<EOL>|385,386
Attending|386,395
:|395,396
_|397,398
_|398,399
_|399,400
<EOL>|400,401
<EOL>|402,403
For|420,423
admission|424,433
:|433,434
elective|435,443
gynecologic|444,455
surgery|456,463
for|464,467
urinary|468,475
<EOL>|476,477
retention|477,486
<EOL>|486,487
For|487,490
MICU|491,495
transfer|496,504
:|504,505
Anaphylaxis|506,517
<EOL>|517,518
<EOL>|519,520
Major|520,525
Surgical|526,534
or|535,537
Invasive|538,546
Procedure|547,556
:|556,557
<EOL>|557,558
Stage|558,563
2|564,565
interstim|566,575
w|576,577
/|577,578
posterior|579,588
colporrhaphy|589,601
for|602,605
rectocele|606,615
+|616,617
<EOL>|618,619
enterocele|619,629
_|630,631
_|631,632
_|632,633
<EOL>|633,634
<EOL>|635,636
History|664,671
of|672,674
Present|675,682
Illness|683,690
:|690,691
Ms.|693,696
_|697,698
_|698,699
_|699,700
is|701,703
a|704,705
_|706,707
_|707,708
_|708,709
w|710,711
/|711,712
Hx|713,715
<EOL>|716,717
of|717,719
cervical|720,728
CA|729,731
s|732,733
/|733,734
p|734,735
radical|736,743
hysterectomy|744,756
c|757,758
/|758,759
b|759,760
chronic|761,768
_|769,770
_|770,771
_|771,772
<EOL>|773,774
lymphedema|774,784
and|785,788
urinary|789,796
retention|797,806
,|806,807
for|808,811
which|812,817
she|818,821
frequently|822,832
<EOL>|833,834
self|834,838
-|838,839
caths|839,844
,|844,845
Asthma|846,852
,|852,853
GERD|854,858
,|858,859
IBS|860,863
,|863,864
anxiety|865,872
/|872,873
depression|873,883
,|883,884
fibromyalgia|885,897
<EOL>|898,899
and|899,902
other|903,908
issues|909,915
who|916,919
was|920,923
admitted|924,932
for|933,936
an|937,939
elective|940,948
gynecologic|949,960
<EOL>|961,962
surgery|962,969
(|970,971
stage|971,976
2|977,978
interstim|979,988
and|989,992
posterior|993,1002
colporrhaphy|1003,1015
w|1016,1017
/|1017,1018
graft|1019,1024
)|1024,1025
<EOL>|1026,1027
for|1027,1030
urinary|1031,1038
retention|1039,1048
and|1049,1052
rectocele|1053,1062
+|1063,1064
enterocele|1065,1075
.|1075,1076
<EOL>|1078,1079
<EOL>|1080,1081
Cervical|1103,1111
CA|1112,1114
s|1115,1116
/|1116,1117
p|1117,1118
radical|1119,1126
hysterectomy|1127,1139
c|1140,1141
/|1141,1142
b|1142,1143
chronic|1144,1151
_|1152,1153
_|1153,1154
_|1154,1155
lymphedema|1156,1166
<EOL>|1166,1167
ADHD|1167,1171
<EOL>|1171,1172
Anxiety|1172,1179
/|1179,1180
Depression|1180,1190
<EOL>|1190,1191
Asthma|1191,1197
<EOL>|1197,1198
Insomnia|1198,1206
<EOL>|1206,1207
GERD|1207,1211
<EOL>|1211,1212
Raynaud|1212,1219
's|1219,1221
<EOL>|1221,1222
IBS|1222,1225
<EOL>|1225,1226
Fibromyalgia|1226,1238
<EOL>|1240,1241
<EOL>|1241,1242
<EOL>|1243,1244
:|1258,1259
<EOL>|1259,1260
_|1260,1261
_|1261,1262
_|1262,1263
<EOL>|1263,1264
:|1278,1279
<EOL>|1279,1280
+|1280,1281
Hx|1281,1283
of|1284,1286
atopy|1287,1292
in|1293,1295
son|1296,1299
,|1299,1300
daughter|1301,1309
;|1309,1310
both|1311,1315
w|1316,1317
/|1317,1318
frequent|1319,1327
allergy|1328,1335
rxns|1336,1340
<EOL>|1341,1342
requiring|1342,1351
epi|1352,1355
pens|1356,1360
<EOL>|1360,1361
<EOL>|1362,1363
MICU|1378,1382
ADMISSION|1383,1392
EXAM|1393,1397
:|1397,1398
<EOL>|1398,1399
-|1399,1400
-|1400,1401
-|1401,1402
-|1402,1403
-|1403,1404
-|1404,1405
-|1405,1406
-|1406,1407
-|1407,1408
-|1408,1409
-|1409,1410
-|1410,1411
-|1411,1412
-|1412,1413
-|1413,1414
-|1414,1415
-|1415,1416
-|1416,1417
-|1417,1418
-|1418,1419
<EOL>|1419,1420
<EOL>|1420,1421
Vitals|1421,1427
:|1427,1428
T|1429,1430
:|1430,1431
98.7|1432,1436
BP|1437,1439
:|1439,1440
113|1441,1444
/|1444,1445
83|1445,1447
P|1448,1449
:|1449,1450
79|1451,1453
R|1454,1455
:|1455,1456
18|1457,1459
O2|1460,1462
:|1462,1463
97|1464,1466
%|1466,1467
_|1468,1469
_|1469,1470
_|1470,1471
<EOL>|1473,1474
_|1474,1475
_|1475,1476
_|1476,1477
:|1477,1478
Well|1479,1483
appearing|1484,1493
female|1494,1500
in|1501,1503
no|1504,1506
acute|1507,1512
distress|1513,1521
,|1521,1522
slightly|1523,1531
<EOL>|1532,1533
muffled|1533,1540
voice|1541,1546
,|1546,1547
somewhat|1548,1556
flushed|1557,1564
skin|1565,1569
<EOL>|1569,1570
HEENT|1570,1575
:|1575,1576
Moist|1577,1582
mucous|1583,1589
membranes|1590,1599
,|1599,1600
mild|1601,1605
lip|1606,1609
swelling|1610,1618
,|1618,1619
tongue|1620,1626
not|1627,1630
<EOL>|1631,1632
grossly|1632,1639
edematous|1640,1649
,|1649,1650
no|1651,1653
angioedema|1654,1664
<EOL>|1664,1665
Neck|1665,1669
:|1669,1670
JVP|1671,1674
non|1675,1678
elevated|1679,1687
<EOL>|1687,1688
CV|1688,1690
:|1690,1691
Regular|1692,1699
rate|1700,1704
and|1705,1708
rhythm|1709,1715
,|1715,1716
normal|1717,1723
S1|1724,1726
S2|1727,1729
,|1729,1730
no|1731,1733
murmurs|1734,1741
<EOL>|1741,1742
Lungs|1742,1747
:|1747,1748
Clear|1749,1754
to|1755,1757
auscultation|1758,1770
bilaterally|1771,1782
,|1782,1783
no|1784,1786
<EOL>|1787,1788
wheezes|1788,1795
/|1795,1796
rales|1796,1801
/|1801,1802
rhonchi|1802,1809
<EOL>|1809,1810
Abdomen|1810,1817
:|1817,1818
Soft|1819,1823
,|1823,1824
normoactive|1825,1836
bowel|1837,1842
sounds|1843,1849
,|1849,1850
nontender|1851,1860
,|1860,1861
<EOL>|1862,1863
nondistended|1863,1875
,|1875,1876
no|1877,1879
rebound|1880,1887
or|1888,1890
guarding|1891,1899
<EOL>|1899,1900
GU|1900,1902
:|1902,1903
Foley|1904,1909
in|1910,1912
place|1913,1918
<EOL>|1918,1919
Ext|1919,1922
:|1922,1923
Warm|1925,1929
,|1929,1930
trace|1931,1936
_|1937,1938
_|1938,1939
_|1939,1940
edema|1941,1946
,|1946,1947
peripheral|1948,1958
pulses|1959,1965
2|1966,1967
+|1967,1968
_|1969,1970
_|1970,1971
_|1971,1972
<EOL>|1972,1973
Neuro|1973,1978
:|1978,1979
alert|1980,1985
and|1986,1989
oriented|1990,1998
to|1999,2001
person|2002,2008
,|2008,2009
hospital|2010,2018
,|2018,2019
and|2020,2023
date|2024,2028
<EOL>|2028,2029
<EOL>|2029,2030
MICU|2030,2034
DISCHARGE|2035,2044
EXAM|2045,2049
:|2049,2050
<EOL>|2050,2051
-|2051,2052
-|2052,2053
-|2053,2054
-|2054,2055
-|2055,2056
-|2056,2057
-|2057,2058
-|2058,2059
-|2059,2060
-|2060,2061
-|2061,2062
-|2062,2063
-|2063,2064
-|2064,2065
-|2065,2066
-|2066,2067
-|2067,2068
-|2068,2069
-|2069,2070
-|2070,2071
<EOL>|2071,2072
<EOL>|2072,2073
Vitals|2073,2079
:|2079,2080
T|2081,2082
:|2082,2083
97.5|2084,2088
BP|2089,2091
:|2091,2092
107|2093,2096
/|2096,2097
62|2097,2099
P|2100,2101
:|2101,2102
84|2103,2105
R|2106,2107
:|2107,2108
16|2109,2111
O2|2112,2114
:|2114,2115
99|2116,2118
%|2118,2119
_|2120,2121
_|2121,2122
_|2122,2123
<EOL>|2125,2126
_|2126,2127
_|2127,2128
_|2128,2129
:|2129,2130
Well|2131,2135
appearing|2136,2145
female|2146,2152
in|2153,2155
no|2156,2158
acute|2159,2164
distress|2165,2173
,|2173,2174
normal|2175,2181
<EOL>|2182,2183
voice|2183,2188
,|2188,2189
somewhat|2190,2198
flushed|2199,2206
skin|2207,2211
,|2211,2212
most|2213,2217
prominent|2218,2227
in|2228,2230
malar|2231,2236
<EOL>|2237,2238
distribution|2238,2250
on|2251,2253
face|2254,2258
<EOL>|2258,2259
HEENT|2259,2264
:|2264,2265
Moist|2266,2271
mucous|2272,2278
membranes|2279,2288
,|2288,2289
appearance|2290,2300
of|2301,2303
face|2304,2308
unchanged|2309,2318
from|2319,2323
<EOL>|2324,2325
yesterday|2325,2334
,|2334,2335
tongue|2336,2342
not|2343,2346
edematous|2347,2356
,|2356,2357
no|2358,2360
angioedema|2361,2371
<EOL>|2371,2372
Neck|2372,2376
:|2376,2377
JVP|2378,2381
non|2382,2385
elevated|2386,2394
<EOL>|2394,2395
CV|2395,2397
:|2397,2398
Regular|2399,2406
rate|2407,2411
and|2412,2415
rhythm|2416,2422
,|2422,2423
normal|2424,2430
S1|2431,2433
S2|2434,2436
,|2436,2437
no|2438,2440
murmurs|2441,2448
<EOL>|2448,2449
Lungs|2449,2454
:|2454,2455
Clear|2456,2461
to|2462,2464
auscultation|2465,2477
bilaterally|2478,2489
,|2489,2490
no|2491,2493
<EOL>|2494,2495
wheezes|2495,2502
/|2502,2503
rales|2503,2508
/|2508,2509
rhonchi|2509,2516
<EOL>|2516,2517
Abdomen|2517,2524
:|2524,2525
Soft|2526,2530
,|2530,2531
normoactive|2532,2543
bowel|2544,2549
sounds|2550,2556
,|2556,2557
nontender|2558,2567
,|2567,2568
<EOL>|2569,2570
nondistended|2570,2582
,|2582,2583
no|2584,2586
rebound|2587,2594
or|2595,2597
guarding|2598,2606
<EOL>|2606,2607
GU|2607,2609
:|2609,2610
Foley|2611,2616
in|2617,2619
place|2620,2625
<EOL>|2625,2626
Ext|2626,2629
:|2629,2630
Warm|2632,2636
,|2636,2637
trace|2638,2643
_|2644,2645
_|2645,2646
_|2646,2647
edema|2648,2653
,|2653,2654
peripheral|2655,2665
pulses|2666,2672
2|2673,2674
+|2674,2675
_|2676,2677
_|2677,2678
_|2678,2679
<EOL>|2679,2680
Neuro|2680,2685
:|2685,2686
alert|2687,2692
and|2693,2696
oriented|2697,2705
to|2706,2708
person|2709,2715
,|2715,2716
hospital|2717,2725
,|2725,2726
and|2727,2730
date|2731,2735
<EOL>|2735,2736
<EOL>|2736,2737
GYN|2737,2740
Floor|2741,2746
discharge|2747,2756
exam|2757,2761
:|2761,2762
<EOL>|2762,2763
VSS|2763,2766
,|2766,2767
AF|2768,2770
<EOL>|2770,2771
Gen|2771,2774
:|2774,2775
NAD|2776,2779
A|2780,2781
&|2781,2782
O|2782,2783
x|2784,2785
3|2786,2787
<EOL>|2787,2788
Resp|2788,2792
:|2792,2793
no|2794,2796
visible|2797,2804
respiratory|2805,2816
distress|2817,2825
,|2825,2826
speaking|2827,2835
in|2836,2838
full|2839,2843
<EOL>|2844,2845
sentences|2845,2854
<EOL>|2854,2855
Abd|2855,2858
:|2858,2859
soft|2860,2864
,|2864,2865
NT|2866,2868
ND|2869,2871
<EOL>|2871,2872
Ext|2872,2875
:|2875,2876
moving|2877,2883
all|2884,2887
4|2888,2889
extremities|2890,2901
<EOL>|2901,2902
<EOL>|2902,2903
<EOL>|2904,2905
Pertinent|2905,2914
Results|2915,2922
:|2922,2923
<EOL>|2923,2924
MICU|2924,2928
ADMISSION|2929,2938
LABS|2939,2943
:|2943,2944
<EOL>|2944,2945
<EOL>|2945,2946
_|2946,2947
_|2947,2948
_|2948,2949
06|2950,2952
:|2952,2953
02PM|2953,2957
BLOOD|2958,2963
WBC|2964,2967
-|2967,2968
17|2968,2970
.|2970,2971
0|2971,2972
*|2972,2973
RBC|2974,2977
-|2977,2978
4|2978,2979
.|2979,2980
33|2980,2982
Hgb|2983,2986
-|2986,2987
13.9|2987,2991
Hct|2992,2995
-|2995,2996
39.1|2996,3000
<EOL>|3001,3002
MCV|3002,3005
-|3005,3006
90|3006,3008
MCH|3009,3012
-|3012,3013
32|3013,3015
.|3015,3016
2|3016,3017
*|3017,3018
MCHC|3019,3023
-|3023,3024
35|3024,3026
.|3026,3027
6|3027,3028
*|3028,3029
RDW|3030,3033
-|3033,3034
11.8|3034,3038
Plt|3039,3042
_|3043,3044
_|3044,3045
_|3045,3046
<EOL>|3046,3047
_|3047,3048
_|3048,3049
_|3049,3050
06|3051,3053
:|3053,3054
02PM|3054,3058
BLOOD|3059,3064
Neuts|3065,3070
-|3070,3071
94|3071,3073
.|3073,3074
5|3074,3075
*|3075,3076
Lymphs|3077,3083
-|3083,3084
4|3084,3085
.|3085,3086
3|3086,3087
*|3087,3088
Monos|3089,3094
-|3094,3095
0|3095,3096
.|3096,3097
7|3097,3098
*|3098,3099
<EOL>|3100,3101
Eos|3101,3104
-|3104,3105
0.1|3105,3108
Baso|3109,3113
-|3113,3114
0.3|3114,3117
<EOL>|3117,3118
_|3118,3119
_|3119,3120
_|3120,3121
06|3122,3124
:|3124,3125
02PM|3125,3129
BLOOD|3130,3135
_|3136,3137
_|3137,3138
_|3138,3139
PTT|3140,3143
-|3143,3144
31.8|3144,3148
_|3149,3150
_|3150,3151
_|3151,3152
<EOL>|3152,3153
_|3153,3154
_|3154,3155
_|3155,3156
06|3157,3159
:|3159,3160
02PM|3160,3164
BLOOD|3165,3170
Glucose|3171,3178
-|3178,3179
146|3179,3182
*|3182,3183
UreaN|3184,3189
-|3189,3190
16|3190,3192
Creat|3193,3198
-|3198,3199
0.8|3199,3202
Na|3203,3205
-|3205,3206
140|3206,3209
<EOL>|3210,3211
K|3211,3212
-|3212,3213
3.9|3213,3216
Cl|3217,3219
-|3219,3220
106|3220,3223
HCO3|3224,3228
-|3228,3229
24|3229,3231
AnGap|3232,3237
-|3237,3238
14|3238,3240
<EOL>|3240,3241
_|3241,3242
_|3242,3243
_|3243,3244
06|3245,3247
:|3247,3248
02PM|3248,3252
BLOOD|3253,3258
Calcium|3259,3266
-|3266,3267
9.1|3267,3270
Phos|3271,3275
-|3275,3276
3.1|3276,3279
Mg|3280,3282
-|3282,3283
1.5|3283,3286
*|3286,3287
<EOL>|3287,3288
_|3288,3289
_|3289,3290
_|3290,3291
06|3292,3294
:|3294,3295
02PM|3295,3299
BLOOD|3300,3305
TRYPTASE|3306,3314
-|3314,3315
PND|3315,3318
<EOL>|3318,3319
<EOL>|3319,3320
MICU|3320,3324
DISCHARGE|3325,3334
LABS|3335,3339
:|3339,3340
<EOL>|3340,3341
<EOL>|3341,3342
_|3342,3343
_|3343,3344
_|3344,3345
02|3346,3348
:|3348,3349
59AM|3349,3353
BLOOD|3354,3359
WBC|3360,3363
-|3363,3364
20|3364,3366
.|3366,3367
1|3367,3368
*|3368,3369
RBC|3370,3373
-|3373,3374
3|3374,3375
.|3375,3376
98|3376,3378
*|3378,3379
Hgb|3380,3383
-|3383,3384
12.6|3384,3388
Hct|3389,3392
-|3392,3393
36.3|3393,3397
<EOL>|3398,3399
MCV|3399,3402
-|3402,3403
91|3403,3405
MCH|3406,3409
-|3409,3410
31.6|3410,3414
MCHC|3415,3419
-|3419,3420
34.7|3420,3424
RDW|3425,3428
-|3428,3429
11.9|3429,3433
Plt|3434,3437
_|3438,3439
_|3439,3440
_|3440,3441
<EOL>|3441,3442
_|3442,3443
_|3443,3444
_|3444,3445
02|3446,3448
:|3448,3449
59AM|3449,3453
BLOOD|3454,3459
Plt|3460,3463
_|3464,3465
_|3465,3466
_|3466,3467
<EOL>|3467,3468
_|3468,3469
_|3469,3470
_|3470,3471
02|3472,3474
:|3474,3475
59AM|3475,3479
BLOOD|3480,3485
Glucose|3486,3493
-|3493,3494
152|3494,3497
*|3497,3498
UreaN|3499,3504
-|3504,3505
18|3505,3507
Creat|3508,3513
-|3513,3514
0.8|3514,3517
Na|3518,3520
-|3520,3521
138|3521,3524
<EOL>|3525,3526
K|3526,3527
-|3527,3528
3.5|3528,3531
Cl|3532,3534
-|3534,3535
102|3535,3538
HCO3|3539,3543
-|3543,3544
24|3544,3546
AnGap|3547,3552
-|3552,3553
16|3553,3555
<EOL>|3555,3556
_|3556,3557
_|3557,3558
_|3558,3559
02|3560,3562
:|3562,3563
59AM|3563,3567
BLOOD|3568,3573
Calcium|3574,3581
-|3581,3582
9.1|3582,3585
Phos|3586,3590
-|3590,3591
4.0|3591,3594
Mg|3595,3597
-|3597,3598
2|3598,3599
.|3599,3600
8|3600,3601
*|3601,3602
<EOL>|3602,3603
<EOL>|3603,3604
PERTINENT|3604,3613
LABS|3614,3618
:|3618,3619
<EOL>|3619,3620
<EOL>|3620,3621
_|3621,3622
_|3622,3623
_|3623,3624
06|3625,3627
:|3627,3628
02PM|3628,3632
BLOOD|3633,3638
WBC|3639,3642
-|3642,3643
17|3643,3645
.|3645,3646
0|3646,3647
*|3647,3648
RBC|3649,3652
-|3652,3653
4|3653,3654
.|3654,3655
33|3655,3657
Hgb|3658,3661
-|3661,3662
13.9|3662,3666
Hct|3667,3670
-|3670,3671
39.1|3671,3675
<EOL>|3676,3677
MCV|3677,3680
-|3680,3681
90|3681,3683
MCH|3684,3687
-|3687,3688
32|3688,3690
.|3690,3691
2|3691,3692
*|3692,3693
MCHC|3694,3698
-|3698,3699
35|3699,3701
.|3701,3702
6|3702,3703
*|3703,3704
RDW|3705,3708
-|3708,3709
11.8|3709,3713
Plt|3714,3717
_|3718,3719
_|3719,3720
_|3720,3721
<EOL>|3721,3722
_|3722,3723
_|3723,3724
_|3724,3725
06|3726,3728
:|3728,3729
02PM|3729,3733
BLOOD|3734,3739
Neuts|3740,3745
-|3745,3746
94|3746,3748
.|3748,3749
5|3749,3750
*|3750,3751
Lymphs|3752,3758
-|3758,3759
4|3759,3760
.|3760,3761
3|3761,3762
*|3762,3763
Monos|3764,3769
-|3769,3770
0|3770,3771
.|3771,3772
7|3772,3773
*|3773,3774
<EOL>|3775,3776
Eos|3776,3779
-|3779,3780
0.1|3780,3783
Baso|3784,3788
-|3788,3789
0.3|3789,3792
<EOL>|3792,3793
_|3793,3794
_|3794,3795
_|3795,3796
06|3797,3799
:|3799,3800
02PM|3800,3804
BLOOD|3805,3810
_|3811,3812
_|3812,3813
_|3813,3814
PTT|3815,3818
-|3818,3819
31.8|3819,3823
_|3824,3825
_|3825,3826
_|3826,3827
<EOL>|3827,3828
_|3828,3829
_|3829,3830
_|3830,3831
06|3832,3834
:|3834,3835
02PM|3835,3839
BLOOD|3840,3845
Glucose|3846,3853
-|3853,3854
146|3854,3857
*|3857,3858
UreaN|3859,3864
-|3864,3865
16|3865,3867
Creat|3868,3873
-|3873,3874
0.8|3874,3877
Na|3878,3880
-|3880,3881
140|3881,3884
<EOL>|3885,3886
K|3886,3887
-|3887,3888
3.9|3888,3891
Cl|3892,3894
-|3894,3895
106|3895,3898
HCO3|3899,3903
-|3903,3904
24|3904,3906
AnGap|3907,3912
-|3912,3913
14|3913,3915
<EOL>|3915,3916
_|3916,3917
_|3917,3918
_|3918,3919
06|3920,3922
:|3922,3923
02PM|3923,3927
BLOOD|3928,3933
Calcium|3934,3941
-|3941,3942
9.1|3942,3945
Phos|3946,3950
-|3950,3951
3.1|3951,3954
Mg|3955,3957
-|3957,3958
1.5|3958,3961
*|3961,3962
<EOL>|3962,3963
_|3963,3964
_|3964,3965
_|3965,3966
06|3967,3969
:|3969,3970
02PM|3970,3974
BLOOD|3975,3980
TRYPTASE|3981,3989
-|3989,3990
PND|3990,3993
<EOL>|3993,3994
<EOL>|3994,3995
PERTINENT|3995,4004
IMAGING|4005,4012
:|4012,4013
<EOL>|4013,4014
<EOL>|4014,4015
None|4015,4019
<EOL>|4019,4020
<EOL>|4020,4021
PERTINENT|4021,4030
MICRO|4031,4036
:|4036,4037
<EOL>|4037,4038
<EOL>|4038,4039
None|4039,4043
<EOL>|4043,4044
<EOL>|4045,4046
Ms.|4069,4072
_|4073,4074
_|4074,4075
_|4075,4076
is|4077,4079
a|4080,4081
_|4082,4083
_|4083,4084
_|4084,4085
y|4086,4087
/|4087,4088
o|4088,4089
F|4090,4091
w|4092,4093
/|4093,4094
Hx|4095,4097
of|4098,4100
cervical|4101,4109
CA|4110,4112
s|4113,4114
/|4114,4115
p|4115,4116
radical|4117,4124
<EOL>|4125,4126
hysterectomy|4126,4138
c|4139,4140
/|4140,4141
b|4141,4142
chronic|4143,4150
_|4151,4152
_|4152,4153
_|4153,4154
lymphedema|4155,4165
and|4166,4169
urinary|4170,4177
retention|4178,4187
,|4187,4188
<EOL>|4189,4190
Asthma|4190,4196
,|4196,4197
GERD|4198,4202
,|4202,4203
anxiety|4204,4211
/|4211,4212
depression|4212,4222
,|4222,4223
fibromyalgia|4224,4236
.|4236,4237
Please|4238,4244
refer|4245,4250
to|4251,4253
<EOL>|4254,4255
the|4255,4258
operative|4259,4268
report|4269,4275
for|4276,4279
full|4280,4284
details|4285,4292
.|4292,4293
<EOL>|4293,4294
<EOL>|4294,4295
Her|4295,4298
post-operative|4299,4313
course|4314,4320
was|4321,4324
uncomplicated|4325,4338
.|4338,4339
Immediately|4340,4351
<EOL>|4352,4353
post-op|4353,4360
,|4360,4361
her|4362,4365
pain|4366,4370
was|4371,4374
controlled|4375,4385
with|4386,4390
IV|4391,4393
dilaudid|4394,4402
and|4403,4406
toradol|4407,4414
.|4414,4415
<EOL>|4416,4417
However|4417,4424
,|4424,4425
in|4426,4428
the|4429,4432
PACU|4433,4437
,|4437,4438
the|4439,4442
patient|4443,4450
started|4451,4458
feeling|4459,4466
itchy|4467,4472
.|4472,4473
Once|4475,4479
<EOL>|4480,4481
the|4481,4484
pt|4485,4487
returned|4488,4496
to|4497,4499
the|4500,4503
floor|4504,4509
,|4509,4510
she|4511,4514
noted|4515,4520
sensation|4521,4530
of|4531,4533
tongue|4534,4540
/|4541,4542
<EOL>|4543,4544
lip|4544,4547
swelling|4548,4556
,|4556,4557
difficulty|4558,4568
swallowing|4569,4579
secretions|4580,4590
,|4590,4591
and|4592,4595
a|4596,4597
change|4598,4604
in|4605,4607
<EOL>|4608,4609
her|4609,4612
voice|4613,4618
.|4618,4619
No|4621,4623
SOB|4624,4627
,|4627,4628
no|4629,4631
flushing|4632,4640
,|4640,4641
no|4642,4644
stridor|4645,4652
or|4653,4655
wheeze|4656,4662
.|4662,4663
She|4665,4668
was|4669,4672
<EOL>|4673,4674
administered|4674,4686
an|4687,4689
Epi|4690,4693
-|4693,4694
pen|4694,4697
,|4697,4698
Solumedrol|4699,4709
100|4710,4713
mg|4714,4716
IV|4717,4719
,|4719,4720
Famotidine|4721,4731
20|4732,4734
mg|4735,4737
<EOL>|4738,4739
IV|4739,4741
,|4741,4742
and|4743,4746
Hydroxyzine|4747,4758
25|4759,4761
mg|4762,4764
IM|4765,4767
.|4767,4768
She|4770,4773
was|4774,4777
transferred|4778,4789
to|4790,4792
the|4793,4796
MICU|4797,4801
<EOL>|4802,4803
for|4803,4806
closer|4807,4813
monitoring|4814,4824
.|4824,4825
<EOL>|4826,4827
<EOL>|4827,4828
The|4828,4831
patient|4832,4839
has|4840,4843
numerous|4844,4852
drug|4853,4857
allergies|4858,4867
and|4868,4871
was|4872,4875
administered|4876,4888
the|4889,4892
<EOL>|4893,4894
following|4894,4903
medications|4904,4915
intra-operatively|4916,4933
:|4933,4934
Midazolam|4935,4944
,|4944,4945
Rocuronium|4946,4956
,|4956,4957
<EOL>|4958,4959
Fentanyl|4959,4967
,|4967,4968
Dexamethasone|4969,4982
,|4982,4983
Hydromorphone|4984,4997
,|4997,4998
Ondansetron|4999,5010
,|5010,5011
Lidocaine|5012,5021
,|5021,5022
<EOL>|5023,5024
Propofol|5024,5032
,|5032,5033
Cefazolin|5034,5043
,|5043,5044
Glycopyrrolate|5045,5059
,|5059,5060
Phenylephrine|5061,5074
,|5074,5075
and|5076,5079
<EOL>|5080,5081
Ketorolac|5081,5090
.|5090,5091
<EOL>|5091,5092
<EOL>|5092,5093
In|5093,5095
the|5096,5099
MICU|5100,5104
,|5104,5105
initial|5106,5113
VS|5114,5116
were|5117,5121
HR|5122,5124
87|5125,5127
,|5127,5128
BP|5129,5131
100|5132,5135
/|5135,5136
63|5136,5138
,|5138,5139
RR|5140,5142
17|5143,5145
,|5145,5146
S|5147,5148
100|5149,5152
%|5152,5153
<EOL>|5154,5155
_|5155,5156
_|5156,5157
_|5157,5158
.|5158,5159
The|5161,5164
patient|5165,5172
was|5173,5176
in|5177,5179
NAD|5180,5183
,|5183,5184
without|5185,5192
wheeze|5193,5199
or|5200,5202
poor|5203,5207
air|5208,5211
<EOL>|5212,5213
movement|5213,5221
on|5222,5224
exam|5225,5229
,|5229,5230
but|5231,5234
complained|5235,5245
of|5246,5248
persistent|5249,5259
voice|5260,5265
change|5266,5272
and|5273,5276
<EOL>|5277,5278
difficulty|5278,5288
swallowing|5289,5299
,|5299,5300
for|5301,5304
which|5305,5310
she|5311,5314
required|5315,5323
2|5324,5325
more|5326,5330
epi|5331,5334
pens|5335,5339
.|5339,5340
<EOL>|5342,5343
Has|5343,5346
remained|5347,5355
hemodynamically|5356,5371
stable|5372,5378
and|5379,5382
without|5383,5390
respiratory|5391,5402
<EOL>|5403,5404
compromise|5404,5414
.|5414,5415
<EOL>|5415,5416
<EOL>|5416,5417
ACTIVE|5417,5423
ISSUES|5424,5430
:|5430,5431
<EOL>|5431,5432
<EOL>|5432,5433
*|5433,5434
)|5434,5435
Post|5436,5440
operative|5441,5450
care|5451,5455
<EOL>|5455,5456
Her|5456,5459
pain|5460,5464
was|5465,5468
controlled|5469,5479
immediately|5480,5491
post-op|5492,5499
with|5500,5504
IV|5505,5507
dilaudid|5508,5516
and|5517,5520
<EOL>|5521,5522
toradol|5522,5529
.|5529,5530
This|5531,5535
was|5536,5539
transitioned|5540,5552
to|5553,5555
po|5556,5558
oxycodone|5559,5568
as|5569,5571
it|5572,5574
was|5575,5578
<EOL>|5579,5580
difficult|5580,5589
to|5590,5592
determine|5593,5602
what|5603,5607
was|5608,5611
causing|5612,5619
an|5620,5622
allergic|5623,5631
reaction|5632,5640
in|5641,5643
<EOL>|5644,5645
Ms.|5645,5648
_|5649,5650
_|5650,5651
_|5651,5652
.|5652,5653
<EOL>|5653,5654
<EOL>|5654,5655
Her|5655,5658
vaginal|5659,5666
packing|5667,5674
was|5675,5678
removed|5679,5686
on|5687,5689
POD|5690,5693
1|5694,5695
,|5695,5696
on|5697,5699
post-operative|5700,5714
day|5715,5718
<EOL>|5719,5720
2|5720,5721
,|5721,5722
her|5723,5726
urine|5727,5732
output|5733,5739
was|5740,5743
adequate|5744,5752
and|5753,5756
her|5757,5760
Foley|5761,5766
was|5767,5770
removed|5771,5778
.|5778,5779
The|5780,5783
<EOL>|5784,5785
patient|5785,5792
was|5793,5796
able|5797,5801
to|5802,5804
void|5805,5809
spontaneously|5810,5823
,|5823,5824
but|5825,5828
did|5829,5832
require|5833,5840
<EOL>|5841,5842
self|5842,5846
-|5846,5847
catheterization|5847,5862
_|5863,5864
_|5864,5865
_|5865,5866
times|5867,5872
a|5873,5874
day|5875,5878
based|5879,5884
on|5885,5887
a|5888,5889
sensation|5890,5899
of|5900,5902
<EOL>|5903,5904
bladder|5904,5911
fullness|5912,5920
.|5920,5921
<EOL>|5922,5923
<EOL>|5923,5924
*|5924,5925
)|5925,5926
Anaphylaxis|5927,5938
:|5938,5939
<EOL>|5940,5941
In|5941,5943
the|5944,5947
PACU|5948,5952
the|5953,5956
patient|5957,5964
awoke|5965,5970
and|5971,5974
started|5975,5982
feeling|5983,5990
pruritis|5991,5999
.|5999,6000
Once|6001,6005
<EOL>|6006,6007
she|6007,6010
arrived|6011,6018
to|6019,6021
the|6022,6025
floor|6026,6031
,|6031,6032
the|6033,6036
patient|6037,6044
noted|6045,6050
difficulty|6051,6061
talking|6062,6069
,|6069,6070
<EOL>|6071,6072
subjectively|6072,6084
swollen|6085,6092
lips|6093,6097
/|6097,6098
tongue|6098,6104
,|6104,6105
and|6106,6109
vocal|6110,6115
changes|6116,6123
.|6123,6124
No|6125,6127
SOB|6128,6131
,|6131,6132
no|6133,6135
<EOL>|6136,6137
flushing|6137,6145
,|6145,6146
no|6147,6149
stridor|6150,6157
or|6158,6160
wheeze|6161,6167
.|6167,6168
A|6169,6170
trigger|6171,6178
was|6179,6182
called|6183,6189
for|6190,6193
<EOL>|6194,6195
anaphyllaxis|6195,6207
and|6208,6211
she|6212,6215
recieved|6216,6224
an|6225,6227
Epi|6228,6231
-|6231,6232
pen|6232,6235
,|6235,6236
Solumedrol|6237,6247
100|6248,6251
mg|6252,6254
IV|6255,6257
,|6257,6258
<EOL>|6259,6260
Famotidine|6260,6270
20|6271,6273
mg|6274,6276
IV|6277,6279
,|6279,6280
and|6281,6284
Hydroxyzine|6285,6296
25|6297,6299
mg|6300,6302
IM|6303,6305
.|6305,6306
She|6308,6311
was|6312,6315
<EOL>|6316,6317
transferred|6317,6328
to|6329,6331
the|6332,6335
MICU|6336,6340
for|6341,6344
closer|6345,6351
monitoring|6352,6362
.|6362,6363
<EOL>|6364,6365
<EOL>|6365,6366
In|6366,6368
the|6369,6372
MICU|6373,6377
,|6377,6378
initial|6379,6386
VS|6387,6389
were|6390,6394
HR|6395,6397
87|6398,6400
,|6400,6401
BP|6402,6404
100|6405,6408
/|6408,6409
63|6409,6411
,|6411,6412
RR|6413,6415
17|6416,6418
,|6418,6419
S|6420,6421
100|6422,6425
%|6425,6426
<EOL>|6427,6428
_|6428,6429
_|6429,6430
_|6430,6431
.|6431,6432
The|6434,6437
patient|6438,6445
was|6446,6449
in|6450,6452
NAD|6453,6456
,|6456,6457
without|6458,6465
wheeze|6466,6472
or|6473,6475
poor|6476,6480
air|6481,6484
<EOL>|6485,6486
movement|6486,6494
on|6495,6497
exam|6498,6502
,|6502,6503
but|6504,6507
complained|6508,6518
of|6519,6521
persistent|6522,6532
voice|6533,6538
change|6539,6545
and|6546,6549
<EOL>|6550,6551
difficulty|6551,6561
swallowing|6562,6572
,|6572,6573
for|6574,6577
which|6578,6583
she|6584,6587
required|6588,6596
2|6597,6598
more|6599,6603
epi|6604,6607
pens|6608,6612
.|6612,6613
<EOL>|6615,6616
Has|6616,6619
remained|6620,6628
hemodynamically|6629,6644
stable|6645,6651
and|6652,6655
without|6656,6663
respiratory|6664,6675
<EOL>|6676,6677
compromise|6677,6687
.|6687,6688
<EOL>|6689,6690
<EOL>|6690,6691
Of|6691,6693
note|6694,6698
,|6698,6699
patient|6700,6707
was|6708,6711
lying|6712,6717
comfortable|6718,6729
in|6730,6732
bed|6733,6736
around|6737,6743
2200|6744,6748
and|6749,6752
<EOL>|6753,6754
continuing|6754,6764
to|6765,6767
inquire|6768,6775
about|6776,6781
more|6782,6786
Epi|6787,6790
-|6790,6791
pens|6791,6795
vs|6796,6798
epinephrine|6799,6810
gtt|6811,6814
<EOL>|6815,6816
despite|6816,6823
comfortable|6824,6835
respiration|6836,6847
,|6847,6848
vocalization|6849,6861
,|6861,6862
non-edematous|6863,6876
<EOL>|6877,6878
oral|6878,6882
structures|6883,6893
.|6893,6894
She|6895,6898
also|6899,6903
perseverated|6904,6916
about|6917,6922
her|6923,6926
Ativan|6927,6933
and|6934,6937
<EOL>|6938,6939
Ambien|6939,6945
,|6945,6946
as|6947,6949
well|6950,6954
as|6955,6957
her|6958,6961
propranolol|6962,6973
for|6974,6977
essential|6978,6987
tremor|6988,6994
despite|6995,7002
<EOL>|7003,7004
explanation|7004,7015
that|7016,7020
beta|7021,7025
blockers|7026,7034
can|7035,7038
worsen|7039,7045
bronchoconstriction|7046,7065
<EOL>|7066,7067
and|7067,7070
respiratory|7071,7082
compromise|7083,7093
in|7094,7096
anaphylaxis|7097,7108
.|7108,7109
<EOL>|7109,7110
<EOL>|7110,7111
On|7111,7113
the|7114,7117
day|7118,7121
she|7122,7125
was|7126,7129
called|7130,7136
out|7137,7140
to|7141,7143
the|7144,7147
floor|7148,7153
,|7153,7154
the|7155,7158
pt|7159,7161
complained|7162,7172
of|7173,7175
<EOL>|7176,7177
persistent|7177,7187
facial|7188,7194
flushing|7195,7203
.|7203,7204
She|7206,7209
was|7210,7213
afebrile|7214,7222
,|7222,7223
hemodynamically|7224,7239
<EOL>|7240,7241
stable|7241,7247
,|7247,7248
and|7249,7252
without|7253,7260
respiratory|7261,7272
compromise|7273,7283
or|7284,7286
systemic|7287,7295
symptoms|7296,7304
.|7304,7305
<EOL>|7306,7307
Symptomatic|7308,7319
care|7320,7324
with|7325,7329
hydroxyzine|7330,7341
and|7342,7345
eucerin|7346,7353
lotion|7354,7360
was|7361,7364
<EOL>|7365,7366
provided|7366,7374
.|7374,7375
<EOL>|7375,7376
<EOL>|7376,7377
Upon|7377,7381
step|7382,7386
down|7387,7391
to|7392,7394
the|7395,7398
floor|7399,7404
,|7404,7405
the|7406,7409
patient|7410,7417
again|7418,7423
reported|7424,7432
to|7433,7435
<EOL>|7436,7437
nursing|7437,7444
that|7445,7449
she|7450,7453
felt|7454,7458
throat|7459,7465
constriction|7466,7478
.|7478,7479
Epinephrine|7480,7491
and|7492,7495
<EOL>|7496,7497
solumedrol|7497,7507
were|7508,7512
given|7513,7518
and|7519,7522
the|7523,7526
patient|7527,7534
felt|7535,7539
relief|7540,7546
.|7546,7547
Allergy|7548,7555
was|7556,7559
<EOL>|7560,7561
consulted|7561,7570
,|7570,7571
and|7572,7575
they|7576,7580
asked|7581,7586
us|7587,7589
to|7590,7592
stop|7593,7597
all|7598,7601
new|7602,7605
medications|7606,7617
given|7618,7623
<EOL>|7624,7625
to|7625,7627
her|7628,7631
while|7632,7637
at|7638,7640
the|7641,7644
hospital|7645,7653
,|7653,7654
and|7655,7658
to|7659,7661
report|7662,7668
all|7669,7672
of|7673,7675
them|7676,7680
as|7681,7683
<EOL>|7684,7685
allergies|7685,7694
.|7694,7695
In|7696,7698
addition|7699,7707
,|7707,7708
we|7709,7711
sent|7712,7716
out|7717,7720
a|7721,7722
tryptase|7723,7731
level|7732,7737
,|7737,7738
as|7739,7741
well|7742,7746
as|7747,7749
<EOL>|7750,7751
coordinated|7751,7762
outpatient|7763,7773
follow|7774,7780
-|7780,7781
up|7781,7783
with|7784,7788
them|7789,7793
.|7793,7794
<EOL>|7795,7796
<EOL>|7796,7797
#|7797,7798
Chronic|7798,7805
_|7806,7807
_|7807,7808
_|7808,7809
edema|7810,7815
:|7815,7816
Continue|7817,7825
home|7826,7830
Metolazone|7831,7841
,|7841,7842
spironolactone|7843,7857
,|7857,7858
<EOL>|7859,7860
potassium|7860,7869
repletion|7870,7879
as|7880,7882
not|7883,7886
hypotensive|7887,7898
.|7898,7899
We|7901,7903
monitored|7904,7913
her|7914,7917
K|7918,7919
<EOL>|7920,7921
during|7921,7927
her|7928,7931
stay|7932,7936
,|7936,7937
which|7938,7943
was|7944,7947
WNL|7948,7951
.|7951,7952
<EOL>|7952,7953
<EOL>|7953,7954
#|7954,7955
Asthma|7955,7961
:|7961,7962
Home|7963,7967
Albuterol|7968,7977
use|7978,7981
_|7982,7983
_|7983,7984
_|7984,7985
per|7986,7989
week|7990,7994
,|7994,7995
did|7996,7999
not|8000,8003
require|8004,8011
in|8012,8014
<EOL>|8015,8016
the|8016,8019
MICU|8020,8024
.|8024,8025
<EOL>|8026,8027
<EOL>|8027,8028
#|8028,8029
GERD|8029,8033
:|8033,8034
Nexium|8035,8041
(|8042,8043
was|8043,8046
initially|8047,8056
held|8057,8061
on|8062,8064
admission|8065,8074
,|8074,8075
but|8076,8079
per|8080,8083
pt|8084,8086
<EOL>|8087,8088
request|8088,8095
was|8096,8099
given|8100,8105
on|8106,8108
_|8109,8110
_|8110,8111
_|8111,8112
prior|8113,8118
to|8119,8121
advancing|8122,8131
diet|8132,8136
)|8136,8137
<EOL>|8137,8138
<EOL>|8138,8139
#|8139,8140
ADHD|8140,8144
:|8144,8145
On|8146,8148
Adderall|8149,8157
,|8157,8158
held|8159,8163
on|8164,8166
admission|8167,8176
<EOL>|8176,8177
<EOL>|8177,8178
#|8178,8179
Anxiety|8180,8187
/|8187,8188
depression|8188,8198
/|8198,8199
fibromyalgia|8199,8211
:|8211,8212
lorazepam|8213,8222
<EOL>|8223,8224
<EOL>|8224,8225
#|8225,8226
Insomnia|8227,8235
:|8235,8236
zolpidem|8237,8245
<EOL>|8245,8246
<EOL>|8246,8247
By|8247,8249
post-operative|8250,8264
day|8265,8268
1|8269,8270
,|8270,8271
she|8272,8275
was|8276,8279
tolerating|8280,8290
a|8291,8292
regular|8293,8300
diet|8301,8305
,|8305,8306
<EOL>|8307,8308
ambulating|8308,8318
independently|8319,8332
,|8332,8333
and|8334,8337
pain|8338,8342
was|8343,8346
controlled|8347,8357
with|8358,8362
oral|8363,8367
<EOL>|8368,8369
medications|8369,8380
.|8380,8381
She|8382,8385
was|8386,8389
the|8390,8393
discharged|8395,8405
home|8406,8410
in|8411,8413
stable|8414,8420
condition|8421,8430
<EOL>|8431,8432
with|8432,8436
outpatient|8437,8447
follow|8448,8454
-|8454,8455
up|8455,8457
scheduled|8458,8467
.|8467,8468
She|8469,8472
was|8473,8476
also|8477,8481
scheduled|8482,8491
to|8492,8494
<EOL>|8495,8496
have|8496,8500
an|8501,8503
appointment|8504,8515
with|8516,8520
Allergy|8521,8528
and|8529,8532
Immunology|8533,8543
.|8543,8544
<EOL>|8544,8545
<EOL>|8545,8546
<EOL>|8547,8548
Medications|8548,8559
on|8560,8562
Admission|8563,8572
:|8572,8573
<EOL>|8573,8574
Albuterol|8574,8583
sulfate|8584,8591
2.5|8592,8595
mg|8596,8598
/|8598,8599
3|8599,8600
mL|8601,8603
(|8604,8605
0.083|8605,8610
%|8611,8612
)|8612,8613
Neb|8614,8617
TID|8618,8621
PRN|8622,8625
<EOL>|8625,8626
Albuterol|8626,8635
ProAir|8636,8642
HFA|8643,8646
90|8647,8649
mcg|8650,8653
INH|8654,8657
1|8658,8659
puff|8660,8664
BID|8665,8668
PRN|8669,8672
<EOL>|8673,8674
Cephalexin|8674,8684
250|8685,8688
mg|8689,8691
Q6H|8692,8695
<EOL>|8695,8696
Adderall|8696,8704
XR|8705,8707
15|8708,8710
mg|8711,8713
BID|8714,8717
<EOL>|8717,8718
Ergocalciferol|8718,8732
(|8733,8734
vitamin|8734,8741
D2|8742,8744
)|8744,8745
50,000|8746,8752
U|8753,8754
Q|8755,8756
week|8757,8761
<EOL>|8761,8762
Nexium|8762,8768
40|8769,8771
mg|8772,8774
_|8775,8776
_|8776,8777
_|8777,8778
QAM|8779,8782
<EOL>|8782,8783
Vivelle|8783,8790
0.075|8791,8796
mg|8797,8799
/|8799,8800
24|8800,8802
hr|8803,8805
Transderm|8806,8815
Patch|8816,8821
2x|8822,8824
/|8825,8826
week|8827,8831
<EOL>|8832,8833
Diflucan|8833,8841
200|8842,8845
mg|8846,8848
Q|8849,8850
_|8851,8852
_|8852,8853
_|8853,8854
<EOL>|8855,8856
Hydroxyzine|8856,8867
HCl|8868,8871
25|8872,8874
mg|8875,8877
QD|8878,8880
PRN|8881,8884
<EOL>|8885,8886
Ibuprofen|8886,8895
600|8896,8899
mg|8900,8902
Q8H|8903,8906
PRN|8907,8910
<EOL>|8910,8911
Linzess|8911,8918
(|8919,8920
linactolide|8920,8931
)|8931,8932
145|8933,8936
mcg|8937,8940
QD|8941,8943
<EOL>|8943,8944
Ativan|8944,8950
1|8951,8952
mg|8953,8955
QD|8956,8958
PRN|8959,8962
<EOL>|8963,8964
Metolazone|8964,8974
2.5|8975,8978
mg|8979,8981
QD|8982,8984
<EOL>|8984,8985
Zofran|8985,8991
8|8992,8993
mg|8994,8996
PO|8997,8999
PRN|9000,9003
<EOL>|9004,9005
Oxycodone|9005,9014
5|9015,9016
mg|9017,9019
PO|9020,9022
Q6H|9023,9026
PRN|9027,9030
<EOL>|9031,9032
Potassium|9032,9041
chloride|9042,9050
10|9051,9053
%|9054,9055
Oral|9056,9060
Liquid|9061,9067
30ml|9068,9072
PO|9073,9075
QID|9076,9079
<EOL>|9079,9080
Propranolol|9080,9091
ER|9092,9094
80|9095,9097
mg|9098,9100
ER|9101,9103
QHS|9104,9107
<EOL>|9107,9108
Spironolactone|9108,9122
100|9123,9126
mg|9127,9129
QD|9130,9132
<EOL>|9132,9133
Trimethoprim|9133,9145
100|9146,9149
mg|9150,9152
tablet|9153,9159
QD|9160,9162
<EOL>|9162,9163
Ambien|9163,9169
10|9170,9172
mg|9173,9175
QHS|9176,9179
<EOL>|9179,9180
#|9180,9181
14|9181,9183
_|9184,9185
_|9185,9186
_|9186,9187
catheter|9188,9196
<EOL>|9197,9198
Docusate|9198,9206
sodium|9207,9213
100|9214,9217
mg|9218,9220
BID|9221,9224
<EOL>|9224,9225
LACTOBACILLUS|9225,9238
COMBINATION|9239,9250
<EOL>|9250,9251
<EOL>|9252,9253
Discharge|9253,9262
Medications|9263,9274
:|9274,9275
<EOL>|9275,9276
1.|9276,9278
Docusate|9279,9287
Sodium|9288,9294
(|9295,9296
Liquid|9296,9302
)|9302,9303
100|9304,9307
mg|9308,9310
PO|9311,9313
BID|9314,9317
<EOL>|9318,9319
RX|9319,9321
*|9322,9323
docusate|9323,9331
sodium|9332,9338
100|9339,9342
mg|9343,9345
1|9346,9347
tablet|9348,9354
by|9355,9357
mouth|9358,9363
twice|9364,9369
a|9370,9371
day|9372,9375
Disp|9376,9380
<EOL>|9381,9382
#|9382,9383
*|9383,9384
60|9384,9386
Capsule|9387,9394
Refills|9395,9402
:|9402,9403
*|9403,9404
0|9404,9405
<EOL>|9405,9406
2.|9406,9408
Bisacodyl|9409,9418
10|9419,9421
mg|9422,9424
PO|9425,9427
/|9427,9428
PR|9428,9430
DAILY|9431,9436
:|9436,9437
PRN|9437,9440
Constipation|9441,9453
<EOL>|9454,9455
RX|9455,9457
*|9458,9459
bisacodyl|9459,9468
5|9469,9470
mg|9471,9473
_|9474,9475
_|9475,9476
_|9476,9477
tablet|9478,9484
,|9484,9485
delayed|9485,9492
release|9493,9500
(|9501,9502
_|9502,9503
_|9503,9504
_|9504,9505
)|9505,9506
by|9507,9509
<EOL>|9510,9511
mouth|9511,9516
constipation|9517,9529
Disp|9530,9534
#|9535,9536
*|9536,9537
20|9537,9539
Tablet|9540,9546
Refills|9547,9554
:|9554,9555
*|9555,9556
0|9556,9557
<EOL>|9557,9558
3.|9558,9560
Metolazone|9561,9571
2.5|9572,9575
mg|9576,9578
PO|9579,9581
DAILY|9582,9587
<EOL>|9588,9589
4.|9589,9591
NexIUM|9592,9598
(|9599,9600
esomeprazole|9600,9612
magnesium|9613,9622
)|9622,9623
40|9624,9626
mg|9627,9629
Oral|9630,9634
once|9635,9639
Duration|9640,9648
:|9648,9649
1|9650,9651
<EOL>|9652,9653
Dose|9653,9657
<EOL>|9658,9659
5.|9659,9661
OxycoDONE|9662,9671
(|9672,9673
Immediate|9673,9682
Release|9683,9690
)|9690,9691
_|9693,9694
_|9694,9695
_|9695,9696
mg|9697,9699
PO|9700,9702
Q6H|9703,9706
:|9706,9707
PRN|9707,9710
pain|9711,9715
<EOL>|9716,9717
do|9717,9719
not|9720,9723
drive|9724,9729
and|9730,9733
drink|9734,9739
on|9740,9742
this|9743,9747
medication|9748,9758
<EOL>|9759,9760
RX|9760,9762
*|9763,9764
oxycodone|9764,9773
5|9774,9775
mg|9776,9778
_|9779,9780
_|9780,9781
_|9781,9782
tablet|9783,9789
(|9789,9790
s|9790,9791
)|9791,9792
by|9793,9795
mouth|9796,9801
every|9802,9807
6|9808,9809
hrs|9810,9813
Disp|9814,9818
#|9819,9820
*|9820,9821
20|9821,9823
<EOL>|9824,9825
Tablet|9825,9831
Refills|9832,9839
:|9839,9840
*|9840,9841
0|9841,9842
<EOL>|9842,9843
6.|9843,9845
Propranolol|9846,9857
LA|9858,9860
80|9861,9863
mg|9864,9866
PO|9867,9869
DAILY|9870,9875
<EOL>|9876,9877
7.|9877,9879
Spironolactone|9880,9894
100|9895,9898
mg|9899,9901
PO|9902,9904
DAILY|9905,9910
<EOL>|9911,9912
8.|9912,9914
Zolpidem|9915,9923
Tartrate|9924,9932
5|9933,9934
mg|9935,9937
PO|9938,9940
HS|9941,9943
<EOL>|9944,9945
9.|9945,9947
Trimethoprim|9948,9960
100|9961,9964
mg|9965,9967
PO|9968,9970
DAILY|9971,9976
<EOL>|9977,9978
10.|9978,9981
Vivelle|9982,9989
(|9990,9991
estradiol|9991,10000
)|10000,10001
0.075|10002,10007
mg|10008,10010
/|10010,10011
24|10011,10013
hr|10014,10016
Transdermal|10017,10028
twice|10029,10034
/|10034,10035
week|10035,10039
<EOL>|10040,10041
11|10041,10043
.|10043,10044
Lorazepam|10045,10054
1|10055,10056
mg|10057,10059
PO|10060,10062
DAILY|10063,10068
:|10068,10069
PRN|10069,10072
anxiety|10073,10080
<EOL>|10081,10082
12.|10082,10085
Potassium|10086,10095
Chloride|10096,10104
40|10105,10107
mEq|10108,10111
PO|10112,10114
DAILY|10115,10120
Duration|10121,10129
:|10129,10130
24|10131,10133
Hours|10134,10139
<EOL>|10140,10141
Hold|10141,10145
for|10146,10149
K|10150,10151
>|10152,10153
<EOL>|10154,10155
<EOL>|10155,10156
<EOL>|10157,10158
Discharge|10158,10167
Disposition|10168,10179
:|10179,10180
<EOL>|10180,10181
Home|10181,10185
<EOL>|10185,10186
<EOL>|10187,10188
Discharge|10188,10197
Diagnosis|10198,10207
:|10207,10208
<EOL>|10208,10209
urinary|10209,10216
retention|10217,10226
,|10226,10227
rectocele|10228,10237
<EOL>|10237,10238
<EOL>|10238,10239
<EOL>|10240,10241
Mental|10262,10268
Status|10269,10275
:|10275,10276
Clear|10277,10282
and|10283,10286
coherent|10287,10295
.|10295,10296
<EOL>|10296,10297
Level|10297,10302
of|10303,10305
Consciousness|10306,10319
:|10319,10320
Alert|10321,10326
and|10327,10330
interactive|10331,10342
.|10342,10343
<EOL>|10343,10344
Activity|10344,10352
Status|10353,10359
:|10359,10360
Ambulatory|10361,10371
-|10372,10373
Independent|10374,10385
.|10385,10386
<EOL>|10386,10387
<EOL>|10387,10388
<EOL>|10389,10390
Dear|10414,10418
_|10419,10420
_|10420,10421
_|10421,10422
,|10422,10423
<EOL>|10423,10424
<EOL>|10424,10425
You|10425,10428
were|10429,10433
admitted|10434,10442
to|10443,10445
the|10446,10449
Gynecology|10450,10460
service|10461,10468
after|10469,10474
your|10475,10479
scheduled|10480,10489
<EOL>|10490,10491
Stage|10491,10496
2|10497,10498
Insterstim|10499,10509
placement|10510,10519
and|10520,10523
posterior|10524,10533
colporrhaphy|10534,10546
with|10547,10551
<EOL>|10552,10553
graft|10553,10558
for|10559,10562
urinary|10563,10570
retention|10571,10580
and|10581,10584
rectocele|10585,10594
and|10595,10598
enterocele|10599,10609
.|10609,10610
You|10612,10615
<EOL>|10616,10617
tolerated|10617,10626
the|10627,10630
procedure|10631,10640
well|10641,10645
.|10645,10646
However|10647,10654
,|10654,10655
after|10656,10661
your|10662,10666
operation|10667,10676
,|10676,10677
you|10678,10681
<EOL>|10682,10683
had|10683,10686
a|10687,10688
severe|10689,10695
allergic|10696,10704
reaction|10705,10713
,|10713,10714
and|10715,10718
had|10719,10722
to|10723,10725
go|10726,10728
to|10729,10731
the|10732,10735
ICU|10736,10739
for|10740,10743
<EOL>|10744,10745
monitoring|10745,10755
.|10755,10756
Since|10757,10762
then|10763,10767
,|10767,10768
you|10769,10772
have|10773,10777
recovered|10778,10787
well|10788,10792
,|10792,10793
and|10794,10797
we|10798,10800
have|10801,10805
<EOL>|10806,10807
determined|10807,10817
that|10818,10822
you|10823,10826
are|10827,10830
in|10831,10833
stable|10834,10840
condition|10841,10850
for|10851,10854
discharge|10855,10864
.|10864,10865
<EOL>|10866,10867
Please|10867,10873
take|10874,10878
your|10879,10883
medication|10884,10894
and|10895,10898
follow|10899,10905
-|10905,10906
up|10906,10908
at|10909,10911
your|10912,10916
appointments|10917,10929
<EOL>|10930,10931
as|10931,10933
scheduled|10934,10943
.|10943,10944
<EOL>|10944,10945
<EOL>|10945,10946
_|10946,10947
_|10947,10948
_|10948,10949
instructions|10950,10962
:|10962,10963
<EOL>|10965,10966
*|10966,10967
Take|10968,10972
your|10973,10977
medications|10978,10989
as|10990,10992
prescribed|10993,11003
.|11003,11004
<EOL>|11006,11007
*|11007,11008
Do|11009,11011
not|11012,11015
drive|11016,11021
while|11022,11027
taking|11028,11034
narcotics|11035,11044
.|11044,11045
<EOL>|11046,11047
*|11047,11048
Take|11049,11053
a|11054,11055
stool|11056,11061
softener|11062,11070
such|11071,11075
as|11076,11078
colace|11079,11085
while|11086,11091
taking|11092,11098
narcotics|11099,11108
to|11109,11111
<EOL>|11112,11113
prevent|11113,11120
constipation|11121,11133
<EOL>|11134,11135
*|11135,11136
Do|11137,11139
not|11140,11143
combine|11144,11151
narcotic|11152,11160
and|11161,11164
sedative|11165,11173
medications|11174,11185
or|11186,11188
alcohol|11189,11196
<EOL>|11198,11199
*|11199,11200
Do|11201,11203
not|11204,11207
take|11208,11212
more|11213,11217
than|11218,11222
4000mg|11223,11229
acetaminophen|11230,11243
(|11244,11245
APAP|11245,11249
)|11249,11250
in|11251,11253
24|11254,11256
hrs|11257,11260
<EOL>|11262,11263
*|11263,11264
No|11265,11267
strenuous|11268,11277
activity|11278,11286
until|11287,11292
your|11293,11297
post-op|11298,11305
appointment|11306,11317
<EOL>|11319,11320
*|11320,11321
Nothing|11322,11329
in|11330,11332
the|11333,11336
vagina|11337,11343
(|11344,11345
no|11345,11347
tampons|11348,11355
,|11355,11356
no|11357,11359
douching|11360,11368
,|11368,11369
no|11370,11372
sex|11373,11376
)|11376,11377
for|11378,11381
6|11382,11383
<EOL>|11384,11385
weeks|11385,11390
<EOL>|11390,11391
*|11391,11392
No|11393,11395
heavy|11396,11401
lifting|11402,11409
of|11410,11412
objects|11413,11420
>|11421,11422
10lbs|11422,11427
for|11428,11431
6|11432,11433
weeks|11434,11439
.|11439,11440
<EOL>|11444,11445
*|11445,11446
You|11447,11450
may|11451,11454
eat|11455,11458
a|11459,11460
regular|11461,11468
diet|11469,11473
<EOL>|11475,11476
*|11476,11477
or|11478,11480
anything|11481,11489
that|11490,11494
concerns|11495,11503
you|11504,11507
<EOL>|11507,11508
<EOL>|11508,11509
Incision|11509,11517
care|11518,11522
:|11522,11523
<EOL>|11525,11526
*|11526,11527
You|11528,11531
may|11532,11535
shower|11536,11542
and|11543,11546
allow|11547,11552
soapy|11553,11558
water|11559,11564
to|11565,11567
run|11568,11571
over|11572,11576
incision|11577,11585
;|11585,11586
no|11587,11589
<EOL>|11590,11591
scrubbing|11591,11600
of|11601,11603
incision|11604,11612
.|11612,11613
No|11614,11616
bath|11617,11621
tubs|11622,11626
for|11627,11630
6|11631,11632
weeks|11633,11638
.|11638,11639
<EOL>|11641,11642
<EOL>|11643,11644
Call|11644,11648
your|11649,11653
doctor|11654,11660
for|11661,11664
:|11664,11665
<EOL>|11667,11668
*|11668,11669
fever|11670,11675
>|11676,11677
100.4|11678,11683
<EOL>|11685,11686
*|11686,11687
severe|11688,11694
abdominal|11695,11704
pain|11705,11709
<EOL>|11711,11712
*|11712,11713
difficulty|11714,11724
urinating|11725,11734
<EOL>|11736,11737
*|11737,11738
vaginal|11739,11746
bleeding|11747,11755
requiring|11756,11765
>|11766,11767
1|11767,11768
pad|11769,11772
/|11772,11773
hr|11773,11775
<EOL>|11777,11778
*|11778,11779
abnormal|11780,11788
vaginal|11789,11796
discharge|11797,11806
<EOL>|11808,11809
*|11809,11810
redness|11811,11818
or|11819,11821
drainage|11822,11830
from|11831,11835
incision|11836,11844
<EOL>|11846,11847
*|11847,11848
nausea|11849,11855
/|11855,11856
vomiting|11856,11864
where|11865,11870
you|11871,11874
are|11875,11878
unable|11879,11885
to|11886,11888
keep|11889,11893
down|11894,11898
fluids|11899,11905
/|11905,11906
food|11906,11910
<EOL>|11911,11912
or|11912,11914
your|11915,11919
medication|11920,11930
<EOL>|11932,11933
*|11933,11934
or|11935,11937
anything|11938,11946
that|11947,11951
concerns|11952,11960
you|11961,11964
<EOL>|11964,11965
<EOL>|11965,11966
To|11966,11968
reach|11969,11974
medical|11975,11982
records|11983,11990
to|11991,11993
get|11994,11997
the|11998,12001
records|12002,12009
from|12010,12014
this|12015,12019
<EOL>|12020,12021
hospitalization|12021,12036
sent|12037,12041
to|12042,12044
your|12045,12049
doctor|12050,12056
at|12057,12059
home|12060,12064
,|12064,12065
call|12066,12070
_|12071,12072
_|12072,12073
_|12073,12074
.|12074,12075
<EOL>|12076,12077
<EOL>|12077,12078
<EOL>|12079,12080
Followup|12080,12088
Instructions|12089,12101
:|12101,12102
<EOL>|12102,12103
_|12103,12104
_|12104,12105
_|12105,12106
<EOL>|12106,12107

