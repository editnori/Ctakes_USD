 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|22,26
No|27,29
:|29,30
_|33,34
_|34,35
_|35,36
<EOL>|36,37
<EOL>|38,39
Admission|39,48
Date|49,53
:|53,54
_|56,57
_|57,58
_|58,59
Discharge|73,82
Date|83,87
:|87,88
_|91,92
_|92,93
_|93,94
<EOL>|94,95
<EOL>|96,97
Date|97,101
of|102,104
Birth|105,110
:|110,111
_|113,114
_|114,115
_|115,116
Sex|129,132
:|132,133
F|136,137
<EOL>|137,138
<EOL>|139,140
Service|140,147
:|147,148
MEDICINE|149,157
<EOL>|157,158
<EOL>|159,160
Allergies|160,169
:|169,170
<EOL>|171,172
No|172,174
Known|175,180
Allergies|181,190
/|191,192
Adverse|193,200
Drug|201,205
Reactions|206,215
<EOL>|215,216
<EOL>|217,218
Attending|218,227
:|227,228
_|229,230
_|230,231
_|231,232
.|232,233
<EOL>|233,234
<EOL>|235,236
Chief|236,241
Complaint|242,251
:|251,252
<EOL>|252,253
fatigue|253,260
,|260,261
anemia|262,268
<EOL>|268,269
<EOL>|270,271
Major|271,276
Surgical|277,285
or|286,288
Invasive|289,297
Procedure|298,307
:|307,308
<EOL>|308,309
None|309,313
<EOL>|313,314
<EOL>|314,315
<EOL>|316,317
History|317,324
of|325,327
Present|328,335
Illness|336,343
:|343,344
<EOL>|344,345
Ms.|345,348
_|349,350
_|350,351
_|351,352
is|353,355
a|356,357
_|358,359
_|359,360
_|360,361
year|362,366
old|367,370
woman|371,376
with|377,381
a|382,383
past|384,388
medical|389,396
<EOL>|397,398
history|398,405
of|406,408
type|409,413
-|413,414
2|414,415
DM|416,418
,|418,419
hypertension|420,432
,|432,433
stage|434,439
IV|440,442
CKD|443,446
,|446,447
CAD|448,451
s|452,453
/|453,454
p|454,455
<EOL>|456,457
distant|457,464
MI|465,467
and|468,471
bare|472,476
metal|477,482
stent|483,488
,|488,489
stroke|490,496
,|496,497
recent|498,504
unprovoked|505,515
DVTs|516,520
<EOL>|521,522
on|522,524
Coumadin|525,533
,|533,534
and|535,538
recent|539,545
upper|546,551
GI|552,554
bleeding|555,563
,|563,564
who|565,568
was|569,572
sent|573,577
to|578,580
_|581,582
_|582,583
_|583,584
<EOL>|585,586
by|586,588
her|589,592
physician|593,602
for|603,606
anemia|607,613
(|614,615
Hgb|615,618
6.5|619,622
)|622,623
.|623,624
<EOL>|624,625
<EOL>|625,626
The|626,629
patient|630,637
was|638,641
admitted|642,650
to|651,653
_|654,655
_|655,656
_|656,657
in|658,660
_|661,662
_|662,663
_|663,664
with|665,669
unprovoked|670,680
<EOL>|681,682
bilateral|682,691
lower|692,697
extremity|698,707
DVTs|708,712
.|712,713
She|714,717
was|718,721
started|722,729
on|730,732
heparin|733,740
as|741,743
an|744,746
<EOL>|747,748
inpatient|748,757
,|757,758
but|759,762
anticoagulation|763,778
was|779,782
complicated|783,794
by|795,797
severely|798,806
<EOL>|807,808
elevated|808,816
PTT|817,820
(|821,822
>|822,823
150|823,826
)|826,827
and|828,831
upper|832,837
GI|838,840
bleed|841,846
.|846,847
Endoscopy|848,857
was|858,861
notable|862,869
<EOL>|870,871
for|871,874
significant|875,886
erythema|887,895
,|895,896
superficial|897,908
ulceration|909,919
,|919,920
and|921,924
gastritis|925,934
<EOL>|935,936
without|936,943
active|944,950
bleeding|951,959
.|959,960
She|961,964
was|965,968
placed|969,975
on|976,978
BID|979,982
PPI|983,986
prophylaxis|987,998
.|998,999
<EOL>|1000,1001
She|1001,1004
was|1005,1008
eventually|1009,1019
bridged|1020,1027
to|1028,1030
Coumadin|1031,1039
for|1040,1043
a|1044,1045
planned|1046,1053
6|1054,1055
month|1056,1061
<EOL>|1062,1063
course|1063,1069
.|1069,1070
Her|1071,1074
INR|1075,1078
is|1079,1081
managed|1082,1089
by|1090,1092
her|1093,1096
rehab|1097,1102
facility|1103,1111
,|1111,1112
and|1113,1116
she|1117,1120
is|1121,1123
<EOL>|1124,1125
followed|1125,1133
by|1134,1136
Dr.|1137,1140
_|1141,1142
_|1142,1143
_|1143,1144
in|1145,1147
_|1148,1149
_|1149,1150
_|1150,1151
clinic|1152,1158
.|1158,1159
<EOL>|1160,1161
<EOL>|1161,1162
For|1162,1165
the|1166,1169
last|1170,1174
two|1175,1178
weeks|1179,1184
she|1185,1188
has|1189,1192
noted|1193,1198
increasing|1199,1209
fatigue|1210,1217
along|1218,1223
<EOL>|1224,1225
with|1225,1229
shortness|1230,1239
of|1240,1242
breath|1243,1249
,|1249,1250
exertional|1251,1261
sub-sternal|1262,1273
chest|1274,1279
pain|1280,1284
<EOL>|1285,1286
relieved|1286,1294
with|1295,1299
rest|1300,1304
,|1304,1305
and|1306,1309
symmetrical|1310,1321
lower|1322,1327
extremity|1328,1337
swelling|1338,1346
.|1346,1347
<EOL>|1348,1349
During|1349,1355
this|1356,1360
period|1361,1367
she|1368,1371
reports|1372,1379
that|1380,1384
her|1385,1388
appetite|1389,1397
remained|1398,1406
good|1407,1411
,|1411,1412
<EOL>|1413,1414
and|1414,1417
he|1418,1420
bowel|1421,1426
function|1427,1435
was|1436,1439
normal|1440,1446
.|1446,1447
She|1448,1451
denies|1452,1458
bloody|1459,1465
stools|1466,1472
or|1473,1475
<EOL>|1476,1477
dark|1477,1481
stool|1482,1487
.|1487,1488
On|1489,1491
_|1492,1493
_|1493,1494
_|1494,1495
she|1496,1499
presented|1500,1509
to|1510,1512
her|1513,1516
PCP|1517,1520
office|1521,1527
from|1528,1532
rehab|1533,1538
<EOL>|1539,1540
reporting|1540,1549
increasing|1550,1560
shortness|1561,1570
of|1571,1573
breath|1574,1580
and|1581,1584
fatigue|1585,1592
.|1592,1593
She|1594,1597
was|1598,1601
<EOL>|1602,1603
found|1603,1608
to|1609,1611
have|1612,1616
a|1617,1618
Hgb|1619,1622
of|1623,1625
6.5|1626,1629
,|1629,1630
with|1631,1635
an|1636,1638
unconcerning|1639,1651
CXR|1652,1655
.|1655,1656
She|1657,1660
was|1661,1664
<EOL>|1665,1666
sent|1666,1670
to|1671,1673
the|1674,1677
_|1678,1679
_|1679,1680
_|1680,1681
ED|1682,1684
.|1684,1685
<EOL>|1685,1686
<EOL>|1686,1687
In|1687,1689
the|1690,1693
ED|1694,1696
,|1696,1697
her|1698,1701
initial|1702,1709
vitals|1710,1716
were|1717,1721
T|1722,1723
:|1723,1724
97.5|1725,1729
P|1730,1731
:|1731,1732
60|1733,1735
BP|1736,1738
:|1738,1739
156|1740,1743
/|1743,1744
76|1744,1746
RR|1747,1749
:|1749,1750
<EOL>|1751,1752
16|1752,1754
SPO2|1755,1759
:|1759,1760
100|1761,1764
%|1764,1765
RA.|1766,1769
Exam|1770,1774
was|1775,1778
notable|1779,1786
for|1787,1790
guiac|1791,1796
negative|1797,1805
stool|1806,1811
.|1811,1812
<EOL>|1813,1814
Imaging|1814,1821
was|1822,1825
notable|1826,1833
for|1834,1837
:|1837,1838
<EOL>|1838,1839
"|1840,1841
1|1841,1842
.|1842,1843
Nonocclusive|1844,1856
deep|1857,1861
vein|1862,1866
thrombosis|1867,1877
of|1878,1880
one|1881,1884
of|1885,1887
the|1888,1891
paired|1892,1898
<EOL>|1899,1900
posterior|1900,1909
tibial|1910,1916
veins|1917,1922
bilaterally|1923,1934
.|1934,1935
The|1936,1939
extent|1940,1946
of|1947,1949
thrombus|1950,1958
<EOL>|1959,1960
bilaterally|1960,1971
has|1972,1975
decreased|1976,1985
.|1985,1986
No|1987,1989
new|1990,1993
deep|1994,1998
venous|1999,2005
thrombosis|2006,2016
in|2017,2019
<EOL>|2020,2021
either|2021,2027
lower|2028,2033
extremity|2034,2043
.|2043,2044
<EOL>|2045,2046
2.|2047,2049
Right|2050,2055
complex|2056,2063
_|2064,2065
_|2065,2066
_|2066,2067
cyst|2068,2072
.|2072,2073
"|2073,2074
<EOL>|2074,2075
<EOL>|2075,2076
The|2076,2079
patient|2080,2087
was|2088,2091
transfused|2092,2102
with|2103,2107
2|2108,2109
units|2110,2115
of|2116,2118
pRBCs|2119,2124
,|2124,2125
with|2126,2130
<EOL>|2131,2132
appropriate|2132,2143
increase|2144,2152
in|2153,2155
Hgb|2156,2159
to|2160,2162
9.0|2163,2166
.|2166,2167
Following|2168,2177
transfusion|2178,2189
,|2189,2190
a|2191,2192
<EOL>|2193,2194
repeat|2194,2200
CXR|2201,2204
was|2205,2208
notable|2209,2216
for|2217,2220
pulmonary|2221,2230
edema|2231,2236
with|2237,2241
bilateral|2242,2251
<EOL>|2252,2253
pleural|2253,2260
effusions|2261,2270
.|2270,2271
She|2272,2275
was|2276,2279
given|2280,2285
20mg|2286,2290
PO|2291,2293
Lasix|2294,2299
and|2300,2303
40mg|2304,2308
IV|2309,2311
Lasix|2312,2317
<EOL>|2318,2319
in|2319,2321
the|2322,2325
ED|2326,2328
.|2328,2329
The|2330,2333
decision|2334,2342
was|2343,2346
made|2347,2351
to|2352,2354
admit|2355,2360
the|2361,2364
patient|2365,2372
for|2373,2376
anemia|2377,2383
<EOL>|2384,2385
and|2385,2388
flash|2389,2394
pulmonary|2395,2404
edema|2405,2410
.|2410,2411
<EOL>|2412,2413
<EOL>|2413,2414
On|2414,2416
the|2417,2420
floor|2421,2426
,|2426,2427
vitals|2428,2434
notable|2435,2442
for|2443,2446
T|2447,2448
:|2448,2449
97.9|2450,2454
BP|2455,2457
:|2457,2458
154|2459,2462
/|2462,2463
75|2463,2465
P|2466,2467
:|2467,2468
65|2469,2471
R|2472,2473
:|2473,2474
20|2475,2477
<EOL>|2478,2479
O2|2479,2481
:|2481,2482
99RA|2483,2487
FSBG|2488,2492
:|2492,2493
76|2494,2496
.|2496,2497
She|2498,2501
reports|2502,2509
no|2510,2512
acute|2513,2518
complaints|2519,2529
,|2529,2530
and|2531,2534
that|2535,2539
her|2540,2543
<EOL>|2544,2545
shortness|2545,2554
of|2555,2557
breath|2558,2564
has|2565,2568
resolved|2569,2577
.|2577,2578
She|2579,2582
denies|2583,2589
chest|2590,2595
pain|2596,2600
,|2600,2601
<EOL>|2602,2603
dizziness|2603,2612
,|2612,2613
lightheadedness|2614,2629
.|2629,2630
<EOL>|2630,2631
<EOL>|2632,2633
Past|2633,2637
Medical|2638,2645
History|2646,2653
:|2653,2654
<EOL>|2654,2655
-|2655,2656
hypertension|2657,2669
<EOL>|2671,2672
-|2672,2673
diabetes|2674,2682
<EOL>|2684,2685
-|2685,2686
hx|2687,2689
CVA|2690,2693
(|2694,2695
cerebellar|2695,2705
-|2705,2706
medullary|2706,2715
stroke|2716,2722
in|2723,2725
_|2726,2727
_|2727,2728
_|2728,2729
<EOL>|2731,2732
-|2732,2733
CAD|2734,2737
(|2738,2739
hx|2739,2741
of|2742,2744
MI|2745,2747
in|2748,2750
_|2751,2752
_|2752,2753
_|2753,2754
BMS|2755,2758
to|2759,2761
circumflex|2762,2772
and|2773,2776
POBA|2777,2781
_|2782,2783
_|2783,2784
_|2784,2785
<EOL>|2787,2788
-|2788,2789
peripheral|2790,2800
arterial|2801,2809
disease|2810,2817
-|2817,2818
claudication|2819,2831
,|2831,2832
followed|2833,2841
by|2842,2844
<EOL>|2845,2846
vascular|2846,2854
,|2854,2855
managed|2856,2863
conservatively|2864,2878
<EOL>|2878,2879
-|2879,2880
stage|2881,2886
IV|2887,2889
CKD|2890,2893
(|2894,2895
baseline|2895,2903
2.1|2904,2907
-|2907,2908
2.6|2908,2911
)|2911,2912
<EOL>|2914,2915
-|2915,2916
GERD|2917,2921
/|2921,2922
esophageal|2922,2932
rings|2933,2938
<EOL>|2938,2939
<EOL>|2940,2941
Social|2941,2947
History|2948,2955
:|2955,2956
<EOL>|2956,2957
_|2957,2958
_|2958,2959
_|2959,2960
<EOL>|2960,2961
Family|2961,2967
History|2968,2975
:|2975,2976
<EOL>|2976,2977
Niece|2977,2982
had|2983,2986
some|2987,2991
sort|2992,2996
of|2997,2999
cancer|3000,3006
.|3006,3007
Father|3008,3014
died|3015,3019
in|3020,3022
his|3023,3026
_|3027,3028
_|3028,3029
_|3029,3030
due|3031,3034
to|3035,3037
<EOL>|3038,3039
lung|3039,3043
disease|3044,3051
.|3051,3052
Mother|3054,3060
died|3061,3065
in|3066,3068
her|3069,3072
_|3073,3074
_|3074,3075
_|3075,3076
due|3077,3080
to|3081,3083
an|3084,3086
unknown|3087,3094
cause|3095,3100
.|3100,3101
<EOL>|3103,3104
No|3104,3106
early|3107,3112
CAD|3113,3116
or|3117,3119
sudden|3120,3126
cardiac|3127,3134
death|3135,3140
.|3140,3141
No|3142,3144
other|3145,3150
known|3151,3156
history|3157,3164
of|3165,3167
<EOL>|3168,3169
cancer|3169,3175
.|3175,3176
<EOL>|3176,3177
<EOL>|3178,3179
Physical|3179,3187
Exam|3188,3192
:|3192,3193
<EOL>|3193,3194
ADMISSION|3194,3203
PHYSICAL|3204,3212
EXAM|3213,3217
:|3217,3218
<EOL>|3220,3221
Vitals|3221,3227
:|3227,3228
T|3229,3230
:|3230,3231
97.9|3232,3236
BP|3237,3239
:|3239,3240
154|3241,3244
/|3244,3245
75|3245,3247
P|3248,3249
:|3249,3250
65|3251,3253
R|3254,3255
:|3255,3256
20|3257,3259
O2|3260,3262
:|3262,3263
99RA|3264,3268
FSBG|3269,3273
:|3273,3274
_|3275,3276
_|3276,3277
_|3277,3278
<EOL>|3279,3280
General|3280,3287
:|3287,3288
Overweight|3289,3299
woman|3300,3305
,|3305,3306
alert|3307,3312
,|3312,3313
oriented|3314,3322
,|3322,3323
no|3324,3326
acute|3327,3332
distress|3333,3341
<EOL>|3343,3344
HEENT|3344,3349
:|3349,3350
Sclera|3351,3357
anicteric|3358,3367
,|3367,3368
MMM|3369,3372
,|3372,3373
oropharynx|3374,3384
clear|3385,3390
<EOL>|3392,3393
Neck|3393,3397
:|3397,3398
supple|3399,3405
,|3405,3406
JVP|3407,3410
not|3411,3414
elevated|3415,3423
<EOL>|3425,3426
Lungs|3426,3431
:|3431,3432
Crackles|3433,3441
to|3442,3444
the|3445,3448
mid-lungs|3449,3458
bilaterally|3459,3470
<EOL>|3472,3473
CV|3473,3475
:|3475,3476
Regular|3477,3484
rate|3485,3489
and|3490,3493
rhythm|3494,3500
,|3500,3501
normal|3502,3508
S1|3509,3511
+|3512,3513
S2|3514,3516
,|3516,3517
no|3518,3520
murmurs|3521,3528
or|3529,3531
<EOL>|3532,3533
gallops|3533,3540
<EOL>|3542,3543
Abdomen|3543,3550
:|3550,3551
soft|3552,3556
,|3556,3557
non-tender|3558,3568
,|3568,3569
non-distended|3570,3583
,|3583,3584
bowel|3585,3590
sounds|3591,3597
present|3598,3605
,|3605,3606
<EOL>|3607,3608
no|3608,3610
rebound|3611,3618
tenderness|3619,3629
or|3630,3632
guarding|3633,3641
,|3641,3642
no|3643,3645
organomegaly|3646,3658
<EOL>|3660,3661
Ext|3661,3664
:|3664,3665
Warm|3666,3670
,|3670,3671
well|3672,3676
perfused|3677,3685
,|3685,3686
2|3687,3688
+|3688,3689
pulses|3690,3696
,|3696,3697
no|3698,3700
clubbing|3701,3709
or|3710,3712
cyanosis|3713,3721
.|3721,3722
2|3723,3724
+|3724,3725
<EOL>|3726,3727
pitting|3727,3734
edema|3735,3740
in|3741,3743
dependent|3744,3753
areas|3754,3759
to|3760,3762
the|3763,3766
buttocks|3767,3775
<EOL>|3777,3778
Skin|3778,3782
:|3782,3783
no|3784,3786
rashes|3787,3793
noted|3794,3799
<EOL>|3799,3800
Neuro|3800,3805
:|3805,3806
_|3807,3808
_|3808,3809
_|3809,3810
strength|3811,3819
in|3820,3822
deltoids|3823,3831
,|3831,3832
biceps|3833,3839
,|3839,3840
triceps|3841,3848
,|3848,3849
wrist|3850,3855
<EOL>|3856,3857
extensors|3857,3866
,|3866,3867
finger|3868,3874
extensors|3875,3884
,|3884,3885
hip|3886,3889
flexors|3890,3897
,|3897,3898
hamstrings|3899,3909
,|3909,3910
<EOL>|3911,3912
quadriceps|3912,3922
,|3922,3923
gastrocs|3924,3932
,|3932,3933
tibialis|3934,3942
anterior|3943,3951
,|3951,3952
bilaterally|3953,3964
.|3964,3965
Sensation|3966,3975
<EOL>|3976,3977
intact|3977,3983
bilaterally|3984,3995
.|3995,3996
<EOL>|3997,3998
PSYCH|3998,4003
:|4003,4004
Alert|4005,4010
and|4011,4014
fully|4015,4020
oriented|4021,4029
;|4029,4030
normal|4031,4037
mood|4038,4042
and|4043,4046
affect|4047,4053
.|4053,4054
<EOL>|4054,4055
sometimes|4055,4064
slow|4065,4069
to|4070,4072
respond|4073,4080
and|4081,4084
responding|4085,4095
with|4096,4100
repetitive|4101,4111
answers|4112,4119
<EOL>|4119,4120
but|4120,4123
otherwise|4124,4133
appropriate|4134,4145
<EOL>|4145,4146
<EOL>|4146,4147
DISCHARGE|4147,4156
PHYSICAL|4157,4165
EXAM|4166,4170
:|4170,4171
<EOL>|4171,4172
VS|4172,4174
:|4174,4175
T|4176,4177
:|4177,4178
97.6|4179,4183
BP|4184,4186
:|4186,4187
150s|4188,4192
-|4192,4193
160s|4193,4197
/|4197,4198
70s|4198,4201
-|4201,4202
80s|4202,4205
P|4206,4207
:|4207,4208
60s|4209,4212
-|4212,4213
70s|4213,4216
RR|4217,4219
:|4219,4220
18|4221,4223
SPO2|4224,4228
:|4228,4229
100RA|4230,4235
<EOL>|4235,4236
General|4236,4243
:|4243,4244
Overweight|4245,4255
woman|4256,4261
,|4261,4262
alert|4263,4268
,|4268,4269
oriented|4270,4278
,|4278,4279
no|4280,4282
acute|4283,4288
distress|4289,4297
<EOL>|4299,4300
HEENT|4300,4305
:|4305,4306
Sclera|4307,4313
anicteric|4314,4323
,|4323,4324
MMM|4325,4328
,|4328,4329
oropharynx|4330,4340
clear|4341,4346
<EOL>|4348,4349
Neck|4349,4353
:|4353,4354
supple|4355,4361
,|4361,4362
JVP|4363,4366
not|4367,4370
elevated|4371,4379
<EOL>|4381,4382
Lungs|4382,4387
:|4387,4388
Clear|4389,4394
to|4395,4397
auscultation|4398,4410
bilaterally|4411,4422
<EOL>|4422,4423
CV|4423,4425
:|4425,4426
Regular|4427,4434
rate|4435,4439
and|4440,4443
rhythm|4444,4450
,|4450,4451
normal|4452,4458
S1|4459,4461
+|4462,4463
S2|4464,4466
,|4466,4467
no|4468,4470
murmurs|4471,4478
or|4479,4481
<EOL>|4482,4483
gallops|4483,4490
<EOL>|4492,4493
Abdomen|4493,4500
:|4500,4501
soft|4502,4506
,|4506,4507
non-tender|4508,4518
,|4518,4519
non-distended|4520,4533
,|4533,4534
bowel|4535,4540
sounds|4541,4547
present|4548,4555
,|4555,4556
<EOL>|4557,4558
no|4558,4560
rebound|4561,4568
tenderness|4569,4579
or|4580,4582
guarding|4583,4591
,|4591,4592
no|4593,4595
organomegaly|4596,4608
<EOL>|4610,4611
Ext|4611,4614
:|4614,4615
Warm|4616,4620
,|4620,4621
well|4622,4626
perfused|4627,4635
,|4635,4636
2|4637,4638
+|4638,4639
pulses|4640,4646
,|4646,4647
no|4648,4650
clubbing|4651,4659
or|4660,4662
cyanosis|4663,4671
.|4671,4672
1|4673,4674
+|4674,4675
<EOL>|4676,4677
pitting|4677,4684
edema|4685,4690
in|4691,4693
shins|4694,4699
bilaterally|4700,4711
<EOL>|4711,4712
Skin|4712,4716
:|4716,4717
no|4718,4720
rashes|4721,4727
noted|4728,4733
<EOL>|4733,4734
<EOL>|4734,4735
<EOL>|4736,4737
Pertinent|4737,4746
Results|4747,4754
:|4754,4755
<EOL>|4755,4756
LABORATORY|4756,4766
STUDIES|4767,4774
ON|4775,4777
ADMISSION|4778,4787
<EOL>|4787,4788
=|4788,4789
=|4789,4790
=|4790,4791
=|4791,4792
=|4792,4793
=|4793,4794
=|4794,4795
=|4795,4796
=|4796,4797
=|4797,4798
=|4798,4799
=|4799,4800
=|4800,4801
=|4801,4802
=|4802,4803
=|4803,4804
=|4804,4805
=|4805,4806
=|4806,4807
=|4807,4808
=|4808,4809
=|4809,4810
=|4810,4811
=|4811,4812
=|4812,4813
=|4813,4814
=|4814,4815
=|4815,4816
=|4816,4817
=|4817,4818
=|4818,4819
=|4819,4820
=|4820,4821
=|4821,4822
=|4822,4823
=|4823,4824
=|4824,4825
=|4825,4826
=|4826,4827
=|4827,4828
=|4828,4829
=|4829,4830
=|4830,4831
=|4831,4832
=|4832,4833
<EOL>|4833,4834
_|4834,4835
_|4835,4836
_|4836,4837
12|4838,4840
:|4840,4841
30PM|4841,4845
WBC|4848,4851
-|4851,4852
4.4|4852,4855
RBC|4856,4859
-|4859,4860
2|4860,4861
.|4861,4862
03|4862,4864
*|4864,4865
HGB|4866,4869
-|4869,4870
6|4870,4871
.|4871,4872
5|4872,4873
*|4873,4874
HCT|4875,4878
-|4878,4879
20|4879,4881
.|4881,4882
6|4882,4883
*|4883,4884
<EOL>|4885,4886
MCV|4886,4889
-|4889,4890
102|4890,4893
*|4893,4894
#|4894,4895
MCH|4896,4899
-|4899,4900
32.0|4900,4904
MCHC|4905,4909
-|4909,4910
31|4910,4912
.|4912,4913
6|4913,4914
*|4914,4915
RDW|4916,4919
-|4919,4920
16|4920,4922
.|4922,4923
3|4923,4924
*|4924,4925
RDWSD|4926,4931
-|4931,4932
59|4932,4934
.|4934,4935
6|4935,4936
*|4936,4937
<EOL>|4937,4938
_|4938,4939
_|4939,4940
_|4940,4941
12|4942,4944
:|4944,4945
30PM|4945,4949
_|4952,4953
_|4953,4954
_|4954,4955
<EOL>|4955,4956
_|4956,4957
_|4957,4958
_|4958,4959
12|4960,4962
:|4962,4963
30PM|4963,4967
ALBUMIN|4970,4977
-|4977,4978
4.1|4978,4981
CALCIUM|4982,4989
-|4989,4990
9.2|4990,4993
PHOSPHATE|4994,5003
-|5003,5004
4|5004,5005
.|5005,5006
7|5006,5007
*|5007,5008
<EOL>|5009,5010
IRON|5010,5014
-|5014,5015
61|5015,5017
<EOL>|5017,5018
_|5018,5019
_|5019,5020
_|5020,5021
12|5022,5024
:|5024,5025
30PM|5025,5029
calTIBC|5032,5039
-|5039,5040
303|5040,5043
FERRITIN|5044,5052
-|5052,5053
155|5053,5056
*|5056,5057
TRF|5058,5061
-|5061,5062
233|5062,5065
<EOL>|5065,5066
_|5066,5067
_|5067,5068
_|5068,5069
12|5070,5072
:|5072,5073
30PM|5073,5077
UREA|5080,5084
N|5085,5086
-|5086,5087
42|5087,5089
*|5089,5090
CREAT|5091,5096
-|5096,5097
2|5097,5098
.|5098,5099
3|5099,5100
*|5100,5101
SODIUM|5102,5108
-|5108,5109
142|5109,5112
<EOL>|5113,5114
POTASSIUM|5114,5123
-|5123,5124
4.7|5124,5127
CHLORIDE|5128,5136
-|5136,5137
109|5137,5140
*|5140,5141
TOTAL|5142,5147
CO2|5148,5151
-|5151,5152
23|5152,5154
ANION|5155,5160
GAP|5161,5164
-|5164,5165
15|5165,5167
<EOL>|5167,5168
_|5168,5169
_|5169,5170
_|5170,5171
04|5172,5174
:|5174,5175
50PM|5175,5179
LD|5182,5184
(|5184,5185
_|5185,5186
_|5186,5187
_|5187,5188
)|5188,5189
-|5189,5190
247|5190,5193
TOT|5194,5197
BILI|5198,5202
-|5202,5203
0.2|5203,5206
<EOL>|5206,5207
_|5207,5208
_|5208,5209
_|5209,5210
04|5211,5213
:|5213,5214
50PM|5214,5218
HAPTOGLOB|5221,5230
-|5230,5231
188|5231,5234
<EOL>|5234,5235
<EOL>|5235,5236
IMAGING|5236,5243
:|5243,5244
<EOL>|5246,5247
=|5247,5248
=|5248,5249
=|5249,5250
=|5250,5251
=|5251,5252
=|5252,5253
=|5253,5254
=|5254,5255
=|5255,5256
=|5256,5257
=|5257,5258
=|5258,5259
=|5259,5260
=|5260,5261
=|5261,5262
=|5262,5263
=|5263,5264
=|5264,5265
=|5265,5266
=|5266,5267
=|5267,5268
=|5268,5269
=|5269,5270
=|5270,5271
=|5271,5272
=|5272,5273
=|5273,5274
=|5274,5275
=|5275,5276
=|5276,5277
=|5277,5278
=|5278,5279
=|5279,5280
=|5280,5281
=|5281,5282
=|5282,5283
=|5283,5284
=|5284,5285
=|5285,5286
=|5286,5287
=|5287,5288
=|5288,5289
=|5289,5290
=|5290,5291
=|5291,5292
=|5292,5293
<EOL>|5293,5294
LENIs|5294,5299
(|5300,5301
_|5301,5302
_|5302,5303
_|5303,5304
)|5304,5305
<EOL>|5305,5306
1.|5306,5308
Nonocclusive|5309,5321
deep|5322,5326
vein|5327,5331
thrombosis|5332,5342
of|5343,5345
one|5346,5349
of|5350,5352
the|5353,5356
paired|5357,5363
<EOL>|5364,5365
posterior|5365,5374
tibial|5375,5381
veins|5382,5387
bilaterally|5388,5399
.|5399,5400
The|5402,5405
extent|5406,5412
of|5413,5415
thrombus|5416,5424
<EOL>|5425,5426
bilaterally|5426,5437
has|5438,5441
decreased|5442,5451
.|5451,5452
No|5454,5456
new|5457,5460
deep|5461,5465
venous|5466,5472
thrombosis|5473,5483
in|5484,5486
<EOL>|5487,5488
either|5488,5494
lower|5495,5500
extremity|5501,5510
.|5510,5511
<EOL>|5512,5513
2.|5513,5515
Right|5516,5521
complex|5522,5529
_|5530,5531
_|5531,5532
_|5532,5533
cyst|5534,5538
.|5538,5539
<EOL>|5540,5541
<EOL>|5541,5542
CXR|5542,5545
(|5546,5547
_|5547,5548
_|5548,5549
_|5549,5550
)|5550,5551
:|5551,5552
<EOL>|5553,5554
1.|5554,5556
New|5557,5560
mild|5561,5565
pulmonary|5566,5575
edema|5576,5581
with|5582,5586
persistent|5587,5597
small|5598,5603
bilateral|5604,5613
<EOL>|5614,5615
pleural|5615,5622
effusions|5623,5632
.|5632,5633
<EOL>|5634,5635
2.|5635,5637
Severe|5638,5644
cardiomegaly|5645,5657
is|5658,5660
likely|5661,5667
accentuated|5668,5679
due|5680,5683
to|5684,5686
low|5687,5690
lung|5691,5695
<EOL>|5696,5697
volumes|5697,5704
and|5705,5708
patient|5709,5716
positioning|5717,5728
.|5728,5729
<EOL>|5730,5731
<EOL>|5731,5732
CXR|5732,5735
(|5736,5737
_|5737,5738
_|5738,5739
_|5739,5740
)|5740,5741
:|5741,5742
<EOL>|5742,5743
As|5743,5745
compared|5746,5754
to|5755,5757
_|5758,5759
_|5759,5760
_|5760,5761
,|5761,5762
the|5763,5766
lung|5767,5771
volumes|5772,5779
have|5780,5784
slightly|5785,5793
<EOL>|5794,5795
decreased|5795,5804
.|5804,5805
Signs|5807,5812
of|5813,5815
mild|5816,5820
overinflation|5821,5834
and|5835,5838
moderate|5839,5847
pleural|5848,5855
<EOL>|5856,5857
effusions|5857,5866
persist|5867,5874
.|5874,5875
Moderate|5877,5885
cardiomegaly|5886,5898
.|5898,5899
Elongation|5901,5911
of|5912,5914
the|5915,5918
<EOL>|5919,5920
descending|5920,5930
aorta|5931,5936
.|5936,5937
No|5939,5941
pneumonia|5942,5951
.|5951,5952
<EOL>|5953,5954
<EOL>|5954,5955
LABORAROTY|5955,5965
STUDIES|5966,5973
ON|5974,5976
DISCHARGE|5977,5986
<EOL>|5986,5987
=|5987,5988
=|5988,5989
=|5989,5990
=|5990,5991
=|5991,5992
=|5992,5993
=|5993,5994
=|5994,5995
=|5995,5996
=|5996,5997
=|5997,5998
=|5998,5999
=|5999,6000
=|6000,6001
=|6001,6002
=|6002,6003
=|6003,6004
=|6004,6005
=|6005,6006
=|6006,6007
=|6007,6008
=|6008,6009
=|6009,6010
=|6010,6011
=|6011,6012
=|6012,6013
=|6013,6014
=|6014,6015
=|6015,6016
=|6016,6017
=|6017,6018
=|6018,6019
=|6019,6020
=|6020,6021
=|6021,6022
=|6022,6023
=|6023,6024
=|6024,6025
=|6025,6026
=|6026,6027
=|6027,6028
=|6028,6029
=|6029,6030
=|6030,6031
=|6031,6032
=|6032,6033
<EOL>|6033,6034
_|6034,6035
_|6035,6036
_|6036,6037
05|6038,6040
:|6040,6041
45AM|6041,6045
BLOOD|6046,6051
WBC|6052,6055
-|6055,6056
3|6056,6057
.|6057,6058
4|6058,6059
*|6059,6060
RBC|6061,6064
-|6064,6065
2|6065,6066
.|6066,6067
93|6067,6069
*|6069,6070
Hgb|6071,6074
-|6074,6075
8|6075,6076
.|6076,6077
9|6077,6078
*|6078,6079
Hct|6080,6083
-|6083,6084
28|6084,6086
.|6086,6087
0|6087,6088
*|6088,6089
<EOL>|6090,6091
MCV|6091,6094
-|6094,6095
96|6095,6097
MCH|6098,6101
-|6101,6102
30.4|6102,6106
MCHC|6107,6111
-|6111,6112
31|6112,6114
.|6114,6115
8|6115,6116
*|6116,6117
RDW|6118,6121
-|6121,6122
17|6122,6124
.|6124,6125
5|6125,6126
*|6126,6127
RDWSD|6128,6133
-|6133,6134
59|6134,6136
.|6136,6137
7|6137,6138
*|6138,6139
Plt|6140,6143
_|6144,6145
_|6145,6146
_|6146,6147
<EOL>|6147,6148
_|6148,6149
_|6149,6150
_|6150,6151
05|6152,6154
:|6154,6155
45AM|6155,6159
BLOOD|6160,6165
_|6166,6167
_|6167,6168
_|6168,6169
PTT|6170,6173
-|6173,6174
30.6|6174,6178
_|6179,6180
_|6180,6181
_|6181,6182
<EOL>|6182,6183
_|6183,6184
_|6184,6185
_|6185,6186
05|6187,6189
:|6189,6190
45AM|6190,6194
BLOOD|6195,6200
Glucose|6201,6208
-|6208,6209
116|6209,6212
*|6212,6213
UreaN|6214,6219
-|6219,6220
41|6220,6222
*|6222,6223
Creat|6224,6229
-|6229,6230
2|6230,6231
.|6231,6232
1|6232,6233
*|6233,6234
Na|6235,6237
-|6237,6238
144|6238,6241
<EOL>|6242,6243
K|6243,6244
-|6244,6245
4.0|6245,6248
Cl|6249,6251
-|6251,6252
108|6252,6255
HCO3|6256,6260
-|6260,6261
25|6261,6263
AnGap|6264,6269
-|6269,6270
15|6270,6272
<EOL>|6272,6273
_|6273,6274
_|6274,6275
_|6275,6276
04|6277,6279
:|6279,6280
50PM|6280,6284
BLOOD|6285,6290
LD|6291,6293
(|6293,6294
LDH|6294,6297
)|6297,6298
-|6298,6299
247|6299,6302
TotBili|6303,6310
-|6310,6311
0.2|6311,6314
<EOL>|6314,6315
_|6315,6316
_|6316,6317
_|6317,6318
05|6319,6321
:|6321,6322
45AM|6322,6326
BLOOD|6327,6332
Calcium|6333,6340
-|6340,6341
9.4|6341,6344
Phos|6345,6349
-|6349,6350
4|6350,6351
.|6351,6352
7|6352,6353
*|6353,6354
Mg|6355,6357
-|6357,6358
1.7|6358,6361
<EOL>|6361,6362
<EOL>|6363,6364
Brief|6364,6369
Hospital|6370,6378
Course|6379,6385
:|6385,6386
<EOL>|6386,6387
Ms.|6387,6390
_|6391,6392
_|6392,6393
_|6393,6394
is|6395,6397
a|6398,6399
_|6400,6401
_|6401,6402
_|6402,6403
year|6404,6408
old|6409,6412
woman|6413,6418
with|6419,6423
a|6424,6425
past|6426,6430
medical|6431,6438
<EOL>|6439,6440
history|6440,6447
of|6448,6450
type|6451,6455
-|6455,6456
2|6456,6457
DM|6458,6460
,|6460,6461
hypertension|6462,6474
,|6474,6475
stage|6476,6481
IV|6482,6484
CKD|6485,6488
,|6488,6489
CAD|6490,6493
s|6494,6495
/|6495,6496
p|6496,6497
<EOL>|6498,6499
distant|6499,6506
MI|6507,6509
and|6510,6513
bare|6514,6518
metal|6519,6524
stent|6525,6530
,|6530,6531
stroke|6532,6538
,|6538,6539
recent|6540,6546
unprovoked|6547,6557
DVTs|6558,6562
<EOL>|6563,6564
on|6564,6566
Coumadin|6567,6575
,|6575,6576
and|6577,6580
recent|6581,6587
upper|6588,6593
GI|6594,6596
bleed|6597,6602
,|6602,6603
who|6604,6607
was|6608,6611
sent|6612,6616
to|6617,6619
_|6620,6621
_|6621,6622
_|6622,6623
by|6624,6626
<EOL>|6627,6628
her|6628,6631
physician|6632,6641
for|6642,6645
anemia|6646,6652
.|6652,6653
<EOL>|6654,6655
<EOL>|6655,6656
#|6656,6657
Anemia|6658,6664
:|6664,6665
<EOL>|6666,6667
Patient|6667,6674
presented|6675,6684
with|6685,6689
Hgb|6690,6693
of|6694,6696
6.5|6697,6700
,|6700,6701
down|6702,6706
from|6707,6711
her|6712,6715
recent|6716,6722
baseline|6723,6731
<EOL>|6732,6733
of|6733,6735
~|6736,6737
7.5|6737,6740
since|6741,6746
her|6747,6750
_|6751,6752
_|6752,6753
_|6753,6754
hospitalization|6755,6770
.|6770,6771
Upon|6772,6776
presentation|6777,6789
she|6790,6793
<EOL>|6794,6795
had|6795,6798
a|6799,6800
new|6801,6804
macrocytic|6805,6815
anemia|6816,6822
.|6822,6823
Hemolysis|6824,6833
labs|6834,6838
were|6839,6843
negative|6844,6852
.|6852,6853
She|6854,6857
<EOL>|6858,6859
received|6859,6867
two|6868,6871
units|6872,6877
of|6878,6880
packed|6881,6887
red|6888,6891
cells|6892,6897
with|6898,6902
an|6903,6905
appropriate|6906,6917
rise|6918,6922
<EOL>|6923,6924
in|6924,6926
her|6927,6930
Hgb|6931,6934
to|6935,6937
9.0|6938,6941
.|6941,6942
Stool|6943,6948
was|6949,6952
guiac|6953,6958
negative|6959,6967
,|6967,6968
with|6969,6973
no|6974,6976
reports|6977,6984
of|6985,6987
<EOL>|6988,6989
dark|6989,6993
stool|6994,6999
or|7000,7002
blood|7003,7008
in|7009,7011
stool|7012,7017
.|7017,7018
Her|7019,7022
hemoglobin|7023,7033
remained|7034,7042
stable|7043,7049
at|7050,7052
<EOL>|7053,7054
this|7054,7058
level|7059,7064
,|7064,7065
there|7066,7071
was|7072,7075
no|7076,7078
overt|7079,7084
bleeding|7085,7093
,|7093,7094
and|7095,7098
her|7099,7102
stool|7103,7108
was|7109,7112
guiac|7113,7118
<EOL>|7119,7120
negative|7120,7128
.|7128,7129
After|7130,7135
transfusion|7136,7147
the|7148,7151
patient|7152,7159
reported|7160,7168
significant|7169,7180
<EOL>|7181,7182
improvement|7182,7193
in|7194,7196
her|7197,7200
shortness|7201,7210
of|7211,7213
breath|7214,7220
and|7221,7224
fatigue|7225,7232
.|7232,7233
Given|7234,7239
her|7240,7243
<EOL>|7244,7245
history|7245,7252
of|7253,7255
gastritis|7256,7265
and|7266,7269
diverticulosis|7270,7284
,|7284,7285
a|7286,7287
GI|7288,7290
bleed|7291,7296
was|7297,7300
believed|7301,7309
<EOL>|7310,7311
responsible|7311,7322
for|7323,7326
her|7327,7330
anemia|7331,7337
.|7337,7338
Patient|7339,7346
should|7347,7353
receive|7354,7361
an|7362,7364
<EOL>|7365,7366
EGD|7366,7369
/|7369,7370
colonoscopy|7370,7381
as|7382,7384
an|7385,7387
outpatient|7388,7398
.|7398,7399
<EOL>|7400,7401
<EOL>|7401,7402
#|7402,7403
Acute|7404,7409
exacerbation|7410,7422
of|7423,7425
heart|7426,7431
failure|7432,7439
with|7440,7444
preserved|7445,7454
ejection|7455,7463
<EOL>|7464,7465
fraction|7465,7473
:|7473,7474
<EOL>|7475,7476
The|7476,7479
patient|7480,7487
was|7488,7491
also|7492,7496
found|7497,7502
to|7503,7505
be|7506,7508
slightly|7509,7517
volume|7518,7524
overloaded|7525,7535
,|7535,7536
and|7537,7540
<EOL>|7541,7542
was|7542,7545
treated|7546,7553
with|7554,7558
2x40mg|7559,7565
IV|7566,7568
Lasix|7569,7574
,|7574,7575
with|7576,7580
good|7581,7585
urine|7586,7591
output|7592,7598
and|7599,7602
<EOL>|7603,7604
symptomatic|7604,7615
improvement|7616,7627
.|7627,7628
Her|7629,7632
pulmonary|7633,7642
edema|7643,7648
and|7649,7652
peripheral|7653,7663
<EOL>|7664,7665
edema|7665,7670
resolved|7671,7679
with|7680,7684
diuresis|7685,7693
.|7693,7694
<EOL>|7694,7695
<EOL>|7695,7696
CHRONIC|7696,7703
ISSUES|7704,7710
:|7710,7711
<EOL>|7711,7712
#|7712,7713
Gastic|7714,7720
ulceration|7721,7731
:|7731,7732
<EOL>|7733,7734
Continued|7734,7743
on|7744,7746
home|7747,7751
pantoprazole|7752,7764
BID|7765,7768
<EOL>|7768,7769
<EOL>|7769,7770
#|7770,7771
Hypertension|7772,7784
:|7784,7785
<EOL>|7785,7786
Continued|7786,7795
on|7796,7798
home|7799,7803
nifedipine|7804,7814
,|7814,7815
carvadilol|7816,7826
,|7826,7827
lisinopril|7828,7838
.|7838,7839
<EOL>|7839,7840
<EOL>|7840,7841
#|7841,7842
Stage|7843,7848
IV|7849,7851
Chronic|7852,7859
Kidney|7860,7866
Disease|7867,7874
:|7874,7875
<EOL>|7876,7877
Creatinine|7877,7887
remained|7888,7896
at|7897,7899
baseline|7900,7908
(|7909,7910
b|7910,7911
/|7911,7912
l|7912,7913
Cr|7914,7916
2.1|7917,7920
-|7920,7921
2.6|7921,7924
)|7924,7925
during|7926,7932
<EOL>|7933,7934
admission|7934,7943
.|7943,7944
<EOL>|7944,7945
<EOL>|7945,7946
TRANSITIONAL|7946,7958
ISSUES|7959,7965
<EOL>|7965,7966
=|7966,7967
=|7967,7968
=|7968,7969
=|7969,7970
=|7970,7971
=|7971,7972
=|7972,7973
=|7973,7974
=|7974,7975
=|7975,7976
=|7976,7977
=|7977,7978
=|7978,7979
=|7979,7980
=|7980,7981
=|7981,7982
=|7982,7983
=|7983,7984
=|7984,7985
=|7985,7986
=|7986,7987
=|7987,7988
<EOL>|7988,7989
-|7989,7990
-|7990,7991
Patient|7991,7998
's|7998,8000
Anemia|8001,8007
is|8008,8010
thought|8011,8018
to|8019,8021
be|8022,8024
due|8025,8028
to|8029,8031
slow|8032,8036
GI|8037,8039
bleed|8040,8045
given|8046,8051
<EOL>|8052,8053
history|8053,8060
of|8061,8063
gastritis|8064,8073
and|8074,8077
diverticulosis|8078,8092
.|8092,8093
Please|8094,8100
schedule|8101,8109
<EOL>|8110,8111
EGD|8111,8114
/|8114,8115
colonoscopy|8115,8126
within|8127,8133
the|8134,8137
next|8138,8142
month|8143,8148
<EOL>|8148,8149
-|8149,8150
-|8150,8151
Patient|8151,8158
continued|8159,8168
on|8169,8171
Coumadin|8172,8180
for|8181,8184
bilateral|8185,8194
DVTs|8195,8199
;|8199,8200
please|8201,8207
<EOL>|8208,8209
continue|8209,8217
to|8218,8220
weigh|8221,8226
the|8227,8230
risks|8231,8236
and|8237,8240
benefits|8241,8249
of|8250,8252
anticoagulation|8253,8268
<EOL>|8269,8270
given|8270,8275
history|8276,8283
of|8284,8286
bleed|8287,8292
.|8292,8293
<EOL>|8293,8294
-|8294,8295
-|8295,8296
Discharge|8296,8305
weight|8306,8312
:|8312,8313
167.7|8314,8319
<EOL>|8319,8320
<EOL>|8320,8321
#|8321,8322
CONTACT|8323,8330
:|8330,8331
_|8332,8333
_|8333,8334
_|8334,8335
_|8336,8337
_|8337,8338
_|8338,8339
<EOL>|8339,8340
#|8340,8341
CODE|8342,8346
:|8346,8347
full|8348,8352
,|8352,8353
confirmed|8354,8363
<EOL>|8363,8364
<EOL>|8365,8366
Medications|8366,8377
on|8378,8380
Admission|8381,8390
:|8390,8391
<EOL>|8391,8392
The|8392,8395
Preadmission|8396,8408
Medication|8409,8419
list|8420,8424
may|8425,8428
be|8429,8431
inaccurate|8432,8442
and|8443,8446
requires|8447,8455
<EOL>|8456,8457
futher|8457,8463
investigation|8464,8477
.|8477,8478
<EOL>|8478,8479
1.|8479,8481
Allopurinol|8482,8493
_|8494,8495
_|8495,8496
_|8496,8497
mg|8498,8500
PO|8501,8503
EVERY|8504,8509
OTHER|8510,8515
DAY|8516,8519
<EOL>|8520,8521
2.|8521,8523
Aspirin|8524,8531
81|8532,8534
mg|8535,8537
PO|8538,8540
DAILY|8541,8546
<EOL>|8547,8548
3.|8548,8550
Atorvastatin|8551,8563
80|8564,8566
mg|8567,8569
PO|8570,8572
QPM|8573,8576
<EOL>|8577,8578
4.|8578,8580
Carvedilol|8581,8591
12.5|8592,8596
mg|8597,8599
PO|8600,8602
BID|8603,8606
<EOL>|8607,8608
5.|8608,8610
Lisinopril|8611,8621
40|8622,8624
mg|8625,8627
PO|8628,8630
DAILY|8631,8636
<EOL>|8637,8638
6.|8638,8640
Multivitamins|8641,8654
1|8655,8656
TAB|8657,8660
PO|8661,8663
DAILY|8664,8669
<EOL>|8670,8671
7.|8671,8673
NIFEdipine|8674,8684
CR|8685,8687
30|8688,8690
mg|8691,8693
PO|8694,8696
BID|8697,8700
<EOL>|8701,8702
8.|8702,8704
Vitamin|8705,8712
D|8713,8714
_|8715,8716
_|8716,8717
_|8717,8718
UNIT|8719,8723
PO|8724,8726
DAILY|8727,8732
<EOL>|8733,8734
9.|8734,8736
Docusate|8737,8745
Sodium|8746,8752
100|8753,8756
mg|8757,8759
PO|8760,8762
BID|8763,8766
<EOL>|8767,8768
10.|8768,8771
Gabapentin|8772,8782
100|8783,8786
mg|8787,8789
PO|8790,8792
QHS|8793,8796
neuropathic|8797,8808
pain|8809,8813
<EOL>|8814,8815
11|8815,8817
.|8817,8818
Pantoprazole|8819,8831
40|8832,8834
mg|8835,8837
PO|8838,8840
Q12H|8841,8845
<EOL>|8846,8847
12.|8847,8850
Senna|8851,8856
8.6|8857,8860
mg|8861,8863
PO|8864,8866
BID|8867,8870
constipation|8871,8883
<EOL>|8884,8885
13.|8885,8888
Warfarin|8889,8897
4|8898,8899
mg|8900,8902
PO|8903,8905
3X|8906,8908
/|8908,8909
WEEK|8909,8913
(|8914,8915
_|8915,8916
_|8916,8917
_|8917,8918
)|8918,8919
<EOL>|8920,8921
14.|8921,8924
Nitroglycerin|8925,8938
SL|8939,8941
0.3|8942,8945
mg|8946,8948
SL|8949,8951
Q5MIN|8952,8957
:|8957,8958
PRN|8958,8961
chest|8962,8967
pain|8968,8972
<EOL>|8973,8974
15|8974,8976
.|8976,8977
Furosemide|8978,8988
20|8989,8991
mg|8992,8994
PO|8995,8997
DAILY|8998,9003
<EOL>|9004,9005
16|9005,9007
.|9007,9008
Polyethylene|9009,9021
Glycol|9022,9028
17|9029,9031
g|9032,9033
PO|9034,9036
DAILY|9037,9042
<EOL>|9043,9044
17.|9044,9047
Acetaminophen|9048,9061
325|9062,9065
-|9065,9066
650|9066,9069
mg|9070,9072
PO|9073,9075
Q6H|9076,9079
:|9079,9080
PRN|9080,9083
pain|9084,9088
or|9089,9091
fever|9092,9097
<EOL>|9098,9099
18.|9099,9102
Warfarin|9103,9111
3|9112,9113
mg|9114,9116
PO|9117,9119
4X|9120,9122
/|9122,9123
WEEK|9123,9127
(|9128,9129
_|9129,9130
_|9130,9131
_|9131,9132
)|9132,9133
<EOL>|9134,9135
19.|9135,9138
70|9139,9141
/|9141,9142
30|9142,9144
30|9145,9147
Units|9148,9153
Dinner|9154,9160
<EOL>|9160,9161
<EOL>|9161,9162
<EOL>|9163,9164
Discharge|9164,9173
Medications|9174,9185
:|9185,9186
<EOL>|9186,9187
1.|9187,9189
Acetaminophen|9190,9203
325|9204,9207
-|9207,9208
650|9208,9211
mg|9212,9214
PO|9215,9217
Q6H|9218,9221
:|9221,9222
PRN|9222,9225
pain|9226,9230
or|9231,9233
fever|9234,9239
<EOL>|9240,9241
RX|9241,9243
*|9244,9245
acetaminophen|9245,9258
325|9259,9262
mg|9263,9265
_|9266,9267
_|9267,9268
_|9268,9269
tablet|9270,9276
(|9276,9277
s|9277,9278
)|9278,9279
by|9280,9282
mouth|9283,9288
Q6H|9289,9292
:|9292,9293
PRN|9293,9296
Disp|9297,9301
<EOL>|9302,9303
#|9303,9304
*|9304,9305
120|9305,9308
Tablet|9309,9315
Refills|9316,9323
:|9323,9324
*|9324,9325
0|9325,9326
<EOL>|9326,9327
2.|9327,9329
Aspirin|9330,9337
81|9338,9340
mg|9341,9343
PO|9344,9346
DAILY|9347,9352
<EOL>|9353,9354
RX|9354,9356
*|9357,9358
aspirin|9358,9365
81|9366,9368
mg|9369,9371
1|9372,9373
tablet|9374,9380
(|9380,9381
s|9381,9382
)|9382,9383
by|9384,9386
mouth|9387,9392
daily|9393,9398
Disp|9399,9403
#|9404,9405
*|9405,9406
30|9406,9408
Tablet|9409,9415
<EOL>|9416,9417
Refills|9417,9424
:|9424,9425
*|9425,9426
0|9426,9427
<EOL>|9427,9428
3.|9428,9430
Atorvastatin|9431,9443
80|9444,9446
mg|9447,9449
PO|9450,9452
QPM|9453,9456
<EOL>|9457,9458
RX|9458,9460
*|9461,9462
atorvastatin|9462,9474
80|9475,9477
mg|9478,9480
1|9481,9482
tablet|9483,9489
(|9489,9490
s|9490,9491
)|9491,9492
by|9493,9495
mouth|9496,9501
QPM|9502,9505
Disp|9506,9510
#|9511,9512
*|9512,9513
30|9513,9515
Tablet|9516,9522
<EOL>|9523,9524
Refills|9524,9531
:|9531,9532
*|9532,9533
0|9533,9534
<EOL>|9534,9535
4.|9535,9537
Carvedilol|9538,9548
12.5|9549,9553
mg|9554,9556
PO|9557,9559
BID|9560,9563
<EOL>|9564,9565
RX|9565,9567
*|9568,9569
carvedilol|9569,9579
12.5|9580,9584
mg|9585,9587
1|9588,9589
tablet|9590,9596
(|9596,9597
s|9597,9598
)|9598,9599
by|9600,9602
mouth|9603,9608
twice|9609,9614
a|9615,9616
day|9617,9620
Disp|9621,9625
<EOL>|9626,9627
#|9627,9628
*|9628,9629
60|9629,9631
Tablet|9632,9638
Refills|9639,9646
:|9646,9647
*|9647,9648
0|9648,9649
<EOL>|9649,9650
5.|9650,9652
Docusate|9653,9661
Sodium|9662,9668
100|9669,9672
mg|9673,9675
PO|9676,9678
BID|9679,9682
<EOL>|9683,9684
RX|9684,9686
*|9687,9688
docusate|9688,9696
sodium|9697,9703
100|9704,9707
mg|9708,9710
1|9711,9712
capsule|9713,9720
(|9720,9721
s|9721,9722
)|9722,9723
by|9724,9726
mouth|9727,9732
twice|9733,9738
a|9739,9740
day|9741,9744
<EOL>|9745,9746
Disp|9746,9750
#|9751,9752
*|9752,9753
60|9753,9755
Capsule|9756,9763
Refills|9764,9771
:|9771,9772
*|9772,9773
0|9773,9774
<EOL>|9774,9775
6.|9775,9777
Gabapentin|9778,9788
100|9789,9792
mg|9793,9795
PO|9796,9798
QHS|9799,9802
neuropathic|9803,9814
pain|9815,9819
<EOL>|9820,9821
RX|9821,9823
*|9824,9825
gabapentin|9825,9835
100|9836,9839
mg|9840,9842
1|9843,9844
capsule|9845,9852
(|9852,9853
s|9853,9854
)|9854,9855
by|9856,9858
mouth|9859,9864
at|9865,9867
bedtime|9868,9875
Disp|9876,9880
#|9881,9882
*|9882,9883
30|9883,9885
<EOL>|9886,9887
Capsule|9887,9894
Refills|9895,9902
:|9902,9903
*|9903,9904
0|9904,9905
<EOL>|9905,9906
7.|9906,9908
Lisinopril|9909,9919
40|9920,9922
mg|9923,9925
PO|9926,9928
DAILY|9929,9934
<EOL>|9935,9936
RX|9936,9938
*|9939,9940
lisinopril|9940,9950
40|9951,9953
mg|9954,9956
1|9957,9958
tablet|9959,9965
(|9965,9966
s|9966,9967
)|9967,9968
by|9969,9971
mouth|9972,9977
daily|9978,9983
Disp|9984,9988
#|9989,9990
*|9990,9991
30|9991,9993
Tablet|9994,10000
<EOL>|10001,10002
Refills|10002,10009
:|10009,10010
*|10010,10011
0|10011,10012
<EOL>|10012,10013
8.|10013,10015
Multivitamins|10016,10029
1|10030,10031
TAB|10032,10035
PO|10036,10038
DAILY|10039,10044
<EOL>|10045,10046
RX|10046,10048
*|10049,10050
multivitamin|10050,10062
1|10064,10065
capsule|10066,10073
(|10073,10074
s|10074,10075
)|10075,10076
by|10077,10079
mouth|10080,10085
daily|10086,10091
Disp|10092,10096
#|10097,10098
*|10098,10099
30|10099,10101
Capsule|10102,10109
<EOL>|10110,10111
Refills|10111,10118
:|10118,10119
*|10119,10120
0|10120,10121
<EOL>|10121,10122
9.|10122,10124
NIFEdipine|10125,10135
CR|10136,10138
30|10139,10141
mg|10142,10144
PO|10145,10147
BID|10148,10151
<EOL>|10152,10153
RX|10153,10155
*|10156,10157
nifedipine|10157,10167
30|10168,10170
mg|10171,10173
1|10174,10175
tablet|10176,10182
(|10182,10183
s|10183,10184
)|10184,10185
by|10186,10188
mouth|10189,10194
twice|10195,10200
a|10201,10202
day|10203,10206
Disp|10207,10211
#|10212,10213
*|10213,10214
60|10214,10216
<EOL>|10217,10218
Tablet|10218,10224
Refills|10225,10232
:|10232,10233
*|10233,10234
0|10234,10235
<EOL>|10235,10236
10.|10236,10239
Nitroglycerin|10240,10253
SL|10254,10256
0.3|10257,10260
mg|10261,10263
SL|10264,10266
Q5MIN|10267,10272
:|10272,10273
PRN|10273,10276
chest|10277,10282
pain|10283,10287
<EOL>|10288,10289
RX|10289,10291
*|10292,10293
nitroglycerin|10293,10306
[|10307,10308
Nitrostat|10308,10317
]|10317,10318
0.3|10319,10322
mg|10323,10325
1|10326,10327
tablet|10328,10334
(|10334,10335
s|10335,10336
)|10336,10337
sublingually|10338,10350
<EOL>|10351,10352
Q5MIN|10352,10357
:|10357,10358
PRN|10358,10361
Disp|10362,10366
#|10367,10368
*|10368,10369
10|10369,10371
Tablet|10372,10378
Refills|10379,10386
:|10386,10387
*|10387,10388
0|10388,10389
<EOL>|10389,10390
11.|10390,10393
Pantoprazole|10394,10406
40|10407,10409
mg|10410,10412
PO|10413,10415
Q12H|10416,10420
<EOL>|10421,10422
RX|10422,10424
*|10425,10426
pantoprazole|10426,10438
40|10439,10441
mg|10442,10444
1|10445,10446
tablet|10447,10453
(|10453,10454
s|10454,10455
)|10455,10456
by|10457,10459
mouth|10460,10465
every|10466,10471
twelve|10472,10478
(|10479,10480
12|10480,10482
)|10482,10483
<EOL>|10484,10485
hours|10485,10490
Disp|10491,10495
#|10496,10497
*|10497,10498
60|10498,10500
Tablet|10501,10507
Refills|10508,10515
:|10515,10516
*|10516,10517
0|10517,10518
<EOL>|10518,10519
12.|10519,10522
Polyethylene|10523,10535
Glycol|10536,10542
17|10543,10545
g|10546,10547
PO|10548,10550
DAILY|10551,10556
<EOL>|10557,10558
RX|10558,10560
*|10561,10562
polyethylene|10562,10574
glycol|10575,10581
3350|10582,10586
17|10587,10589
gram|10590,10594
/|10594,10595
dose|10595,10599
1|10600,10601
powder|10602,10608
(|10608,10609
s|10609,10610
)|10610,10611
by|10612,10614
mouth|10615,10620
<EOL>|10621,10622
daily|10622,10627
Refills|10628,10635
:|10635,10636
*|10636,10637
0|10637,10638
<EOL>|10638,10639
13.|10639,10642
Senna|10643,10648
8.6|10649,10652
mg|10653,10655
PO|10656,10658
BID|10659,10662
constipation|10663,10675
<EOL>|10676,10677
RX|10677,10679
*|10680,10681
sennosides|10681,10691
[|10692,10693
senna|10693,10698
]|10698,10699
8.6|10700,10703
mg|10704,10706
1|10707,10708
capsule|10709,10716
by|10717,10719
mouth|10720,10725
twice|10726,10731
a|10732,10733
day|10734,10737
<EOL>|10738,10739
Disp|10739,10743
#|10744,10745
*|10745,10746
60|10746,10748
Capsule|10749,10756
Refills|10757,10764
:|10764,10765
*|10765,10766
0|10766,10767
<EOL>|10767,10768
14.|10768,10771
Vitamin|10772,10779
D|10780,10781
_|10782,10783
_|10783,10784
_|10784,10785
UNIT|10786,10790
PO|10791,10793
DAILY|10794,10799
<EOL>|10800,10801
RX|10801,10803
*|10804,10805
ergocalciferol|10805,10819
(|10820,10821
vitamin|10821,10828
D2|10829,10831
)|10831,10832
2,000|10833,10838
unit|10839,10843
1|10844,10845
tablet|10846,10852
(|10852,10853
s|10853,10854
)|10854,10855
by|10856,10858
mouth|10859,10864
<EOL>|10865,10866
daily|10866,10871
Disp|10872,10876
#|10877,10878
*|10878,10879
30|10879,10881
Tablet|10882,10888
Refills|10889,10896
:|10896,10897
*|10897,10898
0|10898,10899
<EOL>|10899,10900
15.|10900,10903
Warfarin|10904,10912
4|10913,10914
mg|10915,10917
PO|10918,10920
3X|10921,10923
/|10923,10924
WEEK|10924,10928
(|10929,10930
_|10930,10931
_|10931,10932
_|10932,10933
)|10933,10934
<EOL>|10935,10936
RX|10936,10938
*|10939,10940
warfarin|10940,10948
4|10949,10950
mg|10951,10953
1|10954,10955
tablet|10956,10962
(|10962,10963
s|10963,10964
)|10964,10965
by|10966,10968
mouth|10969,10974
3X|10975,10977
/|10977,10978
WEEK|10978,10982
Disp|10983,10987
#|10988,10989
*|10989,10990
30|10990,10992
Tablet|10993,10999
<EOL>|11000,11001
Refills|11001,11008
:|11008,11009
*|11009,11010
0|11010,11011
<EOL>|11011,11012
16|11012,11014
.|11014,11015
Warfarin|11016,11024
3|11025,11026
mg|11027,11029
PO|11030,11032
4X|11033,11035
/|11035,11036
WEEK|11036,11040
(|11041,11042
_|11042,11043
_|11043,11044
_|11044,11045
)|11045,11046
<EOL>|11047,11048
RX|11048,11050
*|11051,11052
warfarin|11052,11060
3|11061,11062
mg|11063,11065
1|11066,11067
tablet|11068,11074
(|11074,11075
s|11075,11076
)|11076,11077
by|11078,11080
mouth|11081,11086
4X|11087,11089
/|11089,11090
WEEK|11090,11094
Disp|11095,11099
#|11100,11101
*|11101,11102
30|11102,11104
Tablet|11105,11111
<EOL>|11112,11113
Refills|11113,11120
:|11120,11121
*|11121,11122
0|11122,11123
<EOL>|11123,11124
17.|11124,11127
Furosemide|11128,11138
20|11139,11141
mg|11142,11144
PO|11145,11147
DAILY|11148,11153
<EOL>|11154,11155
RX|11155,11157
*|11158,11159
furosemide|11159,11169
20|11170,11172
mg|11173,11175
1|11176,11177
tablet|11178,11184
(|11184,11185
s|11185,11186
)|11186,11187
by|11188,11190
mouth|11191,11196
daily|11197,11202
Disp|11203,11207
#|11208,11209
*|11209,11210
30|11210,11212
Tablet|11213,11219
<EOL>|11220,11221
Refills|11221,11228
:|11228,11229
*|11229,11230
0|11230,11231
<EOL>|11231,11232
18.|11232,11235
Allopurinol|11236,11247
_|11248,11249
_|11249,11250
_|11250,11251
mg|11252,11254
PO|11255,11257
EVERY|11258,11263
OTHER|11264,11269
DAY|11270,11273
<EOL>|11274,11275
RX|11275,11277
*|11278,11279
allopurinol|11279,11290
_|11291,11292
_|11292,11293
_|11293,11294
mg|11295,11297
1|11298,11299
tablet|11300,11306
(|11306,11307
s|11307,11308
)|11308,11309
by|11310,11312
mouth|11313,11318
EVERY|11319,11324
OTHER|11325,11330
DAY|11331,11334
Disp|11335,11339
<EOL>|11340,11341
#|11341,11342
*|11342,11343
30|11343,11345
Tablet|11346,11352
Refills|11353,11360
:|11360,11361
*|11361,11362
0|11362,11363
<EOL>|11363,11364
19.|11364,11367
70|11368,11370
/|11370,11371
30|11371,11373
30|11374,11376
Units|11377,11382
Dinner|11383,11389
<EOL>|11389,11390
RX|11390,11392
*|11393,11394
insulin|11394,11401
NPH|11402,11405
and|11406,11409
regular|11410,11417
human|11418,11423
[|11424,11425
Humulin|11425,11432
70|11433,11435
/|11435,11436
30|11436,11438
KwikPen|11439,11446
]|11446,11447
100|11448,11451
<EOL>|11452,11453
unit|11453,11457
/|11457,11458
mL|11458,11460
(|11461,11462
70|11462,11464
-|11464,11465
30|11465,11467
)|11467,11468
30|11469,11471
units|11472,11477
SC|11478,11480
Take|11481,11485
30|11486,11488
Units|11489,11494
before|11495,11501
DINER|11502,11507
Disp|11508,11512
#|11513,11514
*|11514,11515
2|11515,11516
<EOL>|11517,11518
Package|11518,11525
Refills|11526,11533
:|11533,11534
*|11534,11535
0|11535,11536
<EOL>|11536,11537
<EOL>|11537,11538
<EOL>|11539,11540
Discharge|11540,11549
Disposition|11550,11561
:|11561,11562
<EOL>|11562,11563
Home|11563,11567
With|11568,11572
Service|11573,11580
<EOL>|11580,11581
<EOL>|11582,11583
Facility|11583,11591
:|11591,11592
<EOL>|11592,11593
_|11593,11594
_|11594,11595
_|11595,11596
<EOL>|11596,11597
<EOL>|11598,11599
Discharge|11599,11608
Diagnosis|11609,11618
:|11618,11619
<EOL>|11619,11620
Primary|11620,11627
diagnosis|11628,11637
:|11637,11638
<EOL>|11638,11639
Anemia|11639,11645
<EOL>|11645,11646
Congestive|11646,11656
heart|11657,11662
failure|11663,11670
exacerbation|11671,11683
<EOL>|11683,11684
<EOL>|11684,11685
Secondary|11685,11694
diagnosis|11695,11704
:|11704,11705
<EOL>|11705,11706
Hypertension|11706,11718
<EOL>|11719,11720
DMII|11720,11724
on|11725,11727
insulin|11728,11735
<EOL>|11736,11737
Coronary|11737,11745
artery|11746,11752
disease|11753,11760
<EOL>|11761,11762
Stage|11762,11767
IV|11768,11770
chronic|11771,11778
kidney|11779,11785
disease|11786,11793
<EOL>|11793,11794
Deep|11794,11798
vein|11799,11803
thrombosis|11804,11814
<EOL>|11814,11815
<EOL>|11815,11816
<EOL>|11817,11818
Discharge|11818,11827
Condition|11828,11837
:|11837,11838
<EOL>|11838,11839
Mental|11839,11845
Status|11846,11852
:|11852,11853
Clear|11854,11859
and|11860,11863
coherent|11864,11872
.|11872,11873
<EOL>|11873,11874
Level|11874,11879
of|11880,11882
Consciousness|11883,11896
:|11896,11897
Alert|11898,11903
and|11904,11907
interactive|11908,11919
.|11919,11920
<EOL>|11920,11921
Activity|11921,11929
Status|11930,11936
:|11936,11937
Ambulatory|11938,11948
-|11949,11950
requires|11951,11959
assistance|11960,11970
or|11971,11973
aid|11974,11977
(|11978,11979
walker|11979,11985
<EOL>|11986,11987
or|11987,11989
cane|11990,11994
)|11994,11995
.|11995,11996
<EOL>|11996,11997
<EOL>|11997,11998
<EOL>|11999,12000
Discharge|12000,12009
Instructions|12010,12022
:|12022,12023
<EOL>|12023,12024
Dear|12024,12028
_|12029,12030
_|12030,12031
_|12031,12032
,|12032,12033
<EOL>|12033,12034
<EOL>|12034,12035
It|12035,12037
was|12038,12041
a|12042,12043
pleasure|12044,12052
caring|12053,12059
for|12060,12063
you|12064,12067
.|12067,12068
You|12069,12072
were|12073,12077
admitted|12078,12086
to|12087,12089
the|12090,12093
<EOL>|12094,12095
hospital|12095,12103
with|12104,12108
fatigue|12109,12116
,|12116,12117
chest|12118,12123
pain|12124,12128
,|12128,12129
and|12130,12133
shortness|12134,12143
of|12144,12146
breath|12147,12153
.|12153,12154
You|12155,12158
<EOL>|12159,12160
were|12160,12164
found|12165,12170
to|12171,12173
have|12174,12178
too|12179,12182
few|12183,12186
red|12187,12190
blood|12191,12196
cells|12197,12202
(|12203,12204
anemia|12204,12210
)|12210,12211
.|12211,12212
We|12213,12215
gave|12216,12220
you|12221,12224
<EOL>|12225,12226
blood|12226,12231
,|12231,12232
and|12233,12236
your|12237,12241
symptoms|12242,12250
improved|12251,12259
.|12259,12260
Additionally|12261,12273
,|12273,12274
you|12275,12278
were|12279,12283
found|12284,12289
<EOL>|12290,12291
to|12291,12293
have|12294,12298
too|12299,12302
much|12303,12307
fluid|12308,12313
in|12314,12316
your|12317,12321
legs|12322,12326
and|12327,12330
lungs|12331,12336
.|12336,12337
We|12338,12340
treated|12341,12348
you|12349,12352
<EOL>|12353,12354
with|12354,12358
a|12359,12360
diuretic|12361,12369
,|12369,12370
which|12371,12376
helped|12377,12383
eliminate|12384,12393
the|12394,12397
fluid|12398,12403
.|12403,12404
<EOL>|12405,12406
<EOL>|12406,12407
Weigh|12407,12412
yourself|12413,12421
every|12422,12427
morning|12428,12435
,|12435,12436
call|12437,12441
MD|12442,12444
if|12445,12447
weight|12448,12454
goes|12455,12459
up|12460,12462
more|12463,12467
<EOL>|12468,12469
than|12469,12473
3|12474,12475
lbs|12476,12479
.|12479,12480
<EOL>|12480,12481
<EOL>|12481,12482
Sincerely|12482,12491
,|12491,12492
<EOL>|12492,12493
Your|12493,12497
_|12498,12499
_|12499,12500
_|12500,12501
Team|12502,12506
<EOL>|12506,12507
<EOL>|12508,12509
Followup|12509,12517
Instructions|12518,12530
:|12530,12531
<EOL>|12531,12532
_|12532,12533
_|12533,12534
_|12534,12535
<EOL>|12535,12536

