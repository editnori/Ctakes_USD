 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|184,193|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|184,193|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|196,218|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|204,208|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|204,208|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|204,218|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|221,230|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|256,261|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Chief Complaint|256,261|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Chief Complaint|256,266|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Chief Complaint|256,266|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Chief Complaint|262,266|false|true|false|C2598155||Pain
Finding|Functional Concept|Chief Complaint|262,266|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Chief Complaint|262,266|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Classification|Chief Complaint|271,276|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|277,285|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|289,307|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|298,307|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|298,307|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|298,307|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|298,307|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|381,388|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|381,391|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|393,405|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|History of Present Illness|407,413|false|false|false|C0004096|Asthma|asthma
Attribute|Clinical Attribute|History of Present Illness|425,434|false|false|false|C0945731||diagnosis
Finding|Classification|History of Present Illness|425,434|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|History of Present Illness|425,434|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|History of Present Illness|425,434|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|History of Present Illness|438,441|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|438,441|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|438,441|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|438,441|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|438,441|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|438,441|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|438,441|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|History of Present Illness|451,457|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|History of Present Illness|451,457|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|History of Present Illness|451,457|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|History of Present Illness|451,457|false|false|false|C0038435|Stress|stress
Procedure|Health Care Activity|History of Present Illness|459,463|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|459,463|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Idea or Concept|History of Present Illness|477,484|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|History of Present Illness|477,484|false|false|false|C0039869;C4319827|Thought|thought
Finding|Finding|History of Present Illness|491,497|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Disorder|Disease or Syndrome|History of Present Illness|491,512|false|false|false|C0856737|Single vessel disease|single vessel disease
Anatomy|Body Location or Region|History of Present Illness|498,504|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|498,504|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|History of Present Illness|505,512|false|true|false|C0012634|Disease|disease
Anatomy|Body Location or Region|History of Present Illness|545,550|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|545,550|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|545,555|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|545,555|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|551,555|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|551,555|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|551,555|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|573,582|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|History of Present Illness|573,582|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|History of Present Illness|573,582|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|History of Present Illness|573,582|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|History of Present Illness|603,625|false|false|false|C0745043|History of recent hospitalization|recent hospitalization
Procedure|Health Care Activity|History of Present Illness|610,625|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Classification|History of Present Illness|666,674|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|666,674|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|666,674|false|false|false|C5237010|Expression Negative|negative
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|683,690|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|History of Present Illness|683,690|false|false|false|C1314974|Cardiac attachment|cardiac
Attribute|Clinical Attribute|History of Present Illness|683,698|false|false|false|C2926589||cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|683,698|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Drug|Enzyme|History of Present Illness|683,698|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Procedure|Laboratory Procedure|History of Present Illness|683,698|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|691,698|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|History of Present Illness|691,698|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|History of Present Illness|691,698|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Finding|Functional Concept|History of Present Illness|691,698|false|false|false|C0014445|enzymology|enzymes
Attribute|Clinical Attribute|History of Present Illness|711,717|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|History of Present Illness|711,717|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|History of Present Illness|711,717|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|History of Present Illness|711,717|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|History of Present Illness|711,722|false|false|false|C0920208|Echocardiography, Stress|stress echo
Procedure|Health Care Activity|History of Present Illness|718,722|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|718,722|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Functional Concept|History of Present Illness|736,745|false|false|false|C0205263|Induce (action)|inducible
Finding|Pathologic Function|History of Present Illness|746,754|false|true|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|746,754|false|true|false|C4321499|Ischemia Procedure|ischemia
Finding|Finding|History of Present Illness|762,770|false|false|false|C5453128|Achieved|achieved
Finding|Idea or Concept|History of Present Illness|782,789|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|History of Present Illness|782,789|false|false|false|C0039869;C4319827|Thought|thought
Finding|Finding|History of Present Illness|796,802|false|false|false|C0087136;C1549113|Marital Status - Single;Unmarried|single
Disorder|Disease or Syndrome|History of Present Illness|796,817|false|false|false|C0856737|Single vessel disease|single vessel disease
Anatomy|Body Location or Region|History of Present Illness|803,809|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|803,809|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|History of Present Illness|810,817|false|true|false|C0012634|Disease|disease
Procedure|Health Care Activity|History of Present Illness|826,830|false|true|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|826,830|false|true|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Attribute|Clinical Attribute|History of Present Illness|832,838|false|false|false|C4255046||report
Finding|Intellectual Product|History of Present Illness|832,838|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|832,838|false|false|false|C0700287|Reporting|report
Finding|Finding|History of Present Illness|848,852|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|848,852|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|848,852|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|History of Present Illness|857,861|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|History of Present Illness|857,861|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|History of Present Illness|857,861|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|History of Present Illness|857,861|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Functional Concept|History of Present Illness|870,877|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|History of Present Illness|870,877|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|History of Present Illness|870,877|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|History of Present Illness|870,877|false|false|false|C0199168|Medical service|medical
Event|Occupational Activity|History of Present Illness|878,888|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|878,888|false|false|false|C0376636|Disease Management|management
Finding|Finding|History of Present Illness|901,907|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|901,907|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|919,928|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|History of Present Illness|919,928|false|false|false|C2707265||pulmonary
Finding|Finding|History of Present Illness|919,928|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Disorder|Disease or Syndrome|History of Present Illness|919,936|false|false|false|C0024115|Lung diseases|pulmonary disease
Finding|Finding|History of Present Illness|919,936|false|false|false|C0455540|History of - respiratory disease|pulmonary disease
Disorder|Disease or Syndrome|History of Present Illness|929,936|false|false|false|C0012634|Disease|disease
Finding|Intellectual Product|History of Present Illness|963,967|false|false|false|C0439096|Greek letter beta|beta
Drug|Pharmacologic Substance|History of Present Illness|963,975|false|false|false|C0001645|Adrenergic beta-Antagonists|beta blocker
Drug|Organic Chemical|History of Present Illness|996,1005|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|History of Present Illness|996,1005|false|false|false|C0012373|diltiazem|diltiazem
Procedure|Health Care Activity|History of Present Illness|1037,1046|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|History of Present Illness|1095,1098|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Gene or Genome|History of Present Illness|1095,1098|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Intellectual Product|History of Present Illness|1095,1098|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Molecular Function|History of Present Illness|1095,1098|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Idea or Concept|History of Present Illness|1121,1126|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Intellectual Product|History of Present Illness|1121,1126|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Idea or Concept|History of Present Illness|1140,1144|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|1140,1144|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Finding|History of Present Illness|1163,1172|false|false|false|C3842677|Very hard|very hard
Finding|Finding|History of Present Illness|1176,1183|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|History of Present Illness|1176,1183|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Idea or Concept|History of Present Illness|1263,1268|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Finding|Intellectual Product|History of Present Illness|1263,1268|false|false|false|C1515258;C1547567;C1548343;C1576870|Authorization Mode - Phone;MDFAttributeType - Phone;Telephone Number;Visit User Code - Phone|phone
Anatomy|Body Location or Region|History of Present Illness|1299,1304|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1299,1304|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1299,1309|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1299,1309|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1305,1309|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1305,1309|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1305,1309|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1315,1319|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1315,1319|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1315,1319|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|1342,1347|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1342,1347|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|1354,1358|false|false|false|C0278144|Dull pain|dull
Finding|Sign or Symptom|History of Present Illness|1354,1363|false|false|false|C0278144|Dull pain|dull pain
Attribute|Clinical Attribute|History of Present Illness|1359,1363|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1359,1363|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1359,1363|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|History of Present Illness|1364,1368|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Functional Concept|History of Present Illness|1385,1389|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|1391,1399|false|false|false|C0037004;C4299050|Shoulder;Upper extremity>Shoulder|shoulder
Procedure|Diagnostic Procedure|History of Present Illness|1391,1399|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1391,1399|false|false|false|C0221590;C0869975|Examination of shoulder(s);Procedures on Shoulder|shoulder
Finding|Functional Concept|History of Present Illness|1414,1418|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1414,1425|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1419,1425|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|1419,1425|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|1419,1425|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1419,1425|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|History of Present Illness|1478,1485|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|History of Present Illness|1481,1485|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1481,1485|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1481,1485|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|History of Present Illness|1497,1502|false|false|false|C1446899|minor (disease)|minor
Finding|Gene or Genome|History of Present Illness|1497,1502|false|false|false|C1417837;C3272493|NR4A3 gene;NR4A3 wt Allele|minor
Finding|Conceptual Entity|History of Present Illness|1503,1514|false|false|false|C2986411|Improvement|improvement
Finding|Sign or Symptom|History of Present Illness|1624,1627|false|false|false|C0013404|Dyspnea|SOB
Attribute|Clinical Attribute|History of Present Illness|1630,1636|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|1630,1636|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|1630,1645|false|false|false|C0027498|Nausea and vomiting|nausea/vomiting
Finding|Sign or Symptom|History of Present Illness|1637,1645|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|History of Present Illness|1662,1671|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|1662,1671|true|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Disorder|Disease or Syndrome|History of Present Illness|1673,1676|true|false|false|C1956415|Paroxysmal nocturnal dyspnea|PND
Finding|Gene or Genome|History of Present Illness|1673,1676|true|false|false|C1417807;C4552608|NPPA gene;NPPA wt Allele|PND
Attribute|Clinical Attribute|History of Present Illness|1682,1687|true|false|false|C1717255||edema
Finding|Pathologic Function|History of Present Illness|1682,1687|true|false|false|C0013604|Edema|edema
Finding|Finding|History of Present Illness|1692,1704|false|false|false|C0030252|Palpitations|palpitations
Finding|Idea or Concept|History of Present Illness|1723,1730|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Intellectual Product|History of Present Illness|1781,1784|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1781,1784|false|false|false|C1623258|Electrocardiography|EKG
Disorder|Disease or Syndrome|History of Present Illness|1791,1795|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Lab|Laboratory or Test Result|History of Present Illness|1791,1795|false|false|false|C0344420||LBBB
Finding|Finding|History of Present Illness|1805,1814|false|false|false|C0442739||unchanged
Procedure|Diagnostic Procedure|History of Present Illness|1827,1830|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|History of Present Illness|1840,1845|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1846,1853|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|History of Present Illness|1846,1853|false|false|false|C1951340|Process Pharmacologic Substance|process
Finding|Functional Concept|History of Present Illness|1846,1853|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|History of Present Illness|1846,1853|false|false|false|C1522240|Process|process
Finding|Body Substance|History of Present Illness|1855,1862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|1855,1862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|1855,1862|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|History of Present Illness|1869,1876|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|History of Present Illness|1869,1876|false|false|false|C0004057|aspirin|aspirin
Drug|Organic Chemical|History of Present Illness|1920,1927|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|History of Present Illness|1920,1927|false|false|false|C0004057|aspirin|aspirin
Finding|Finding|History of Present Illness|1928,1935|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|History of Present Illness|1931,1935|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1931,1935|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1931,1935|false|false|false|C1553498|home health encounter|home
Anatomy|Body Location or Region|History of Present Illness|1985,1990|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1985,1990|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1985,1995|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1985,1995|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1991,1995|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1991,1995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1991,1995|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Health Care Activity|History of Present Illness|2030,2042|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2030,2042|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Functional Concept|History of Present Illness|2054,2062|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2054,2062|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2054,2062|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|2106,2113|false|false|false|C1706079||arrival
Finding|Functional Concept|History of Present Illness|2106,2113|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2121,2126|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|2128,2135|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2128,2135|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2128,2135|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2138,2145|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Finding|History of Present Illness|2227,2235|false|false|false|C2984078;C3889124|A little bit;Only a Little|a little
Finding|Finding|History of Present Illness|2227,2239|false|false|false|C2984078|A little bit|a little bit
Disorder|Disease or Syndrome|History of Present Illness|2229,2235|false|false|false|C0023882|Little's Disease|little
Finding|Finding|History of Present Illness|2229,2235|false|false|false|C3889124|Only a Little|little
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2236,2239|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Organic Chemical|History of Present Illness|2236,2239|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Drug|Pharmacologic Substance|History of Present Illness|2236,2239|false|false|false|C0045724;C0671702|2-(4-ethoxybenzyl)-1-diethylaminoethyl-5-isothiocyanatobenzimidazole;PTPNS1 protein, human|bit
Finding|Gene or Genome|History of Present Illness|2236,2239|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Intellectual Product|History of Present Illness|2236,2239|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Receptor|History of Present Illness|2236,2239|false|false|false|C0671702;C1705300;C1822726;C4321288|Breast-Impact of Treatment Scale;PTPNS1 protein, human;SIRPA gene;SIRPA wt Allele|bit
Finding|Finding|History of Present Illness|2274,2278|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|History of Present Illness|2291,2301|false|false|false|C5441521|Complaint (finding)|complaints
Disorder|Disease or Syndrome|Past Medical History|2329,2332|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Past Medical History|2335,2341|false|false|false|C0004096|Asthma|Asthma
Disorder|Disease or Syndrome|Past Medical History|2344,2358|false|false|false|C0012813|Diverticulitis|Diverticulitis
Finding|Gene or Genome|Past Medical History|2373,2376|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Anatomy|Body Location or Region|Past Medical History|2379,2384|false|false|false|C0524470|Right hip region structure|R hip
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2381,2384|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2381,2384|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Past Medical History|2381,2384|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Past Medical History|2381,2384|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Past Medical History|2381,2384|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2381,2384|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2381,2396|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Finding|Functional Concept|Past Medical History|2385,2396|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|2385,2396|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2385,2396|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Finding|Sign or Symptom|Past Medical History|2406,2416|false|false|false|C0239313|exercise induced|Exertional
Finding|Finding|Past Medical History|2417,2425|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Past Medical History|2417,2436|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|Past Medical History|2426,2431|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|2426,2431|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Past Medical History|2426,2436|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Past Medical History|2426,2436|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Past Medical History|2432,2436|false|true|false|C2598155||Pain
Finding|Functional Concept|Past Medical History|2432,2436|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Past Medical History|2432,2436|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Idea or Concept|Family Medical History|2475,2481|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|2488,2491|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Conceptual Entity|Family Medical History|2494,2500|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|2494,2500|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Conceptual Entity|Family Medical History|2511,2518|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2511,2518|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Conceptual Entity|Family Medical History|2526,2533|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|2526,2533|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Finding|Family Medical History|2544,2552|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|2544,2552|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|2544,2552|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|2561,2570|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Finding|Classification|Family Medical History|2624,2631|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|Family Medical History|2624,2631|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|Family Medical History|2648,2651|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|2648,2651|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|2648,2651|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|2648,2651|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|2648,2651|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|Family Medical History|2648,2651|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|Family Medical History|2653,2661|false|false|false|C1961028|Oriented to place|Oriented
Attribute|Clinical Attribute|Family Medical History|2666,2670|false|false|false|C2713234||Mood
Finding|Conceptual Entity|Family Medical History|2666,2670|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Finding|Family Medical History|2666,2670|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|Family Medical History|2666,2670|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|Mood
Finding|Mental Process|Family Medical History|2672,2678|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|Family Medical History|2672,2678|false|false|false|C2237113|assessment of affect|affect
Anatomy|Body Location or Region|Family Medical History|2695,2700|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2708,2714|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|Family Medical History|2708,2714|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|Family Medical History|2708,2714|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|Family Medical History|2715,2724|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2726,2737|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|Conjunctiva
Disorder|Disease or Syndrome|Family Medical History|2726,2737|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Disorder|Neoplastic Process|Family Medical History|2726,2737|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|Conjunctiva
Finding|Body Substance|Family Medical History|2726,2737|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Finding|Intellectual Product|Family Medical History|2726,2737|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|Conjunctiva
Procedure|Health Care Activity|Family Medical History|2726,2737|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|Conjunctiva
Finding|Finding|Family Medical History|2752,2758|true|false|false|C0241137|Pallor of skin|pallor
Finding|Sign or Symptom|Family Medical History|2763,2771|false|false|false|C0010520|Cyanosis|cyanosis
Anatomy|Body Space or Junction|Family Medical History|2779,2783|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Family Medical History|2779,2783|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Family Medical History|2779,2783|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Family Medical History|2779,2783|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2779,2790|false|false|false|C0026639|Oral mucous membrane structure|oral mucosa
Anatomy|Tissue|Family Medical History|2784,2790|false|false|false|C0026724|Mucous Membrane|mucosa
Finding|Intellectual Product|Family Medical History|2784,2790|false|false|false|C1561514||mucosa
Anatomy|Body Location or Region|Family Medical History|2810,2814|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|Family Medical History|2810,2814|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|Family Medical History|2810,2814|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|Family Medical History|2816,2822|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2825,2832|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|Family Medical History|2825,2832|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|Family Medical History|2866,2873|true|false|false|C0232269|Cardiac thrill (finding)|thrills
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2898,2903|false|false|false|C0024109|Lung|LUNGS
Anatomy|Body Location or Region|Family Medical History|2908,2913|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Family Medical History|2908,2913|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Location or Region|Family Medical History|2908,2918|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2908,2918|false|false|false|C0205076;C4266615|Chest wall structure;Chest>Chest wall|chest wall
Disorder|Anatomical Abnormality|Family Medical History|2908,2930|true|false|false|C3164427|Deformity of chest wall|chest wall deformities
Disorder|Congenital Abnormality|Family Medical History|2919,2930|true|false|false|C0000768|Congenital Abnormality|deformities
Disorder|Acquired Abnormality|Family Medical History|2932,2941|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Congenital Abnormality|Family Medical History|2932,2941|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Disease or Syndrome|Family Medical History|2932,2941|true|false|false|C0036439;C0559260;C0700208|Acquired scoliosis;Congenital scoliosis|scoliosis
Disorder|Acquired Abnormality|Family Medical History|2945,2953|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Anatomical Abnormality|Family Medical History|2945,2953|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Disorder|Congenital Abnormality|Family Medical History|2945,2953|true|false|false|C0022821;C0022822;C0265673|Acquired kyphosis;Congenital kyphosis;Kyphosis deformity of spine|kyphosis
Finding|Finding|Family Medical History|2945,2953|true|false|false|C2115817|kyphosis|kyphosis
Attribute|Clinical Attribute|Family Medical History|2955,2959|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|Family Medical History|2955,2959|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Finding|Functional Concept|Family Medical History|2966,2975|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|Family Medical History|2980,2996|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|Family Medical History|2980,3000|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2990,2996|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Family Medical History|2990,2996|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|Family Medical History|2997,3000|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Family Medical History|2997,3000|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Finding|Family Medical History|3002,3025|false|false|false|C0238844|Decreased breath sounds|decreased breath sounds
Finding|Body Substance|Family Medical History|3012,3018|false|false|false|C0225386|Breath|breath
Attribute|Clinical Attribute|Family Medical History|3012,3025|false|false|false|C0035234;C3484186|Respiratory Sounds|breath sounds
Phenomenon|Natural Phenomenon or Process|Family Medical History|3019,3025|false|false|false|C0037709||sounds
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3048,3051|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|Family Medical History|3048,3051|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Family Medical History|3048,3051|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Finding|Family Medical History|3056,3064|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Finding|Sign or Symptom|Family Medical History|3066,3073|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|Family Medical History|3077,3084|true|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|Family Medical History|3088,3095|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|Family Medical History|3088,3095|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|Family Medical History|3088,3095|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|Family Medical History|3097,3101|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Finding|Mental Process|Family Medical History|3112,3122|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Family Medical History|3112,3122|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3126,3137|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body System|Family Medical History|3151,3155|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|Family Medical History|3151,3155|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|Family Medical History|3151,3155|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|Family Medical History|3151,3155|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|Family Medical History|3151,3155|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Pathologic Function|Family Medical History|3160,3166|false|false|false|C0333138|Stasis|stasis
Disorder|Disease or Syndrome|Family Medical History|3160,3177|true|false|false|C0011620|Stasis dermatitis|stasis dermatitis
Disorder|Disease or Syndrome|Family Medical History|3167,3177|true|false|false|C0011603|Dermatitis|dermatitis
Finding|Pathologic Function|Family Medical History|3179,3185|true|false|false|C0041582|Ulcer|ulcers
Finding|Finding|Family Medical History|3187,3192|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Finding|Pathologic Function|Family Medical History|3187,3192|true|false|false|C0241158;C2004491|Cicatrix;Scar Tissue|scars
Disorder|Disease or Syndrome|Family Medical History|3197,3206|true|false|false|C0302314|Xanthoma|xanthomas
Drug|Food|Family Medical History|3210,3216|false|false|false|C5890763||PULSES
Finding|Physiologic Function|Family Medical History|3210,3216|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|Family Medical History|3210,3216|false|false|false|C0034107|Pulse taking|PULSES
Finding|Functional Concept|Family Medical History|3220,3225|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Finding|Functional Concept|Family Medical History|3242,3246|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Neoplastic Process|Family Medical History|3303,3306|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Family Medical History|3303,3306|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Procedure|Laboratory Procedure|Family Medical History|3330,3333|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Antibiotic|Family Medical History|3373,3378|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|Family Medical History|3373,3378|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|Family Medical History|3373,3378|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|Family Medical History|3383,3386|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|Family Medical History|3383,3386|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Anatomy|Cell|Family Medical History|3416,3419|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|3424,3427|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|3424,3427|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|3424,3427|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3433,3436|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|Family Medical History|3433,3436|false|false|false|C0019046|Hemoglobin|HGB
Finding|Gene or Genome|Family Medical History|3433,3436|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|Family Medical History|3433,3436|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|Family Medical History|3442,3445|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3442,3445|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|Family Medical History|3451,3454|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Family Medical History|3451,3454|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|3451,3454|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|3451,3454|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|3459,3462|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|3459,3462|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Family Medical History|3459,3462|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|3459,3462|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|3459,3462|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Family Medical History|3468,3472|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Drug|Biologically Active Substance|Family Medical History|3561,3568|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|Family Medical History|3561,3568|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|Family Medical History|3561,3568|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|Family Medical History|3561,3568|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|Family Medical History|3561,3568|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|Family Medical History|3572,3576|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|Family Medical History|3572,3576|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|Family Medical History|3572,3576|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|Family Medical History|3572,3576|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|Family Medical History|3593,3599|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|Family Medical History|3593,3599|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|Family Medical History|3593,3599|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|Family Medical History|3593,3599|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|Family Medical History|3593,3599|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|Family Medical History|3605,3614|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|Family Medical History|3605,3614|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|Family Medical History|3605,3614|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|Family Medical History|3605,3614|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|Family Medical History|3605,3614|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|Family Medical History|3605,3614|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|Family Medical History|3605,3614|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|Family Medical History|3619,3627|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|Family Medical History|3619,3627|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|Family Medical History|3619,3627|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|Family Medical History|3638,3641|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|Family Medical History|3638,3641|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|Family Medical History|3638,3641|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|Family Medical History|3638,3641|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|Family Medical History|3645,3650|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|Family Medical History|3645,3654|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|Family Medical History|3645,3654|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|Family Medical History|3645,3654|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3651,3654|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|Family Medical History|3651,3654|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|Family Medical History|3651,3654|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Drug|Biologically Active Substance|Family Medical History|3672,3679|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|Family Medical History|3672,3679|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|Family Medical History|3672,3679|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|Family Medical History|3672,3679|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|Family Medical History|3672,3679|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3704,3709|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|3704,3709|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|3704,3709|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|3704,3709|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|Family Medical History|3707,3711|false|false|false|C0602254|MB 3|MB-3
Drug|Amino Acid, Peptide, or Protein|Family Medical History|3743,3746|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|Family Medical History|3743,3746|false|false|false|C0010287|Creatine Kinase|CPK
Finding|Gene or Genome|Family Medical History|3743,3746|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|Family Medical History|3743,3746|false|false|false|C0201973|Creatine kinase measurement|CPK
Procedure|Diagnostic Procedure|Family Medical History|3753,3756|false|false|false|C0039985|Plain chest X-ray|CXR
Disorder|Disease or Syndrome|Family Medical History|3758,3767|false|false|false|C0034067|Pulmonary Emphysema|Emphysema
Finding|Pathologic Function|Family Medical History|3758,3767|false|false|false|C0013990|Pathological accumulation of air in tissues|Emphysema
Disorder|Disease or Syndrome|Family Medical History|3789,3798|true|false|false|C0032285|Pneumonia|pneumonia
Anatomy|Body Space or Junction|Family Medical History|3802,3805|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Family Medical History|3802,3805|true|false|false|C0018802|Congestive heart failure|CHF
Event|Activity|Hospital Course|3832,3842|false|false|false|C1516048|Assessed|ASSESSMENT
Finding|Intellectual Product|Hospital Course|3832,3842|false|false|false|C0679207|Knowledge acquisition using a method of assessment|ASSESSMENT
Procedure|Diagnostic Procedure|Hospital Course|3832,3842|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|ASSESSMENT
Procedure|Health Care Activity|Hospital Course|3832,3842|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|ASSESSMENT
Disorder|Disease or Syndrome|Hospital Course|3847,3851|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|PLAN
Finding|Functional Concept|Hospital Course|3847,3851|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Intellectual Product|Hospital Course|3847,3851|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Mental Process|Hospital Course|3847,3851|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|PLAN
Finding|Idea or Concept|Hospital Course|3870,3874|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|3870,3874|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Attribute|Clinical Attribute|Hospital Course|3901,3910|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|3901,3910|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|3901,3910|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|3901,3910|false|false|false|C0011900|Diagnosis|diagnosis
Disorder|Disease or Syndrome|Hospital Course|3914,3917|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3914,3917|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3914,3917|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|3914,3917|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3914,3917|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3914,3917|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3914,3917|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|3919,3922|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Hospital Course|3927,3933|false|false|false|C0004096|Asthma|asthma
Anatomy|Body Location or Region|Hospital Course|3978,3983|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|3978,3983|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|3978,3988|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|3978,3988|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|3984,3988|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|3984,3988|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|3984,3988|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|Hospital Course|4006,4015|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4006,4015|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4006,4015|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4006,4015|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|Hospital Course|4092,4099|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4092,4099|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4092,4099|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|4130,4134|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Hospital Course|4135,4140|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|4135,4140|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|Hospital Course|4142,4149|false|false|false|C0085624|Burning sensation|burning
Attribute|Clinical Attribute|Hospital Course|4175,4181|true|false|false|C2926611||angina
Finding|Finding|Hospital Course|4175,4181|true|false|false|C0002962;C2024883|Angina Pectoris|angina
Finding|Sign or Symptom|Hospital Course|4175,4181|true|false|false|C0002962;C2024883|Angina Pectoris|angina
Procedure|Health Care Activity|Hospital Course|4210,4222|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4210,4222|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Conceptual Entity|Hospital Course|4263,4274|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Mental Process|Hospital Course|4263,4274|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Finding|Social Behavior|Hospital Course|4263,4274|false|false|false|C0004083;C0699792;C1704770;C1704771|Association Class;Mental association;NCI Thesaurus Association;Relationship by association|association
Phenomenon|Phenomenon or Process|Hospital Course|4263,4274|false|false|false|C0596306|Chemical Association|association
Finding|Daily or Recreational Activity|Hospital Course|4280,4288|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4280,4288|false|false|false|C1522704|Exercise Pain Management|exercise
Attribute|Clinical Attribute|Hospital Course|4309,4317|false|false|false|C2926606||findings
Finding|Functional Concept|Hospital Course|4309,4317|false|false|false|C2607943|findings aspects|findings
Attribute|Clinical Attribute|Hospital Course|4333,4339|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|4333,4339|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|4333,4339|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|4333,4339|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|4333,4344|false|false|false|C0920208|Echocardiography, Stress|stress echo
Procedure|Health Care Activity|Hospital Course|4340,4344|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4340,4344|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Functional Concept|Hospital Course|4348,4357|false|false|false|C0205263|Induce (action)|inducible
Finding|Pathologic Function|Hospital Course|4358,4366|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4358,4366|false|false|false|C4321499|Ischemia Procedure|ischemia
Phenomenon|Natural Phenomenon or Process|Hospital Course|4394,4401|false|false|false|C1705970|Electrical Current|current
Finding|Functional Concept|Hospital Course|4402,4410|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|4402,4410|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|Hospital Course|4435,4445|false|false|false|C4722602|Underlying|underlying
Disorder|Disease or Syndrome|Hospital Course|4446,4449|false|true|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4446,4449|false|true|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|4446,4449|false|true|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|4446,4449|false|true|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|4446,4449|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|4446,4449|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4446,4449|false|true|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4456,4465|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|Hospital Course|4456,4465|false|false|false|C0041199|Troponin|troponins
Finding|Classification|Hospital Course|4471,4479|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|4471,4479|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|4471,4479|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|Hospital Course|4492,4500|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Health Care Activity|Hospital Course|4517,4526|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|4547,4552|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|Hospital Course|4547,4552|false|false|false|C0590690|Imdur|Imdur
Finding|Functional Concept|Hospital Course|4556,4570|false|false|false|C0332287|In addition to|in addition to
Finding|Functional Concept|Hospital Course|4559,4567|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Attribute|Clinical Attribute|Hospital Course|4576,4587|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|4576,4587|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|4576,4587|false|false|false|C4284232|Medications|medications
Finding|Body Substance|Hospital Course|4604,4613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|4604,4613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|4604,4613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|4604,4613|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|4651,4657|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Functional Concept|Hospital Course|4658,4665|false|true|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Hospital Course|4658,4665|false|true|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Hospital Course|4658,4665|false|true|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Hospital Course|4658,4665|false|true|false|C0199168|Medical service|medical
Event|Occupational Activity|Hospital Course|4666,4676|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|4666,4676|false|false|false|C0376636|Disease Management|management
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4699,4702|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Hospital Course|4699,4702|false|false|false|C2713669|SERPINA5 protein, human|PCI
Finding|Gene or Genome|Hospital Course|4699,4702|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Hospital Course|4699,4702|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4699,4702|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Event|Occupational Activity|Hospital Course|4754,4768|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4754,4768|false|false|false|C1533734|Administration (procedure)|administration
Drug|Organic Chemical|Hospital Course|4773,4778|false|false|false|C0590690|Imdur|IMDUR
Drug|Pharmacologic Substance|Hospital Course|4773,4778|false|false|false|C0590690|Imdur|IMDUR
Finding|Body Substance|Hospital Course|4794,4801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4794,4801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4794,4801|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|4820,4824|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|4851,4857|false|false|false|C4300351|Prior functioning.stairs|stairs
Finding|Sign or Symptom|Hospital Course|4878,4893|false|false|false|C0013404|Dyspnea|short of breath
Finding|Body Substance|Hospital Course|4887,4893|false|false|false|C0225386|Breath|breath
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4926,4933|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|4926,4933|false|false|false|C1314974|Cardiac attachment|cardiac
Anatomy|Body Location or Region|Hospital Course|4952,4957|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|4952,4957|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|4959,4963|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|4959,4963|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4959,4963|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4968,4972|false|false|false|C5552605|FACT Complex|fact
Drug|Biologically Active Substance|Hospital Course|4968,4972|false|false|false|C5552605|FACT Complex|fact
Finding|Gene or Genome|Hospital Course|4968,4972|false|false|false|C1420522;C5551287|SSRP1 wt Allele;SUPT16H gene|fact
Finding|Finding|Hospital Course|4999,5003|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Hospital Course|5020,5026|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Finding|Physiologic Function|Hospital Course|5020,5026|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|RHYTHM
Disorder|Disease or Syndrome|Hospital Course|5028,5032|false|false|false|C0023211|Left Bundle-Branch Block|LBBB
Lab|Laboratory or Test Result|Hospital Course|5028,5032|false|false|false|C0344420||LBBB
Finding|Intellectual Product|Hospital Course|5036,5039|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Hospital Course|5036,5039|false|false|false|C1623258|Electrocardiography|EKG
Finding|Body Substance|Hospital Course|5065,5072|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|5065,5072|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|5065,5072|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|5081,5084|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|5081,5084|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|5081,5094|false|false|false|C2585997|New diagnosis (finding)|new diagnosis
Procedure|Diagnostic Procedure|Hospital Course|5081,5094|false|false|false|C1882082|New Diagnosis Procedure|new diagnosis
Attribute|Clinical Attribute|Hospital Course|5085,5094|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|5085,5094|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|5085,5094|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|5085,5094|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Finding|Hospital Course|5098,5101|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Gene or Genome|Hospital Course|5098,5101|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Intellectual Product|Hospital Course|5098,5101|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Molecular Function|Hospital Course|5098,5101|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Procedure|Health Care Activity|Hospital Course|5110,5119|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|5142,5151|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|5142,5151|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|5181,5184|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Gene or Genome|Hospital Course|5181,5184|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Intellectual Product|Hospital Course|5181,5184|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Molecular Function|Hospital Course|5181,5184|false|false|false|C0221158;C1151970;C1412111;C1417038;C3714902;C5780814;C5890859|ACAT1 gene;ACAT1 wt Allele;MAT1A gene;MAT1A wt Allele;Multifocal atrial tachycardia;Multinational Association of Supportive Care in Cancer Antiemesis Tool;[acyl-carrier-protein] S-malonyltransferase activity|MAT
Finding|Gene or Genome|Hospital Course|5188,5192|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Intellectual Product|Hospital Course|5188,5192|false|false|false|C1420621;C1515258|TCAP gene;Telephone Number|tele
Finding|Finding|Hospital Course|5203,5215|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Disorder|Disease or Syndrome|Hospital Course|5232,5235|false|false|false|C0030587|Paroxysmal atrial tachycardia|PAT
Drug|Organic Chemical|Hospital Course|5232,5235|false|false|false|C2825250|Fenamole|PAT
Drug|Pharmacologic Substance|Hospital Course|5232,5235|false|false|false|C2825250|Fenamole|PAT
Finding|Molecular Function|Hospital Course|5232,5235|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|PAT
Procedure|Diagnostic Procedure|Hospital Course|5232,5235|false|false|false|C3897364|Thermoacoustic Computed Tomography|PAT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5244,5250|false|false|false|C0018787|Heart|Hearts
Drug|Hazardous or Poisonous Substance|Hospital Course|5251,5258|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|5251,5258|false|false|false|C0728873|Monitor brand of insecticide|monitor
Finding|Body Substance|Hospital Course|5284,5293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|5284,5293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|5284,5293|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|5284,5293|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|Hospital Course|5327,5335|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|5327,5335|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Finding|Hospital Course|5349,5364|false|false|false|C0080203|Tachyarrhythmia|tachyarrhythmia
Finding|Finding|Hospital Course|5413,5421|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|Inactive
Finding|Idea or Concept|Hospital Course|5413,5421|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|Inactive
Disorder|Disease or Syndrome|Hospital Course|5432,5444|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Idea or Concept|Hospital Course|5456,5460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5456,5460|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5456,5460|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|5461,5465|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Hospital Course|5461,5465|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Organic Chemical|Hospital Course|5470,5479|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|5470,5479|false|false|false|C0012373|diltiazem|diltiazem
Disorder|Disease or Syndrome|Hospital Course|5486,5492|false|false|false|C0004096|Asthma|Asthma
Finding|Idea or Concept|Hospital Course|5503,5507|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5503,5507|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5503,5507|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Hospital Course|5508,5519|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5508,5519|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|5508,5519|false|false|false|C4284232|Medications|medications
Disorder|Disease or Syndrome|Hospital Course|5527,5531|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Idea or Concept|Hospital Course|5543,5547|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5543,5547|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5543,5547|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|5548,5558|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|5548,5558|false|false|false|C0028978|omeprazole|omeprazole
Event|Occupational Activity|Hospital Course|5578,5582|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|Hospital Course|5578,5582|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Finding|Idea or Concept|Hospital Course|5625,5637|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Body Substance|Hospital Course|5649,5656|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|5649,5656|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|5649,5656|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|5672,5677|false|false|false|C0590690|Imdur|Imdur
Drug|Pharmacologic Substance|Hospital Course|5672,5677|false|false|false|C0590690|Imdur|Imdur
Attribute|Clinical Attribute|Hospital Course|5714,5725|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|5714,5725|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|5714,5725|false|false|false|C4284232|Medications|medications
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5767,5775|false|false|false|C0018787|Heart|coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5767,5782|false|false|false|C0205042|Coronary artery|coronary artery
Disorder|Disease or Syndrome|Hospital Course|5767,5790|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5776,5782|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|5776,5782|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Hospital Course|5776,5790|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Hospital Course|5783,5790|false|false|false|C0012634|Disease|disease
Finding|Conceptual Entity|Hospital Course|5804,5813|false|true|false|C4527371|Candidate|candidate
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5818,5821|false|false|false|C2713669|SERPINA5 protein, human|PCI
Drug|Biologically Active Substance|Hospital Course|5818,5821|false|false|false|C2713669|SERPINA5 protein, human|PCI
Finding|Gene or Genome|Hospital Course|5818,5821|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Finding|Intellectual Product|Hospital Course|5818,5821|false|false|false|C1418370;C1705930;C4049621|Peritoneal Cancer Index;SERPINA5 gene;SERPINA5 wt Allele|PCI
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5818,5821|false|false|false|C1514496;C1532338;C4724254|Percutaneous Coronary Intervention;Prophylactic Cranial Irradiation;photochemical internalization|PCI
Anatomy|Body Location or Region|Hospital Course|5856,5861|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|5856,5861|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|5856,5866|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|5856,5866|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|5862,5866|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|5862,5866|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5862,5866|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|5888,5893|false|false|false|C0441471|Event|event
Drug|Hazardous or Poisonous Substance|Hospital Course|5894,5901|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|5894,5901|false|false|false|C0728873|Monitor brand of insecticide|monitor
Finding|Idea or Concept|Hospital Course|5906,5916|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|5906,5916|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Disorder|Disease or Syndrome|Hospital Course|5920,5931|false|false|false|C0003811|Cardiac Arrhythmia|arrhythmias
Attribute|Clinical Attribute|Hospital Course|5934,5945|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|5934,5945|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|5934,5945|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|5934,5958|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|5949,5958|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Hospital Course|5961,5974|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5961,5974|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5961,5974|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Attribute|Clinical Attribute|Hospital Course|6000,6004|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6000,6004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6000,6004|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|6009,6018|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|6009,6018|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|6009,6026|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|6009,6026|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|6019,6026|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|6019,6026|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|6019,6026|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|Hospital Course|6048,6058|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6048,6058|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Sign or Symptom|Hospital Course|6094,6097|false|false|false|C0013404|Dyspnea|SOB
Finding|Sign or Symptom|Hospital Course|6101,6107|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|6112,6123|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6112,6123|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6112,6134|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|6124,6134|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|6124,6134|false|false|false|C0073992|salmeterol|salmeterol
Finding|Functional Concept|Hospital Course|6147,6157|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6147,6157|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6158,6161|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6158,6161|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6158,6161|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6158,6161|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|6165,6176|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6165,6176|false|false|false|C0082607|fluticasone|fluticasone
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6189,6194|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|6189,6194|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|6189,6194|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|6189,6194|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|6189,6194|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|6189,6194|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Intellectual Product|Hospital Course|6195,6199|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6195,6205|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6202,6205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6202,6205|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6209,6228|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|6209,6228|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Finding|Intellectual Product|Hospital Course|6235,6239|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6235,6245|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6242,6245|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6242,6245|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6250,6260|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|6250,6260|false|false|false|C0028978|omeprazole|omeprazole
Drug|Organic Chemical|Hospital Course|6276,6287|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|6276,6287|false|false|false|C0074554|simvastatin|simvastatin
Finding|Intellectual Product|Hospital Course|6294,6298|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6294,6304|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6301,6304|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6301,6304|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6309,6319|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Hospital Course|6309,6319|false|false|false|C0213771|tiotropium|tiotropium
Drug|Organic Chemical|Hospital Course|6309,6327|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Hospital Course|6309,6327|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Hospital Course|6320,6327|false|false|false|C0006222|Bromides|bromide
Procedure|Laboratory Procedure|Hospital Course|6320,6327|false|false|false|C0202341|Bromides measurement|bromide
Drug|Organic Chemical|Hospital Course|6344,6351|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|6344,6351|false|false|false|C0004057|aspirin|aspirin
Finding|Intellectual Product|Hospital Course|6358,6362|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|6358,6368|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|6365,6368|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6365,6368|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6373,6385|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|6373,6385|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|6373,6385|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Biomedical or Dental Material|Hospital Course|6388,6394|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|6404,6413|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|6404,6413|false|false|false|C0012373|diltiazem|diltiazem
Drug|Organic Chemical|Hospital Course|6404,6417|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Hospital Course|6404,6417|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Hospital Course|6414,6417|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|6414,6417|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|6414,6417|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|6414,6417|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Biomedical or Dental Material|Hospital Course|6425,6431|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|6442,6449|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|6442,6449|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6442,6449|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|6465,6474|false|false|false|C0595724|Singulair|singulair
Drug|Pharmacologic Substance|Hospital Course|6465,6474|false|false|false|C0595724|Singulair|singulair
Finding|Body Substance|Hospital Course|6488,6497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|6488,6497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|6488,6497|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|6488,6497|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|6488,6509|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|6498,6509|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|6498,6509|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|6498,6509|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|6514,6527|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|6514,6527|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|Hospital Course|6514,6527|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|6535,6541|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|6555,6561|false|false|false|C0039225|Tablet Dosage Form|Tablet
Attribute|Clinical Attribute|Hospital Course|6601,6605|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6601,6605|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6601,6605|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|6612,6621|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|6612,6621|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|6612,6629|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|6612,6629|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|6622,6629|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|6622,6629|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|6622,6629|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Disorder|Disease or Syndrome|Hospital Course|6647,6650|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|6647,6650|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Hospital Course|6651,6658|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Finding|Functional Concept|Hospital Course|6659,6666|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Hospital Course|6686,6696|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6686,6696|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Sign or Symptom|Hospital Course|6731,6734|false|false|false|C0013404|Dyspnea|sob
Finding|Sign or Symptom|Hospital Course|6737,6745|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|Hospital Course|6753,6764|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6753,6764|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6753,6775|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|6765,6775|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|6765,6775|false|false|false|C0073992|salmeterol|salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6792,6796|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|6792,6796|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|6802,6808|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6809,6812|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6809,6812|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|6809,6812|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|6809,6812|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6823,6827|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|6823,6827|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|6833,6839|false|false|false|C1550509|Participation Type - device|Device
Finding|Functional Concept|Hospital Course|6840,6850|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|6840,6850|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6851,6854|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6851,6854|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|6851,6854|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|6851,6854|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|6856,6863|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|6858,6863|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|6866,6869|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6866,6869|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|6877,6888|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|6877,6888|false|false|false|C0082607|fluticasone|fluticasone
Drug|Biomedical or Dental Material|Hospital Course|6906,6911|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|6906,6911|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|6906,6911|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Hospital Course|6906,6923|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Hospital Course|6913,6923|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Hospital Course|6913,6923|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Finding|Functional Concept|Hospital Course|6913,6923|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|Hospital Course|6938,6943|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Hospital Course|6938,6943|false|false|false|C2003858|Spray (action)|Spray
Finding|Functional Concept|Hospital Course|6938,6943|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6944,6949|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|6944,6949|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|6944,6949|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|6944,6949|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|6944,6949|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|6944,6949|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Drug|Organic Chemical|Hospital Course|6970,6989|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|6970,6989|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6998,7005|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|6998,7005|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|6998,7005|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7019,7026|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7019,7026|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7019,7026|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Intellectual Product|Hospital Course|7031,7035|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7031,7041|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7038,7041|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7038,7041|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7048,7058|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|7048,7058|false|false|false|C0028978|omeprazole|omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7065,7072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7065,7072|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7065,7072|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|7074,7081|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|7074,7089|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|Hospital Course|7082,7089|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7082,7089|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7082,7089|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7110,7117|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7110,7117|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7110,7117|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|7119,7126|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|7119,7134|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Finding|Functional Concept|Hospital Course|7127,7134|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7127,7134|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7127,7134|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|7164,7175|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Hospital Course|7164,7175|false|false|false|C0074554|simvastatin|simvastatin
Drug|Biomedical or Dental Material|Hospital Course|7182,7188|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7202,7208|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|7212,7216|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7212,7222|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7219,7222|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7219,7222|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7229,7239|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Hospital Course|7229,7239|false|false|false|C0213771|tiotropium|tiotropium
Drug|Organic Chemical|Hospital Course|7229,7247|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Hospital Course|7229,7247|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Hospital Course|7240,7247|false|false|false|C0006222|Bromides|bromide
Procedure|Laboratory Procedure|Hospital Course|7240,7247|false|false|false|C0202341|Bromides measurement|bromide
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7255,7262|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7255,7262|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7255,7262|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|7266,7276|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|7266,7276|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Functional Concept|Hospital Course|7277,7283|false|false|false|C1550509|Participation Type - device|Device
Disorder|Congenital Abnormality|Hospital Course|7298,7301|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Hospital Course|7298,7301|false|false|false|C0006935|capsule (pharmacologic)|Cap
Finding|Gene or Genome|Hospital Course|7298,7301|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7298,7301|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Finding|Functional Concept|Hospital Course|7302,7312|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|7302,7312|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Drug|Organic Chemical|Hospital Course|7333,7340|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|7333,7340|false|false|false|C0004057|aspirin|aspirin
Drug|Biomedical or Dental Material|Hospital Course|7347,7353|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7367,7373|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|7377,7381|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7377,7387|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7384,7387|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7384,7387|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7395,7407|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|7395,7407|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Hospital Course|7395,7407|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Hospital Course|7395,7418|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Hospital Course|7412,7418|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7432,7438|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|7464,7475|false|false|false|C0298130|montelukast|montelukast
Drug|Pharmacologic Substance|Hospital Course|7464,7475|false|false|false|C0298130|montelukast|montelukast
Drug|Biomedical or Dental Material|Hospital Course|7482,7488|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|7502,7508|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Intellectual Product|Hospital Course|7517,7521|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Idea or Concept|Hospital Course|7525,7528|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7525,7528|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|7550,7560|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Hospital Course|7550,7560|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|Hospital Course|7550,7572|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|Hospital Course|7550,7572|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Biomedical or Dental Material|Hospital Course|7579,7585|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|7596,7603|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7596,7603|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7596,7603|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Biomedical or Dental Material|Hospital Course|7624,7630|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|7641,7648|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7641,7648|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7641,7648|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|Hospital Course|7658,7662|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7658,7668|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7665,7668|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7665,7668|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|Hospital Course|7679,7685|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Functional Concept|Hospital Course|7696,7703|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7696,7703|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7696,7703|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|Hospital Course|7714,7721|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|7730,7739|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|7730,7739|false|false|false|C0012373|diltiazem|diltiazem
Drug|Organic Chemical|Hospital Course|7730,7743|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Hospital Course|7730,7743|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Hospital Course|7740,7743|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Hospital Course|7740,7743|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Hospital Course|7740,7743|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Hospital Course|7740,7743|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7751,7758|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7751,7758|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7751,7758|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|7766,7773|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7766,7773|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7766,7773|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7794,7801|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7794,7801|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7794,7801|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|7809,7816|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7809,7816|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7809,7816|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Intellectual Product|Hospital Course|7826,7830|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Hospital Course|7826,7836|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Hospital Course|7833,7836|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|7833,7836|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7847,7854|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|7847,7854|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|7847,7854|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Hospital Course|7862,7869|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|7862,7869|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7862,7869|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|Hospital Course|7880,7887|false|false|false|C0807726|refill|Refills
Finding|Body Substance|Hospital Course|7895,7904|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7895,7904|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7895,7904|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7895,7904|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|7895,7916|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|7895,7916|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|7905,7916|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|7905,7916|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|7918,7922|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|7918,7922|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|7918,7922|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|Hospital Course|7925,7934|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|7925,7934|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|7925,7934|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|7925,7934|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|7925,7944|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|7935,7944|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|7935,7944|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|7935,7944|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|7935,7944|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Hospital Course|7958,7966|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|Hospital Course|7958,7977|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|Hospital Course|7967,7972|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|7967,7972|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|7967,7977|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|7967,7977|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|7973,7977|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7973,7977|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7973,7977|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Neoplastic Process|Hospital Course|7979,7988|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|7979,7988|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|Hospital Course|7994,8006|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Hospital Course|8010,8016|false|false|false|C0004096|Asthma|Asthma
Disorder|Disease or Syndrome|Hospital Course|8020,8034|false|false|false|C0012813|Diverticulitis|Diverticulitis
Finding|Mental Process|Discharge Condition|8059,8065|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8059,8072|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8059,8072|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8066,8072|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8066,8072|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|8074,8079|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|8084,8092|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|8094,8116|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8094,8116|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|8103,8116|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8103,8116|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8118,8123|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8118,8123|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8118,8123|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|8118,8123|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8118,8123|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8118,8123|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8128,8139|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8141,8149|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8141,8149|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8141,8149|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8150,8156|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8150,8156|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|8158,8168|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8158,8168|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8158,8168|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8158,8168|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|8171,8182|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8171,8182|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Instructions|8236,8244|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|Discharge Instructions|8249,8257|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|Discharge Instructions|8249,8268|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|Discharge Instructions|8258,8263|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|8258,8263|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|8258,8268|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|8258,8268|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|8264,8268|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|8264,8268|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8264,8268|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Diagnostic Procedure|Discharge Instructions|8293,8302|false|false|false|C0039451|Telemetry|telemetry
Finding|Intellectual Product|Discharge Instructions|8309,8312|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Discharge Instructions|8309,8312|false|false|false|C1623258|Electrocardiography|EKG
Finding|Finding|Discharge Instructions|8317,8326|false|false|false|C0442739||unchanged
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8334,8341|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Discharge Instructions|8334,8341|false|false|false|C1314974|Cardiac attachment|cardiac
Attribute|Clinical Attribute|Discharge Instructions|8334,8349|false|false|false|C2926589||cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|8334,8349|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Drug|Enzyme|Discharge Instructions|8334,8349|false|false|false|C0443763|Cardiac enzymes|cardiac enzymes
Procedure|Laboratory Procedure|Discharge Instructions|8334,8349|false|false|false|C0201934|Cardiac enzymes/isoenzymes measurement|cardiac enzymes
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|8342,8349|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Enzyme|Discharge Instructions|8342,8349|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Drug|Pharmacologic Substance|Discharge Instructions|8342,8349|false|false|false|C0014442;C3540017;C3540048;C3540772;C3540790;C3541394;C3542456|ENZYMES FOR TREATMENT OF WOUNDS AND ULCERS;Enzymes;Enzymes FOR DISORDERS OF THE MUSCULO-SKELETAL SYSTEM;Enzymes for ALIMENTARY TRACT AND METABOLISM;Enzymes, antithrombotic;Enzymes, hematological;Enzymes, peripheral vasodilators|enzymes
Finding|Functional Concept|Discharge Instructions|8342,8349|false|false|false|C0014445|enzymology|enzymes
Finding|Idea or Concept|Discharge Instructions|8371,8379|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|8371,8383|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence for
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8384,8389|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8384,8389|true|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8384,8389|true|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|Discharge Instructions|8390,8396|true|false|false|C0010957|Tissue damage|damage
Finding|Functional Concept|Discharge Instructions|8390,8396|true|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Finding|Gene or Genome|Discharge Instructions|8390,8396|true|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8401,8406|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8401,8406|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8401,8406|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|8401,8413|false|false|false|C0027051|Myocardial Infarction|heart attack
Finding|Finding|Discharge Instructions|8407,8413|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Finding|Social Behavior|Discharge Instructions|8407,8413|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|attack
Drug|Element, Ion, or Isotope|Discharge Instructions|8452,8459|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Inorganic Chemical|Discharge Instructions|8452,8459|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|Discharge Instructions|8452,8459|false|false|false|C0028125;C0699857;C3848573|Nitrate;Nitrates;nitrate ion|nitrate
Drug|Pharmacologic Substance|Discharge Instructions|8461,8471|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|8461,8471|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Anatomy|Body Location or Region|Discharge Instructions|8488,8493|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|8488,8493|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|8488,8498|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|8488,8498|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|8494,8498|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|8494,8498|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8494,8498|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8494,8507|false|false|false|C0030193|Pain|pain symptoms
Finding|Functional Concept|Discharge Instructions|8499,8507|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|8499,8507|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|Discharge Instructions|8533,8542|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Discharge Instructions|8533,8542|false|false|false|C0012373|diltiazem|diltiazem
Finding|Idea or Concept|Discharge Instructions|8547,8553|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|Discharge Instructions|8554,8559|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|8554,8559|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|8554,8568|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|8554,8568|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|8554,8568|false|false|false|C0005824|Blood pressure determination|blood pressure
Finding|Finding|Discharge Instructions|8560,8568|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|8560,8568|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|8560,8568|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|8560,8568|false|false|false|C0033095||pressure
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8573,8578|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8573,8578|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8573,8578|false|false|false|C0795691|HEART PROBLEM|heart
Event|Activity|Discharge Instructions|8580,8584|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Discharge Instructions|8580,8584|false|false|false|C1549480|Amount type - Rate|rate
Finding|Functional Concept|Discharge Instructions|8580,8592|false|false|false|C0489879|rate control|rate control
Drug|Organic Chemical|Discharge Instructions|8585,8592|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Discharge Instructions|8585,8592|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Discharge Instructions|8585,8592|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|Discharge Instructions|8585,8592|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Discharge Instructions|8585,8592|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Discharge Instructions|8585,8592|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Procedure|Diagnostic Procedure|Discharge Instructions|8639,8653|false|false|false|C0013801|Holter Electrocardiography|holter monitor
Drug|Hazardous or Poisonous Substance|Discharge Instructions|8646,8653|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Discharge Instructions|8646,8653|false|false|false|C0728873|Monitor brand of insecticide|monitor
Finding|Idea or Concept|Discharge Instructions|8664,8670|false|false|false|C1550462|Observation Interpretation - better|better
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8684,8689|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8684,8689|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8684,8689|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|Discharge Instructions|8684,8696|false|false|false|C0232187|Cardiac rhythm type|heart rhythm
Finding|Finding|Discharge Instructions|8690,8696|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Discharge Instructions|8690,8696|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|Discharge Instructions|8702,8706|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|8702,8706|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|8702,8706|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body System|Discharge Instructions|8770,8780|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Activity|Discharge Instructions|8781,8792|false|false|false|C0003629|Appointments|appointment
Drug|Pharmacologic Substance|Discharge Instructions|8796,8806|false|false|false|C0013227|Pharmaceutical Preparations|MEDICATION
Finding|Intellectual Product|Discharge Instructions|8796,8806|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|MEDICATION
Finding|Functional Concept|Discharge Instructions|8807,8814|false|false|false|C0392747|Changing|CHANGES
Drug|Food|Discharge Instructions|8818,8823|false|false|false|C0452588|Start brand of breakfast cereal|START
Finding|Intellectual Product|Discharge Instructions|8818,8823|false|false|false|C1552850|start - HtmlLinkType|START
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8818,8823|false|false|false|C5447432|Collagen Tile Brachytherapy|START
Finding|Functional Concept|Discharge Instructions|8844,8852|false|false|false|C0442805|Increase|INCREASE
Drug|Organic Chemical|Discharge Instructions|8853,8862|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Discharge Instructions|8853,8862|false|false|false|C0012373|diltiazem|diltiazem
Attribute|Clinical Attribute|Discharge Instructions|8908,8919|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|8908,8919|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|8908,8919|false|false|false|C4284232|Medications|medications
Finding|Functional Concept|Discharge Instructions|8949,8956|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|8949,8956|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|8949,8956|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|8949,8956|false|false|false|C0199168|Medical service|medical
Finding|Intellectual Product|Discharge Instructions|8957,8966|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Discharge Instructions|8957,8966|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Anatomy|Body Location or Region|Discharge Instructions|8981,8986|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Discharge Instructions|8981,8986|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Discharge Instructions|8981,8991|false|true|false|C2926613||chest pain
Finding|Sign or Symptom|Discharge Instructions|8981,8991|false|true|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Discharge Instructions|8987,8991|false|true|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|8987,8991|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|8987,8991|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|Discharge Instructions|8994,9013|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|8994,9013|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|9007,9013|false|false|false|C0225386|Breath|breath
Finding|Functional Concept|Discharge Instructions|9028,9036|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|9028,9036|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Procedure|Health Care Activity|Discharge Instructions|9040,9048|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9049,9061|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|9049,9061|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

