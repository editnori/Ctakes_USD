 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
<EOL>|206,207
<EOL>|208,209
Chest|226,231
pain|232,236
<EOL>|236,237
<EOL>|238,239
Major|239,244
Surgical|245,253
or|254,256
Invasive|257,265
Procedure|266,275
:|275,276
<EOL>|276,277
None|277,281
<EOL>|281,282
<EOL>|283,284
Ms.|312,315
_|316,317
_|317,318
_|318,319
is|320,322
a|323,324
_|325,326
_|326,327
_|327,328
year|329,333
old|334,337
woman|338,343
with|344,348
extensive|349,358
cardiac|359,366
history|367,374
<EOL>|375,376
including|376,385
multivessel|386,397
vessel|398,404
CAD|405,408
S|409,410
/|410,411
P|411,412
stenting|413,421
of|422,424
the|425,428
LAD|429,432
with|433,437
<EOL>|438,439
in|439,441
-|441,442
stent|442,447
restenosis|448,458
and|459,462
stenting|463,471
of|472,474
the|475,478
CX|479,481
,|481,482
S|483,484
/|484,485
P|485,486
CABG|487,491
in|492,494
_|495,496
_|496,497
_|497,498
with|499,503
known|504,509
occluded|510,518
SVG|519,522
-|522,523
D1|523,525
with|526,530
patent|531,537
LIMA|538,542
-|542,543
LAD|543,546
and|547,550
SVG|551,554
-|554,555
OM|555,557
<EOL>|558,559
in|559,561
_|562,563
_|563,564
_|564,565
,|565,566
poorly|567,573
controlled|574,584
type|585,589
2|590,591
diabetes|592,600
mellitus|601,609
,|609,610
<EOL>|611,612
hypertension|612,624
,|624,625
COPD|626,630
,|630,631
GERD|632,636
,|636,637
now|638,641
presenting|642,652
with|653,657
new|658,661
chest|662,667
pain|668,672
.|672,673
<EOL>|673,674
At|676,678
5|679,680
pm|681,683
on|684,686
the|687,690
day|691,694
of|695,697
presentation|698,710
,|710,711
she|712,715
was|716,719
resting|720,727
at|728,730
home|731,735
<EOL>|736,737
when|737,741
she|742,745
had|746,749
onset|750,755
of|756,758
severe|759,765
stabbing|766,774
pain|775,779
left|780,784
of|785,787
the|788,791
sternum|792,799
.|799,800
<EOL>|801,802
This|802,806
pain|807,811
radiated|812,820
across|821,827
her|828,831
chest|832,837
but|838,841
not|842,845
to|846,848
the|849,852
arm|853,856
or|857,859
jaw|860,863
.|863,864
<EOL>|865,866
She|866,869
took|870,874
1|875,876
nitroglycerin|877,890
,|890,891
which|892,897
improved|898,906
her|907,910
pain|911,915
slightly|916,924
.|924,925
She|926,929
<EOL>|930,931
reports|931,938
that|939,943
the|944,947
pain|948,952
came|953,957
in|958,960
waves|961,966
lasting|967,974
5|975,976
minutes|977,984
.|984,985
She|986,989
also|990,994
<EOL>|995,996
endorsed|996,1004
left|1005,1009
chest|1010,1015
wall|1016,1020
tenderness|1021,1031
.|1031,1032
She|1033,1036
did|1037,1040
not|1041,1044
remember|1045,1053
when|1054,1058
<EOL>|1059,1060
she|1060,1063
last|1064,1068
had|1069,1072
chest|1073,1078
pain|1079,1083
prior|1084,1089
to|1090,1092
this|1093,1097
.|1097,1098
The|1099,1102
pain|1103,1107
was|1108,1111
not|1112,1115
clearly|1116,1123
<EOL>|1124,1125
exertional|1125,1135
.|1135,1136
The|1137,1140
sharp|1141,1146
pains|1147,1152
occurred|1153,1161
when|1162,1166
she|1167,1170
was|1171,1174
lying|1175,1180
down|1181,1185
.|1185,1186
<EOL>|1187,1188
She|1188,1191
says|1192,1196
the|1197,1200
area|1201,1205
is|1206,1208
very|1209,1213
tender|1214,1220
.|1220,1221
Lying|1222,1227
on|1228,1230
the|1231,1234
left|1235,1239
side|1240,1244
causes|1245,1251
<EOL>|1252,1253
pain|1253,1257
.|1257,1258
She|1259,1262
did|1263,1266
have|1267,1271
nausea|1272,1278
the|1279,1282
past|1283,1287
3|1288,1289
mornings|1290,1298
which|1299,1304
resolved|1305,1313
.|1313,1314
<EOL>|1315,1316
She|1316,1319
denied|1320,1326
vomiting|1327,1335
,|1335,1336
diaphoresis|1337,1348
,|1348,1349
fevers|1350,1356
or|1357,1359
chills|1360,1366
.|1366,1367
She|1368,1371
had|1372,1375
an|1376,1378
<EOL>|1379,1380
episode|1380,1387
of|1388,1390
diarrhea|1391,1399
yesterday|1400,1409
,|1409,1410
but|1411,1414
no|1415,1417
abdominal|1418,1427
pain|1428,1432
.|1432,1433
She|1434,1437
<EOL>|1438,1439
already|1439,1446
took|1447,1451
a|1452,1453
full|1454,1458
dose|1459,1463
aspirin|1464,1471
on|1472,1474
the|1475,1478
day|1479,1482
of|1483,1485
presentation|1486,1498
.|1498,1499
<EOL>|1501,1502
In|1504,1506
the|1507,1510
ED|1511,1513
,|1513,1514
initial|1515,1522
vitals|1523,1529
were|1530,1534
:|1534,1535
T|1536,1537
98.0|1538,1542
,|1542,1543
HR|1544,1546
88|1547,1549
,|1549,1550
BP|1551,1553
127|1554,1557
/|1557,1558
65|1558,1560
,|1560,1561
RR|1562,1564
<EOL>|1565,1566
16|1566,1568
,|1568,1569
SaO2|1570,1574
100|1575,1578
%|1578,1579
on|1580,1582
RA|1583,1585
.|1585,1586
FSBG|1587,1591
302|1592,1595
-|1595,1596
>|1596,1597
94|1597,1599
.|1599,1600
Labs|1601,1605
notable|1606,1613
for|1614,1617
Troponin|1618,1626
-|1626,1627
T|1627,1628
<|1629,1630
<EOL>|1631,1632
0.01|1632,1636
,|1636,1637
CK|1638,1640
-|1640,1641
MB|1641,1643
<|1644,1645
1|1646,1647
,|1647,1648
D|1649,1650
-|1650,1651
Dimer|1651,1656
268|1657,1660
,|1660,1661
Cr|1662,1664
1.2|1665,1668
,|1668,1669
Mg|1670,1672
1.4|1673,1676
.|1676,1677
Normal|1678,1684
LFTs|1685,1689
;|1689,1690
CBC|1691,1694
,|1694,1695
<EOL>|1696,1697
Chem|1697,1701
7|1702,1703
,|1703,1704
coags|1705,1710
WNL|1711,1714
.|1714,1715
CXR|1716,1719
showed|1720,1726
no|1727,1729
acute|1730,1735
cardiopulmonary|1736,1751
<EOL>|1752,1753
abnormality|1753,1764
.|1764,1765
Bedside|1766,1773
echocardiogram|1774,1788
showed|1789,1795
no|1796,1798
substantial|1799,1810
<EOL>|1811,1812
pericardial|1812,1823
effusion|1824,1832
or|1833,1835
tamponade|1836,1845
.|1845,1846
Patient|1847,1854
was|1855,1858
given|1859,1864
fluticasone|1865,1876
<EOL>|1877,1878
propionate|1878,1888
inhaled|1889,1896
,|1896,1897
OxyCODONE|1898,1907
-|1907,1908
-|1908,1909
Acetaminophen|1909,1922
(|1923,1924
5mg|1924,1927
-|1927,1928
325mg|1928,1933
)|1933,1934
,|1934,1935
<EOL>|1936,1937
Magnesium|1937,1946
Sulfate|1947,1954
2|1955,1956
gm|1957,1959
IV|1960,1962
.|1962,1963
<EOL>|1964,1965
<EOL>|1965,1966
On|1966,1968
arrival|1969,1976
to|1977,1979
the|1980,1983
cardiology|1984,1994
ward|1995,1999
,|1999,2000
the|2001,2004
patient|2005,2012
reported|2013,2021
that|2022,2026
her|2027,2030
<EOL>|2031,2032
pain|2032,2036
was|2037,2040
still|2041,2046
there|2047,2052
but|2053,2056
it|2057,2059
felt|2060,2064
"|2065,2066
slow|2066,2070
"|2070,2071
_|2073,2074
_|2074,2075
_|2075,2076
but|2077,2080
at|2081,2083
its|2084,2087
worse|2088,2093
<EOL>|2094,2095
was|2095,2098
_|2099,2100
_|2100,2101
_|2101,2102
.|2102,2103
The|2104,2107
area|2108,2112
was|2113,2116
tender|2117,2123
.|2123,2124
She|2125,2128
had|2129,2132
no|2133,2135
breathing|2136,2145
complaints|2146,2156
.|2156,2157
<EOL>|2158,2159
She|2159,2162
felt|2163,2167
a|2168,2169
little|2170,2176
congested|2177,2186
this|2187,2191
evening|2192,2199
when|2200,2204
the|2205,2208
pain|2209,2213
started|2214,2221
.|2221,2222
<EOL>|2222,2223
<EOL>|2224,2225
-|2247,2248
COPD|2248,2252
<EOL>|2252,2253
-|2253,2254
CAD|2254,2257
s|2258,2259
/|2259,2260
p|2260,2261
CABG|2262,2266
and|2267,2270
stenting|2271,2279
,|2279,2280
as|2281,2283
above|2284,2289
<EOL>|2289,2290
-|2290,2291
Depression|2291,2301
<EOL>|2303,2304
-|2304,2305
DM|2305,2307
<EOL>|2309,2310
-|2310,2311
GERD|2311,2315
<EOL>|2317,2318
-|2318,2319
Hypertension|2319,2331
<EOL>|2331,2332
-|2332,2333
Migraines|2333,2342
<EOL>|2342,2343
-|2343,2344
Chronic|2344,2351
shoulder|2352,2360
pain|2361,2365
on|2366,2368
narcotics|2369,2378
<EOL>|2378,2379
-|2379,2380
OSA|2380,2383
<EOL>|2383,2384
-|2384,2385
Peripheral|2385,2395
neuropathy|2396,2406
<EOL>|2406,2407
-|2407,2408
Restless|2408,2416
leg|2417,2420
<EOL>|2420,2421
<EOL>|2422,2423
:|2437,2438
<EOL>|2438,2439
_|2439,2440
_|2440,2441
_|2441,2442
<EOL>|2442,2443
:|2457,2458
<EOL>|2458,2459
Patient|2459,2466
was|2467,2470
ward|2471,2475
of|2476,2478
the|2479,2482
_|2483,2484
_|2484,2485
_|2485,2486
,|2486,2487
does|2488,2492
n't|2492,2495
know|2496,2500
full|2501,2505
details|2506,2513
of|2514,2516
<EOL>|2517,2518
.|2532,2533
Mother|2534,2540
with|2541,2545
possible|2546,2554
alcohol|2555,2562
abuse|2563,2568
.|2568,2569
Father|2570,2576
<EOL>|2577,2578
deceased|2578,2586
at|2587,2589
_|2590,2591
_|2591,2592
_|2592,2593
from|2594,2598
Hodgkin|2599,2606
's|2606,2608
Disease|2609,2616
per|2617,2620
old|2621,2624
records|2625,2632
.|2632,2633
<EOL>|2633,2634
<EOL>|2635,2636
On|2651,2653
admission|2654,2663
<EOL>|2663,2664
General|2664,2671
:|2671,2672
Obese|2673,2678
middle|2679,2685
aged|2686,2690
_|2691,2692
_|2692,2693
_|2693,2694
woman|2695,2700
,|2700,2701
alert|2702,2707
,|2707,2708
oriented|2709,2717
,|2717,2718
in|2719,2721
no|2722,2724
<EOL>|2725,2726
acute|2726,2731
distress|2732,2740
<EOL>|2740,2741
Vital|2741,2746
Signs|2747,2752
:|2752,2753
T|2754,2755
98.7|2756,2760
,|2760,2761
BP|2762,2764
98|2765,2767
/|2767,2768
65|2768,2770
,|2770,2771
HR|2772,2774
79|2775,2777
,|2777,2778
RR|2779,2781
18|2782,2784
,|2784,2785
SaO2|2786,2790
95|2791,2793
%|2793,2794
on|2795,2797
RA|2798,2800
<EOL>|2800,2801
Weight|2801,2807
:|2807,2808
89|2809,2811
kg|2812,2814
<EOL>|2814,2815
HEENT|2815,2820
:|2820,2821
Sclera|2822,2828
anicteric|2829,2838
,|2838,2839
mucous|2840,2846
membranes|2847,2856
moist|2857,2862
,|2862,2863
oropharynx|2864,2874
<EOL>|2875,2876
clear|2876,2881
<EOL>|2881,2882
NECK|2882,2886
:|2886,2887
difficult|2888,2897
to|2898,2900
appreciate|2901,2911
JVP|2912,2915
<EOL>|2915,2916
CV|2916,2918
:|2918,2919
Regular|2920,2927
rate|2928,2932
and|2933,2936
rhythm|2937,2943
,|2943,2944
normal|2945,2951
S1|2952,2954
+|2955,2956
S2|2957,2959
;|2959,2960
no|2961,2963
murmurs|2964,2971
,|2971,2972
rubs|2973,2977
,|2977,2978
<EOL>|2979,2980
gallops|2980,2987
<EOL>|2987,2988
Chest|2988,2993
:|2993,2994
Tenderness|2995,3005
to|3006,3008
palpation|3009,3018
of|3019,3021
the|3022,3025
left|3026,3030
anterior|3031,3039
chest|3040,3045
wall|3046,3050
<EOL>|3050,3051
Lungs|3051,3056
:|3056,3057
Clear|3058,3063
to|3064,3066
auscultation|3067,3079
bilaterally|3080,3091
-|3091,3092
-|3092,3093
no|3093,3095
wheezes|3096,3103
,|3103,3104
rales|3105,3110
,|3110,3111
<EOL>|3112,3113
rhonchi|3113,3120
<EOL>|3120,3121
Abdomen|3121,3128
:|3128,3129
Soft|3130,3134
,|3134,3135
non-tender|3136,3146
,|3146,3147
non-distended|3148,3161
,|3161,3162
obese|3163,3168
<EOL>|3168,3169
GU|3169,3171
:|3171,3172
No|3173,3175
Foley|3176,3181
<EOL>|3181,3182
Ext|3182,3185
:|3185,3186
Warm|3187,3191
,|3191,3192
well|3193,3197
perfused|3198,3206
;|3206,3207
no|3208,3210
clubbing|3211,3219
,|3219,3220
cyanosis|3221,3229
or|3230,3232
edema|3233,3238
<EOL>|3238,3239
<EOL>|3239,3240
Exam|3240,3244
unchanged|3245,3254
at|3255,3257
discharge|3258,3267
,|3267,3268
left|3269,3273
chest|3274,3279
wall|3280,3284
tender|3285,3291
with|3292,3296
<EOL>|3297,3298
palpation|3298,3307
with|3308,3312
pain|3313,3317
after|3318,3323
change|3324,3330
in|3331,3333
position|3334,3342
<EOL>|3342,3343
<EOL>|3344,3345
Pertinent|3345,3354
Results|3355,3362
:|3362,3363
<EOL>|3363,3364
_|3364,3365
_|3365,3366
_|3366,3367
10|3368,3370
:|3370,3371
31PM|3371,3375
BLOOD|3376,3381
WBC|3382,3385
-|3385,3386
9.4|3386,3389
RBC|3390,3393
-|3393,3394
3|3394,3395
.|3395,3396
51|3396,3398
*|3398,3399
Hgb|3400,3403
-|3403,3404
12.0|3404,3408
Hct|3409,3412
-|3412,3413
34.3|3413,3417
<EOL>|3418,3419
MCV|3419,3422
-|3422,3423
98|3423,3425
MCH|3426,3429
-|3429,3430
34|3430,3432
.|3432,3433
2|3433,3434
*|3434,3435
MCHC|3436,3440
-|3440,3441
35.0|3441,3445
RDW|3446,3449
-|3449,3450
11.8|3450,3454
RDWSD|3455,3460
-|3460,3461
42.3|3461,3465
Plt|3466,3469
_|3470,3471
_|3471,3472
_|3472,3473
<EOL>|3473,3474
<EOL>|3474,3475
_|3475,3476
_|3476,3477
_|3477,3478
10|3479,3481
:|3481,3482
31PM|3482,3486
BLOOD|3487,3492
Glucose|3493,3500
-|3500,3501
105|3501,3504
*|3504,3505
UreaN|3506,3511
-|3511,3512
21|3512,3514
*|3514,3515
Creat|3516,3521
-|3521,3522
1|3522,3523
.|3523,3524
2|3524,3525
*|3525,3526
Na|3527,3529
-|3529,3530
137|3530,3533
<EOL>|3534,3535
K|3535,3536
-|3536,3537
3.4|3537,3540
Cl|3541,3543
-|3543,3544
97|3544,3546
HCO3|3547,3551
-|3551,3552
24|3552,3554
AnGap|3555,3560
-|3560,3561
19|3561,3563
<EOL>|3563,3564
_|3564,3565
_|3565,3566
_|3566,3567
10|3568,3570
:|3570,3571
31PM|3571,3575
BLOOD|3576,3581
ALT|3582,3585
-|3585,3586
15|3586,3588
AST|3589,3592
-|3592,3593
16|3593,3595
CK|3596,3598
(|3598,3599
CPK|3599,3602
)|3602,3603
-|3603,3604
39|3604,3606
AlkPhos|3607,3614
-|3614,3615
53|3615,3617
<EOL>|3618,3619
TotBili|3619,3626
-|3626,3627
0.3|3627,3630
<EOL>|3630,3631
_|3631,3632
_|3632,3633
_|3633,3634
10|3635,3637
:|3637,3638
31PM|3638,3642
BLOOD|3643,3648
Albumin|3649,3656
-|3656,3657
3.9|3657,3660
Calcium|3661,3668
-|3668,3669
9.1|3669,3672
Phos|3673,3677
-|3677,3678
4.4|3678,3681
Mg|3682,3684
-|3684,3685
1.4|3685,3688
*|3688,3689
<EOL>|3689,3690
<EOL>|3690,3691
_|3691,3692
_|3692,3693
_|3693,3694
10|3695,3697
:|3697,3698
57PM|3698,3702
BLOOD|3703,3708
D|3709,3710
-|3710,3711
Dimer|3711,3716
-|3716,3717
268|3717,3720
<EOL>|3720,3721
_|3721,3722
_|3722,3723
_|3723,3724
10|3725,3727
:|3727,3728
31PM|3728,3732
BLOOD|3733,3738
CK|3739,3741
-|3741,3742
MB|3742,3744
-|3744,3745
1|3745,3746
cTropnT|3748,3755
-|3755,3756
<|3756,3757
0|3757,3758
.|3758,3759
01|3759,3761
<EOL>|3761,3762
_|3762,3763
_|3763,3764
_|3764,3765
06|3766,3768
:|3768,3769
00AM|3769,3773
BLOOD|3774,3779
CK|3780,3782
-|3782,3783
MB|3783,3785
-|3785,3786
<|3786,3787
1|3787,3788
cTropnT|3789,3796
-|3796,3797
<|3797,3798
0|3798,3799
.|3799,3800
01|3800,3802
<EOL>|3802,3803
<EOL>|3803,3804
_|3804,3805
_|3805,3806
_|3806,3807
06|3808,3810
:|3810,3811
00AM|3811,3815
BLOOD|3816,3821
WBC|3822,3825
-|3825,3826
9.3|3826,3829
RBC|3830,3833
-|3833,3834
3|3834,3835
.|3835,3836
44|3836,3838
*|3838,3839
Hgb|3840,3843
-|3843,3844
11.8|3844,3848
Hct|3849,3852
-|3852,3853
33|3853,3855
.|3855,3856
1|3856,3857
*|3857,3858
<EOL>|3859,3860
MCV|3860,3863
-|3863,3864
96|3864,3866
MCH|3867,3870
-|3870,3871
34|3871,3873
.|3873,3874
3|3874,3875
*|3875,3876
MCHC|3877,3881
-|3881,3882
35.6|3882,3886
RDW|3887,3890
-|3890,3891
11.9|3891,3895
RDWSD|3896,3901
-|3901,3902
41.3|3902,3906
Plt|3907,3910
_|3911,3912
_|3912,3913
_|3913,3914
<EOL>|3914,3915
_|3915,3916
_|3916,3917
_|3917,3918
06|3919,3921
:|3921,3922
00AM|3922,3926
BLOOD|3927,3932
Glucose|3933,3940
-|3940,3941
147|3941,3944
*|3944,3945
UreaN|3946,3951
-|3951,3952
21|3952,3954
*|3954,3955
Creat|3956,3961
-|3961,3962
1|3962,3963
.|3963,3964
2|3964,3965
*|3965,3966
Na|3967,3969
-|3969,3970
139|3970,3973
<EOL>|3974,3975
K|3975,3976
-|3976,3977
3|3977,3978
.|3978,3979
0|3979,3980
*|3980,3981
Cl|3982,3984
-|3984,3985
99|3985,3987
HCO3|3988,3992
-|3992,3993
24|3993,3995
AnGap|3996,4001
-|4001,4002
19|4002,4004
<EOL>|4004,4005
_|4005,4006
_|4006,4007
_|4007,4008
06|4009,4011
:|4011,4012
00AM|4012,4016
BLOOD|4017,4022
Calcium|4023,4030
-|4030,4031
8.7|4031,4034
Phos|4035,4039
-|4039,4040
4.4|4040,4043
Mg|4044,4046
-|4046,4047
2.0|4047,4050
<EOL>|4050,4051
<EOL>|4051,4052
ECG|4052,4055
_|4056,4057
_|4057,4058
_|4058,4059
8|4060,4061
:|4061,4062
33|4062,4064
:|4064,4065
29|4065,4067
_|4068,4069
_|4069,4070
_|4070,4071
<EOL>|4071,4072
Baseline|4072,4080
artifact|4081,4089
.|4089,4090
Sinus|4091,4096
rhythm|4097,4103
.|4103,4104
Borderline|4105,4115
P|4116,4117
-|4117,4118
R|4118,4119
interval|4120,4128
<EOL>|4129,4130
prolongation|4130,4142
.|4142,4143
Prominent|4144,4153
voltage|4154,4161
in|4162,4164
leads|4165,4170
I|4171,4172
and|4173,4176
aVL|4177,4180
but|4181,4184
does|4185,4189
not|4190,4193
<EOL>|4194,4195
meet|4195,4199
criteria|4200,4208
for|4209,4212
left|4213,4217
ventricular|4218,4229
hypertrophy|4230,4241
.|4241,4242
There|4243,4248
are|4249,4252
marked|4253,4259
<EOL>|4260,4261
ST|4261,4263
segment|4264,4271
depressions|4272,4283
and|4284,4287
T|4288,4289
wave|4290,4294
inversions|4295,4305
in|4306,4308
leads|4309,4314
I|4315,4316
,|4316,4317
II|4318,4320
,|4320,4321
aVL|4322,4325
<EOL>|4326,4327
and|4327,4330
apical|4331,4337
lateral|4338,4345
leads|4346,4351
.|4351,4352
Compared|4353,4361
to|4362,4364
the|4365,4368
previous|4369,4377
tracing|4378,4385
of|4386,4388
<EOL>|4389,4390
_|4390,4391
_|4391,4392
_|4392,4393
the|4394,4397
rate|4398,4402
then|4403,4407
was|4408,4411
faster|4412,4418
.|4418,4419
ST|4420,4422
-|4422,4423
T|4423,4424
wave|4425,4429
abnormalities|4430,4443
were|4444,4448
<EOL>|4449,4450
similar|4450,4457
.|4457,4458
Consider|4459,4467
left|4468,4472
ventricular|4473,4484
hypertrophy|4485,4496
as|4497,4499
before|4500,4506
.|4506,4507
<EOL>|4508,4509
Clinical|4509,4517
correlation|4518,4529
is|4530,4532
suggested|4533,4542
.|4542,4543
<EOL>|4543,4544
<EOL>|4544,4545
CXR|4545,4548
_|4549,4550
_|4550,4551
_|4551,4552
<EOL>|4552,4553
Patient|4553,4560
is|4561,4563
status|4564,4570
post|4571,4575
median|4576,4582
sternotomy|4583,4593
and|4594,4597
CABG|4598,4602
.|4602,4603
Heart|4604,4609
size|4610,4614
is|4615,4617
<EOL>|4618,4619
normal|4619,4625
.|4625,4626
Mediastinal|4627,4638
and|4639,4642
hilar|4643,4648
contours|4649,4657
are|4658,4661
unchanged|4662,4671
.|4671,4672
Pulmonary|4673,4682
<EOL>|4683,4684
vasculature|4684,4695
is|4696,4698
normal|4699,4705
.|4705,4706
No|4707,4709
focal|4710,4715
consolidation|4716,4729
,|4729,4730
pleural|4731,4738
effusion|4739,4747
<EOL>|4748,4749
or|4749,4751
pneumothorax|4752,4764
is|4765,4767
seen|4768,4772
.|4772,4773
No|4774,4776
acute|4777,4782
osseous|4783,4790
abnormality|4791,4802
is|4803,4805
<EOL>|4806,4807
detected|4807,4815
.|4815,4816
<EOL>|4816,4817
IMPRESSION|4817,4827
:|4827,4828
No|4829,4831
acute|4832,4837
cardiopulmonary|4838,4853
abnormality|4854,4865
.|4865,4866
<EOL>|4866,4867
<EOL>|4867,4868
Dipyridamole|4868,4880
-|4880,4881
MIBI|4881,4885
Stress|4886,4892
test|4893,4897
_|4898,4899
_|4899,4900
_|4900,4901
<EOL>|4901,4902
_|4902,4903
_|4903,4904
_|4904,4905
yp|4906,4908
woman|4909,4914
with|4915,4919
HL|4920,4922
,|4922,4923
HTN|4924,4927
,|4927,4928
DM|4929,4931
,|4931,4932
PVD|4933,4936
and|4937,4940
diastolic|4941,4950
CHF|4951,4954
;|4954,4955
s|4956,4957
/|4957,4958
p|4958,4959
MI|4960,4962
and|4963,4966
<EOL>|4967,4968
multiple|4968,4976
PCIs|4977,4981
f|4982,4983
/|4983,4984
b|4984,4985
CABG|4986,4990
x|4991,4992
3|4993,4994
in|4995,4997
_|4998,4999
_|4999,5000
_|5000,5001
with|5002,5006
known|5007,5012
SVG|5013,5016
-|5016,5017
OM|5017,5019
occlusion|5020,5029
<EOL>|5030,5031
was|5031,5034
referred|5035,5043
to|5044,5046
evaluate|5047,5055
an|5056,5058
atypical|5059,5067
chest|5068,5073
discomfort|5074,5084
.|5084,5085
The|5086,5089
<EOL>|5090,5091
patient|5091,5098
was|5099,5102
administered|5103,5115
0.142|5116,5121
mg|5122,5124
/|5124,5125
kg|5125,5127
/|5127,5128
min|5128,5131
of|5132,5134
Persantine|5135,5145
over|5146,5150
4|5151,5152
<EOL>|5153,5154
minutes|5154,5161
.|5161,5162
Prior|5163,5168
to|5169,5171
the|5172,5175
procedure|5176,5185
the|5186,5189
patient|5190,5197
reported|5198,5206
an|5207,5209
isolated|5210,5218
<EOL>|5219,5220
left|5220,5224
-|5224,5225
sided|5225,5230
chest|5231,5236
discomfort|5237,5247
that|5248,5252
had|5253,5256
been|5257,5261
present|5262,5269
since|5270,5275
<EOL>|5276,5277
admission|5277,5286
and|5287,5290
was|5291,5294
tender|5295,5301
to|5302,5304
mild|5305,5309
palpation|5310,5319
;|5319,5320
_|5321,5322
_|5322,5323
_|5323,5324
.|5324,5325
This|5326,5330
<EOL>|5331,5332
discomfort|5332,5342
did|5343,5346
not|5347,5350
change|5351,5357
in|5358,5360
intensity|5361,5370
during|5371,5377
the|5378,5381
procedure|5382,5391
.|5391,5392
In|5393,5395
<EOL>|5396,5397
the|5397,5400
presence|5401,5409
of|5410,5412
diffuse|5413,5420
ST|5421,5423
-|5423,5424
T|5424,5425
wave|5426,5430
changes|5431,5438
,|5438,5439
no|5440,5442
additional|5443,5453
ECG|5454,5457
<EOL>|5458,5459
changes|5459,5466
were|5467,5471
noted|5472,5477
during|5478,5484
the|5485,5488
procedure|5489,5498
.|5498,5499
The|5500,5503
hemodynamic|5504,5515
<EOL>|5516,5517
response|5517,5525
to|5526,5528
the|5529,5532
Persantine|5533,5543
infusion|5544,5552
was|5553,5556
appropriate|5557,5568
.|5568,5569
<EOL>|5570,5571
Post-infusion|5571,5584
,|5584,5585
the|5586,5589
patient|5590,5597
was|5598,5601
administered|5602,5614
125|5615,5618
mg|5619,5621
Aminophylline|5622,5635
<EOL>|5636,5637
IV|5637,5639
.|5639,5640
<EOL>|5640,5641
IMPRESSION|5641,5651
:|5651,5652
Non-anginal|5653,5664
type|5665,5669
symptoms|5670,5678
with|5679,5683
no|5684,5686
additional|5687,5697
ST|5698,5700
<EOL>|5701,5702
segment|5702,5709
changes|5710,5717
from|5718,5722
baseline|5723,5731
.|5731,5732
<EOL>|5732,5733
Imaging|5733,5740
:|5740,5741
<EOL>|5741,5742
Left|5744,5748
ventricular|5749,5760
cavity|5761,5767
size|5768,5772
is|5773,5775
normal|5776,5782
.|5782,5783
<EOL>|5783,5784
Rest|5786,5790
and|5791,5794
stress|5795,5801
perfusion|5802,5811
images|5812,5818
reveal|5819,5825
uniform|5826,5833
tracer|5834,5840
uptake|5841,5847
<EOL>|5848,5849
throughout|5849,5859
the|5860,5863
left|5864,5868
ventricular|5869,5880
myocardium|5881,5891
.|5891,5892
The|5894,5897
previously|5898,5908
<EOL>|5909,5910
noted|5910,5915
perfusion|5916,5925
defect|5926,5932
involving|5933,5942
the|5943,5946
inferolateral|5947,5960
wall|5961,5965
has|5966,5969
<EOL>|5970,5971
resolved|5971,5979
.|5979,5980
<EOL>|5980,5981
Gated|5983,5988
images|5989,5995
reveal|5996,6002
normal|6003,6009
wall|6010,6014
motion|6015,6021
.|6021,6022
The|6023,6026
calculated|6027,6037
left|6038,6042
<EOL>|6043,6044
ventricular|6044,6055
ejection|6056,6064
fraction|6065,6073
is|6074,6076
64|6077,6079
%|6079,6080
.|6080,6081
<EOL>|6081,6082
IMPRESSION|6082,6092
:|6092,6093
Normal|6094,6100
myocardial|6101,6111
perfusion|6112,6121
study|6122,6127
.|6127,6128
Interval|6129,6137
<EOL>|6138,6139
normalization|6139,6152
of|6153,6155
prior|6156,6161
LCx|6162,6165
territory|6166,6175
perfusion|6176,6185
defect|6186,6192
.|6192,6193
<EOL>|6193,6194
<EOL>|6195,6196
This|6219,6223
is|6224,6226
a|6227,6228
_|6229,6230
_|6230,6231
_|6231,6232
with|6233,6237
type|6238,6242
2|6243,6244
diabetes|6245,6253
mellitus|6254,6262
on|6263,6265
insulin|6266,6273
,|6273,6274
CAD|6275,6278
s|6279,6280
/|6280,6281
p|6281,6282
<EOL>|6283,6284
MI|6284,6286
,|6286,6287
S|6288,6289
/|6289,6290
P|6290,6291
multiple|6292,6300
PCIs|6301,6305
and|6306,6309
CABG|6310,6314
_|6315,6316
_|6316,6317
_|6317,6318
(|6319,6320
LIMA|6320,6324
-|6324,6325
LAD|6325,6328
,|6328,6329
SVG|6330,6333
-|6333,6334
OM1|6334,6337
;|6337,6338
also|6339,6343
<EOL>|6344,6345
SVG|6345,6348
-|6348,6349
D1|6349,6351
known|6352,6357
occluded|6358,6366
_|6367,6368
_|6368,6369
_|6369,6370
with|6371,6375
chronic|6376,6383
stable|6384,6390
angina|6391,6397
<EOL>|6398,6399
admitted|6399,6407
with|6408,6412
atypical|6413,6421
,|6421,6422
stabbing|6423,6431
,|6431,6432
focal|6433,6438
chest|6439,6444
pain|6445,6449
.|6449,6450
<EOL>|6450,6451
<EOL>|6451,6452
#|6452,6453
Chest|6454,6459
pain|6460,6464
:|6464,6465
Initially|6466,6475
the|6476,6479
patient|6480,6487
was|6488,6491
started|6492,6499
on|6500,6502
a|6503,6504
heparin|6505,6512
<EOL>|6513,6514
drip|6514,6518
and|6519,6522
other|6523,6528
ACS|6529,6532
protocol|6533,6541
medications|6542,6553
.|6553,6554
Her|6555,6558
home|6559,6563
losartan|6564,6572
and|6573,6576
<EOL>|6577,6578
furosemide|6578,6588
were|6589,6593
held|6594,6598
due|6599,6602
to|6603,6605
low|6606,6609
blood|6610,6615
pressures|6616,6625
.|6625,6626
Suspicion|6627,6636
for|6637,6640
<EOL>|6641,6642
cardiac|6642,6649
etiology|6650,6658
of|6659,6661
chest|6662,6667
pain|6668,6672
was|6673,6676
ultimately|6677,6687
not|6688,6691
high|6692,6696
.|6696,6697
She|6698,6701
had|6702,6705
<EOL>|6706,6707
an|6707,6709
isolated|6710,6718
ongoing|6719,6726
_|6727,6728
_|6728,6729
_|6729,6730
left|6731,6735
-|6735,6736
sided|6736,6741
chest|6742,6747
discomfort|6748,6758
exacerbated|6759,6770
<EOL>|6771,6772
by|6772,6774
changes|6775,6782
in|6783,6785
position|6786,6794
and|6795,6798
with|6799,6803
chest|6804,6809
wall|6810,6814
tenderness|6815,6825
to|6826,6828
light|6829,6834
<EOL>|6835,6836
palpation|6836,6845
.|6845,6846
Despite|6847,6854
prolonged|6855,6864
chest|6865,6870
pain|6871,6875
,|6875,6876
troponin|6877,6885
-|6885,6886
T|6886,6887
and|6888,6891
CK|6892,6894
-|6894,6895
MB|6895,6897
<EOL>|6898,6899
negative|6899,6907
x2|6908,6910
and|6911,6914
EKGs|6915,6919
mostly|6920,6926
unchanged|6927,6936
from|6937,6941
prior|6942,6947
.|6947,6948
Given|6949,6954
known|6955,6960
<EOL>|6961,6962
H|6962,6963
/|6963,6964
O|6964,6965
CAD|6966,6969
,|6969,6970
a|6971,6972
vasodilator|6973,6984
nuclear|6985,6992
stress|6993,6999
test|7000,7004
was|7005,7008
performed|7009,7018
and|7019,7022
was|7023,7026
<EOL>|7027,7028
reassuring|7028,7038
.|7038,7039
Her|7040,7043
discomfort|7044,7054
did|7055,7058
not|7059,7062
change|7063,7069
in|7070,7072
intensity|7073,7082
during|7083,7089
<EOL>|7090,7091
the|7091,7094
stress|7095,7101
test|7102,7106
drug|7107,7111
infusion|7112,7120
.|7120,7121
In|7122,7124
the|7125,7128
presence|7129,7137
of|7138,7140
diffuse|7141,7148
ST|7149,7151
-|7151,7152
T|7152,7153
<EOL>|7154,7155
wave|7155,7159
changes|7160,7167
,|7167,7168
no|7169,7171
additional|7172,7182
ECG|7183,7186
changes|7187,7194
were|7195,7199
noted|7200,7205
during|7206,7212
the|7213,7216
<EOL>|7217,7218
procedure|7218,7227
.|7227,7228
The|7229,7232
hemodynamic|7233,7244
response|7245,7253
to|7254,7256
the|7257,7260
Persantine|7261,7271
infusion|7272,7280
<EOL>|7281,7282
was|7282,7285
appropriate|7286,7297
.|7297,7298
Her|7299,7302
perfusion|7303,7312
study|7313,7318
was|7319,7322
normal|7323,7329
with|7330,7334
interval|7335,7343
<EOL>|7344,7345
normalization|7345,7358
of|7359,7361
prior|7362,7367
LCx|7368,7371
territory|7372,7381
perfusion|7382,7391
defect|7392,7398
.|7398,7399
Given|7400,7405
the|7406,7409
<EOL>|7410,7411
stabbing|7411,7419
quality|7420,7427
and|7428,7431
tenderness|7432,7442
to|7443,7445
palpation|7446,7455
of|7456,7458
the|7459,7462
area|7463,7467
of|7468,7470
<EOL>|7471,7472
discomfort|7472,7482
,|7482,7483
her|7484,7487
symptoms|7488,7496
were|7497,7501
most|7502,7506
likely|7507,7513
related|7514,7521
to|7522,7524
<EOL>|7525,7526
costochondritis|7526,7541
or|7542,7544
other|7545,7550
musculoskeletal|7551,7566
causes|7567,7573
.|7573,7574
She|7575,7578
was|7579,7582
started|7583,7590
<EOL>|7591,7592
on|7592,7594
aspirin|7595,7602
650|7603,7606
mg|7607,7609
q6h|7610,7613
with|7614,7618
plans|7619,7624
to|7625,7627
trial|7628,7633
for|7634,7637
2|7638,7639
days|7640,7644
and|7645,7648
<EOL>|7649,7650
continue|7650,7658
through|7659,7666
the|7667,7670
week|7671,7675
if|7676,7678
symptoms|7679,7687
improve|7688,7695
.|7695,7696
<EOL>|7696,7697
<EOL>|7697,7698
Chronic|7698,7705
medical|7706,7713
problems|7714,7722
:|7722,7723
<EOL>|7723,7724
#|7724,7725
Diabetes|7726,7734
mellitus|7735,7743
:|7743,7744
Continued|7745,7754
levemir|7755,7762
and|7763,7766
was|7767,7770
switched|7771,7779
to|7780,7782
a|7783,7784
<EOL>|7785,7786
sliding|7786,7793
scale|7794,7799
of|7800,7802
Humalog|7803,7810
.|7810,7811
<EOL>|7811,7812
#|7812,7813
Hypertension|7814,7826
:|7826,7827
Losartan|7828,7836
was|7837,7840
held|7841,7845
as|7846,7848
above|7849,7854
due|7855,7858
to|7859,7861
hypotension|7862,7873
<EOL>|7874,7875
and|7875,7878
once|7879,7883
daily|7884,7889
isosorbide|7890,7900
mononitrate|7901,7912
was|7913,7916
switched|7917,7925
temporarily|7926,7937
<EOL>|7938,7939
to|7939,7941
isosorbide|7942,7952
dinitrate|7953,7962
TID|7963,7966
.|7966,7967
<EOL>|7968,7969
#|7969,7970
For|7971,7974
her|7975,7978
hyperlipidemia|7979,7993
,|7993,7994
COPD|7995,7999
and|8000,8003
GERD|8004,8008
,|8008,8009
her|8010,8013
home|8014,8018
regimens|8019,8027
were|8028,8032
<EOL>|8033,8034
continued|8034,8043
.|8043,8044
<EOL>|8046,8047
<EOL>|8047,8048
TRANSITIONAL|8048,8060
ISSUES|8061,8067
:|8067,8068
<EOL>|8068,8069
-|8069,8070
Patient|8071,8078
had|8079,8082
low|8083,8086
blood|8087,8092
pressures|8093,8102
initially|8103,8112
(|8113,8114
88|8114,8116
-|8116,8117
92|8117,8119
systolic|8120,8128
)|8128,8129
.|8129,8130
<EOL>|8131,8132
Would|8132,8137
benefit|8138,8145
from|8146,8150
close|8151,8156
monitoring|8157,8167
and|8168,8171
titration|8172,8181
of|8182,8184
blood|8185,8190
<EOL>|8191,8192
pressure|8192,8200
medications|8201,8212
as|8213,8215
an|8216,8218
outpatient|8219,8229
<EOL>|8229,8230
-|8230,8231
She|8232,8235
was|8236,8239
hypokalemic|8240,8251
(|8252,8253
K|8253,8254
3.0|8255,8258
)|8258,8259
during|8260,8266
admission|8267,8276
(|8277,8278
with|8278,8282
_|8283,8284
_|8284,8285
_|8285,8286
and|8287,8290
<EOL>|8291,8292
furosemide|8292,8302
already|8303,8310
held|8311,8315
)|8315,8316
.|8316,8317
Please|8318,8324
recheck|8325,8332
CHEM|8333,8337
-|8337,8338
10|8338,8340
at|8341,8343
_|8344,8345
_|8345,8346
_|8346,8347
_|8348,8349
_|8349,8350
_|8350,8351
<EOL>|8352,8353
visit|8353,8358
on|8359,8361
_|8362,8363
_|8363,8364
_|8364,8365
to|8366,8368
determine|8369,8378
whether|8379,8386
she|8387,8390
might|8391,8396
benefit|8397,8404
from|8405,8409
K|8410,8411
<EOL>|8412,8413
supplementation|8413,8428
<EOL>|8428,8429
-|8429,8430
Cr|8431,8433
elevated|8434,8442
to|8443,8445
1.2|8446,8449
on|8450,8452
discharge|8453,8462
(|8463,8464
up|8464,8466
from|8467,8471
most|8472,8476
recent|8477,8483
1.1|8484,8487
.1|8487,8489
)|8489,8490
.|8490,8491
<EOL>|8492,8493
Please|8493,8499
recheck|8500,8507
at|8508,8510
_|8511,8512
_|8512,8513
_|8513,8514
office|8515,8521
on|8522,8524
_|8525,8526
_|8526,8527
_|8527,8528
<EOL>|8528,8529
-|8529,8530
Full|8531,8535
code|8536,8540
<EOL>|8540,8541
<EOL>|8542,8543
Medications|8543,8554
on|8555,8557
Admission|8558,8567
:|8567,8568
<EOL>|8568,8569
The|8569,8572
Preadmission|8573,8585
Medication|8586,8596
list|8597,8601
is|8602,8604
accurate|8605,8613
and|8614,8617
complete|8618,8626
.|8626,8627
<EOL>|8627,8628
1.|8628,8630
Oxycodone|8631,8640
-|8640,8641
Acetaminophen|8641,8654
(|8655,8656
5mg|8656,8659
-|8659,8660
325mg|8660,8665
)|8665,8666
1|8667,8668
TAB|8669,8672
PO|8673,8675
Q8H|8676,8679
:|8679,8680
PRN|8680,8683
pain|8684,8688
<EOL>|8689,8690
2.|8690,8692
Nitroglycerin|8693,8706
SL|8707,8709
0.3|8710,8713
mg|8714,8716
SL|8717,8719
Q5MIN|8720,8725
:|8725,8726
PRN|8726,8729
pain|8730,8734
<EOL>|8735,8736
3.|8736,8738
Metoprolol|8739,8749
Succinate|8750,8759
XL|8760,8762
250|8763,8766
mg|8767,8769
PO|8770,8772
DAILY|8773,8778
<EOL>|8779,8780
4.|8780,8782
Levemir|8783,8790
Flexpen|8791,8798
(|8799,8800
insulin|8800,8807
detemir|8808,8815
)|8815,8816
90|8817,8819
units|8820,8825
subcutaneous|8826,8838
in|8839,8841
<EOL>|8842,8843
the|8843,8846
evening|8847,8854
<EOL>|8855,8856
5.|8856,8858
albuterol|8859,8868
sulfate|8869,8876
90|8877,8879
mcg|8880,8883
/|8883,8884
actuation|8884,8893
inhalation|8894,8904
q4hrs|8905,8910
wheezing|8911,8919
<EOL>|8920,8921
6.|8921,8923
Vitamin|8924,8931
D|8932,8933
1000|8934,8938
UNIT|8939,8943
PO|8944,8946
DAILY|8947,8952
<EOL>|8953,8954
7.|8954,8956
TraZODone|8957,8966
100|8967,8970
mg|8971,8973
PO|8974,8976
HS|8977,8979
<EOL>|8980,8981
8.|8981,8983
Isosorbide|8984,8994
Mononitrate|8995,9006
(|9007,9008
Extended|9008,9016
Release|9017,9024
)|9024,9025
120|9026,9029
mg|9030,9032
PO|9033,9035
DAILY|9036,9041
<EOL>|9042,9043
9.|9043,9045
Aspirin|9046,9053
325|9054,9057
mg|9058,9060
PO|9061,9063
DAILY|9064,9069
<EOL>|9070,9071
10.|9071,9074
Atorvastatin|9075,9087
80|9088,9090
mg|9091,9093
PO|9094,9096
HS|9097,9099
<EOL>|9100,9101
11.|9101,9104
Fluticasone|9105,9116
Propionate|9117,9127
110mcg|9128,9134
2|9135,9136
PUFF|9137,9141
IH|9142,9144
BID|9145,9148
<EOL>|9149,9150
12.|9150,9153
Pantoprazole|9154,9166
40|9167,9169
mg|9170,9172
PO|9173,9175
Q12H|9176,9180
<EOL>|9181,9182
13.|9182,9185
Ropinirole|9186,9196
0.5|9197,9200
mg|9201,9203
PO|9204,9206
QPM|9207,9210
<EOL>|9211,9212
14.|9212,9215
HumaLOG|9216,9223
KwikPen|9224,9231
(|9232,9233
insulin|9233,9240
lispro|9241,9247
)|9247,9248
0|9249,9250
SUBCUTANEOUS|9253,9265
AS|9266,9268
<EOL>|9269,9270
DIRECTED|9270,9278
<EOL>|9279,9280
15.|9280,9283
Albuterol|9284,9293
0.083|9294,9299
%|9299,9300
Neb|9301,9304
Soln|9305,9309
1|9310,9311
NEB|9312,9315
IH|9316,9318
Q6H|9319,9322
:|9322,9323
PRN|9323,9326
wheeze|9327,9333
<EOL>|9334,9335
16|9335,9337
.|9337,9338
Methocarbamol|9339,9352
500|9353,9356
mg|9357,9359
PO|9360,9362
TID|9363,9366
:|9366,9367
PRN|9367,9370
muscle|9371,9377
pain|9378,9382
<EOL>|9383,9384
17|9384,9386
.|9386,9387
Losartan|9388,9396
Potassium|9397,9406
25|9407,9409
mg|9410,9412
PO|9413,9415
DAILY|9416,9421
<EOL>|9422,9423
18.|9423,9426
Furosemide|9427,9437
20|9438,9440
mg|9441,9443
PO|9444,9446
DAILY|9447,9452
<EOL>|9453,9454
19.|9454,9457
diclofenac|9458,9468
sodium|9469,9475
1|9476,9477
%|9478,9479
topical|9480,9487
TID|9488,9491
:|9491,9492
PRN|9492,9495
pain|9496,9500
<EOL>|9500,9501
<EOL>|9502,9503
Discharge|9503,9512
Medications|9513,9524
:|9524,9525
<EOL>|9525,9526
1.|9526,9528
Albuterol|9529,9538
0.083|9539,9544
%|9544,9545
Neb|9546,9549
Soln|9550,9554
1|9555,9556
NEB|9557,9560
IH|9561,9563
Q6H|9564,9567
:|9567,9568
PRN|9568,9571
wheeze|9572,9578
<EOL>|9579,9580
2.|9580,9582
Atorvastatin|9583,9595
80|9596,9598
mg|9599,9601
PO|9602,9604
HS|9605,9607
<EOL>|9608,9609
3.|9609,9611
Fluticasone|9612,9623
Propionate|9624,9634
110mcg|9635,9641
2|9642,9643
PUFF|9644,9648
IH|9649,9651
BID|9652,9655
<EOL>|9656,9657
4.|9657,9659
Methocarbamol|9660,9673
500|9674,9677
mg|9678,9680
PO|9681,9683
TID|9684,9687
:|9687,9688
PRN|9688,9691
muscle|9692,9698
pain|9699,9703
<EOL>|9704,9705
5.|9705,9707
Nitroglycerin|9708,9721
SL|9722,9724
0.3|9725,9728
mg|9729,9731
SL|9732,9734
Q5MIN|9735,9740
:|9740,9741
PRN|9741,9744
pain|9745,9749
<EOL>|9750,9751
6.|9751,9753
Pantoprazole|9754,9766
40|9767,9769
mg|9770,9772
PO|9773,9775
Q12H|9776,9780
<EOL>|9781,9782
7.|9782,9784
Ropinirole|9785,9795
0.5|9796,9799
mg|9800,9802
PO|9803,9805
QPM|9806,9809
<EOL>|9810,9811
8.|9811,9813
TraZODone|9814,9823
100|9824,9827
mg|9828,9830
PO|9831,9833
HS|9834,9836
<EOL>|9837,9838
9.|9838,9840
Vitamin|9841,9848
D|9849,9850
1000|9851,9855
UNIT|9856,9860
PO|9861,9863
DAILY|9864,9869
<EOL>|9870,9871
10.|9871,9874
albuterol|9875,9884
sulfate|9885,9892
90|9893,9895
mcg|9896,9899
/|9899,9900
actuation|9900,9909
INHALATION|9910,9920
Q4HRS|9921,9926
wheezing|9927,9935
<EOL>|9935,9936
11.|9936,9939
diclofenac|9940,9950
sodium|9951,9957
1|9958,9959
%|9960,9961
topical|9962,9969
TID|9970,9973
:|9973,9974
PRN|9974,9977
pain|9978,9982
<EOL>|9983,9984
12.|9984,9987
Furosemide|9988,9998
20|9999,10001
mg|10002,10004
PO|10005,10007
DAILY|10008,10013
<EOL>|10014,10015
13.|10015,10018
Isosorbide|10019,10029
Mononitrate|10030,10041
(|10042,10043
Extended|10043,10051
Release|10052,10059
)|10059,10060
120|10061,10064
mg|10065,10067
PO|10068,10070
DAILY|10071,10076
<EOL>|10077,10078
14.|10078,10081
Metoprolol|10082,10092
Succinate|10093,10102
XL|10103,10105
250|10106,10109
mg|10110,10112
PO|10113,10115
DAILY|10116,10121
<EOL>|10122,10123
15.|10123,10126
HumaLOG|10127,10134
KwikPen|10135,10142
(|10143,10144
insulin|10144,10151
lispro|10152,10158
)|10158,10159
0|10160,10161
SUBCUTANEOUS|10164,10176
AS|10177,10179
<EOL>|10180,10181
DIRECTED|10181,10189
<EOL>|10190,10191
16|10191,10193
.|10193,10194
Levemir|10195,10202
Flexpen|10203,10210
(|10211,10212
insulin|10212,10219
detemir|10220,10227
)|10227,10228
90|10229,10231
units|10232,10237
subcutaneous|10238,10250
in|10251,10253
<EOL>|10254,10255
the|10255,10258
evening|10259,10266
<EOL>|10267,10268
17.|10268,10271
Losartan|10272,10280
Potassium|10281,10290
25|10291,10293
mg|10294,10296
PO|10297,10299
DAILY|10300,10305
<EOL>|10306,10307
18.|10307,10310
Oxycodone|10311,10320
-|10320,10321
Acetaminophen|10321,10334
(|10335,10336
5mg|10336,10339
-|10339,10340
325mg|10340,10345
)|10345,10346
1|10347,10348
TAB|10349,10352
PO|10353,10355
Q8H|10356,10359
:|10359,10360
PRN|10360,10363
pain|10364,10368
<EOL>|10369,10370
19|10370,10372
.|10372,10373
Aspirin|10374,10381
650|10382,10385
mg|10386,10388
PO|10389,10391
Q6H|10392,10395
<EOL>|10396,10397
RX|10397,10399
*|10400,10401
aspirin|10401,10408
650|10409,10412
mg|10413,10415
1|10416,10417
tablet|10418,10424
(|10424,10425
s|10425,10426
)|10426,10427
by|10428,10430
mouth|10431,10436
every|10437,10442
six|10443,10446
(|10447,10448
6|10448,10449
)|10449,10450
hours|10451,10456
Disp|10457,10461
<EOL>|10462,10463
#|10463,10464
*|10464,10465
28|10465,10467
Tablet|10468,10474
Refills|10475,10482
:|10482,10483
*|10483,10484
0|10484,10485
<EOL>|10485,10486
<EOL>|10487,10488
Discharge|10488,10497
Disposition|10498,10509
:|10509,10510
<EOL>|10510,10511
Home|10511,10515
<EOL>|10515,10516
<EOL>|10517,10518
Discharge|10518,10527
Diagnosis|10528,10537
:|10537,10538
<EOL>|10538,10539
-|10539,10540
Chest|10541,10546
wall|10547,10551
pain|10552,10556
atypical|10557,10565
for|10566,10569
angina|10570,10576
<EOL>|10576,10577
-|10577,10578
Musculoskeletal|10579,10594
pain|10595,10599
<EOL>|10599,10600
-|10600,10601
Known|10602,10607
native|10608,10614
coronary|10615,10623
artery|10624,10630
and|10631,10634
bypass|10635,10641
graft|10642,10647
disease|10648,10655
<EOL>|10655,10656
-|10656,10657
Type|10658,10662
2|10663,10664
Diabetes|10665,10673
mellitus|10674,10682
,|10682,10683
with|10684,10688
<EOL>|10688,10689
-|10689,10690
Chronic|10691,10698
kidney|10699,10705
disease|10706,10713
,|10713,10714
stage|10715,10720
3|10721,10722
<EOL>|10722,10723
-|10723,10724
Acute|10725,10730
kidney|10731,10737
injury|10738,10744
<EOL>|10744,10745
-|10745,10746
Chronic|10747,10754
obstructive|10755,10766
pulmonary|10767,10776
disease|10777,10784
<EOL>|10784,10785
-|10785,10786
Hypertension|10787,10799
<EOL>|10799,10800
-|10800,10801
Hypotension|10802,10813
<EOL>|10813,10814
-|10814,10815
Hypokalemia|10816,10827
<EOL>|10827,10828
-|10828,10829
Chronic|10830,10837
shoulder|10838,10846
pain|10847,10851
on|10852,10854
narcotics|10855,10864
<EOL>|10864,10865
-|10865,10866
Obstructive|10867,10878
sleep|10879,10884
apnea|10885,10890
<EOL>|10890,10891
-|10891,10892
Gastroseophageal|10893,10909
reflux|10910,10916
disease|10917,10924
<EOL>|10924,10925
<EOL>|10926,10927
Mental|10948,10954
Status|10955,10961
:|10961,10962
Clear|10963,10968
and|10969,10972
coherent|10973,10981
.|10981,10982
<EOL>|10982,10983
Level|10983,10988
of|10989,10991
Consciousness|10992,11005
:|11005,11006
Alert|11007,11012
and|11013,11016
interactive|11017,11028
.|11028,11029
<EOL>|11029,11030
Activity|11030,11038
Status|11039,11045
:|11045,11046
Ambulatory|11047,11057
-|11058,11059
Independent|11060,11071
.|11071,11072
<EOL>|11072,11073
<EOL>|11073,11074
<EOL>|11075,11076
Dear|11100,11104
Ms.|11105,11108
_|11109,11110
_|11110,11111
_|11111,11112
,|11112,11113
<EOL>|11113,11114
It|11114,11116
was|11117,11120
our|11121,11124
pleasure|11125,11133
participating|11134,11147
in|11148,11150
your|11151,11155
care|11156,11160
here|11161,11165
at|11166,11168
_|11169,11170
_|11170,11171
_|11171,11172
.|11172,11173
<EOL>|11174,11175
You|11175,11178
were|11179,11183
admitted|11184,11192
with|11193,11197
severe|11198,11204
chest|11205,11210
pain|11211,11215
.|11215,11216
You|11217,11220
underwent|11221,11230
a|11231,11232
stress|11233,11239
<EOL>|11240,11241
test|11241,11245
that|11246,11250
showed|11251,11257
the|11258,11261
pain|11262,11266
is|11267,11269
unlikely|11270,11278
from|11279,11283
a|11284,11285
big|11286,11289
blockage|11290,11298
in|11299,11301
the|11302,11305
<EOL>|11306,11307
arteries|11307,11315
that|11316,11320
feed|11321,11325
your|11326,11330
heart|11331,11336
.|11336,11337
Your|11338,11342
lab|11343,11346
work|11347,11351
also|11352,11356
did|11357,11360
not|11361,11364
<EOL>|11365,11366
suggest|11366,11373
injury|11374,11380
to|11381,11383
the|11384,11387
heart|11388,11393
.|11393,11394
<EOL>|11394,11395
<EOL>|11395,11396
The|11396,11399
pain|11400,11404
you|11405,11408
are|11409,11412
experiencing|11413,11425
is|11426,11428
most|11429,11433
likely|11434,11440
musculoskeletal|11441,11456
and|11457,11460
<EOL>|11461,11462
should|11462,11468
hopefully|11469,11478
improve|11479,11486
with|11487,11491
supportive|11492,11502
measures|11503,11511
such|11512,11516
as|11517,11519
<EOL>|11520,11521
Tylenol|11521,11528
(|11529,11530
maximum|11530,11537
3|11538,11539
grams|11540,11545
per|11546,11549
day|11550,11553
)|11553,11554
and|11555,11558
time|11559,11563
.|11563,11564
You|11565,11568
will|11569,11573
also|11574,11578
be|11579,11581
<EOL>|11582,11583
prescribed|11583,11593
high|11594,11598
dose|11599,11603
aspirin|11604,11611
(|11612,11613
650mg|11613,11618
)|11618,11619
.|11619,11620
Please|11621,11627
try|11628,11631
this|11632,11636
for|11637,11640
two|11641,11644
<EOL>|11645,11646
days|11646,11650
and|11651,11654
if|11655,11657
there|11658,11663
is|11664,11666
improvement|11667,11678
in|11679,11681
your|11682,11686
symptoms|11687,11695
continue|11696,11704
it|11705,11707
<EOL>|11708,11709
for|11709,11712
the|11713,11716
week|11717,11721
.|11721,11722
<EOL>|11723,11724
<EOL>|11724,11725
If|11725,11727
your|11728,11732
symptoms|11733,11741
worsen|11742,11748
,|11748,11749
you|11750,11753
develop|11754,11761
shortness|11762,11771
of|11772,11774
breath|11775,11781
or|11782,11784
any|11785,11788
<EOL>|11789,11790
other|11790,11795
concerning|11796,11806
symptom|11807,11814
,|11814,11815
please|11816,11822
let|11823,11826
your|11827,11831
doctor|11832,11838
know|11839,11843
right|11844,11849
<EOL>|11850,11851
away|11851,11855
.|11855,11856
<EOL>|11856,11857
<EOL>|11857,11858
Again|11858,11863
,|11863,11864
it|11865,11867
was|11868,11871
our|11872,11875
pleasure|11876,11884
participating|11885,11898
in|11899,11901
your|11902,11906
care|11907,11911
.|11911,11912
<EOL>|11912,11913
<EOL>|11913,11914
We|11914,11916
wish|11917,11921
you|11922,11925
the|11926,11929
very|11930,11934
_|11935,11936
_|11936,11937
_|11937,11938
,|11938,11939
<EOL>|11939,11940
Your|11940,11944
_|11945,11946
_|11946,11947
_|11947,11948
Cardiology|11949,11959
Team|11960,11964
<EOL>|11964,11965
<EOL>|11966,11967
Followup|11967,11975
Instructions|11976,11988
:|11988,11989
<EOL>|11989,11990
_|11990,11991
_|11991,11992
_|11992,11993
<EOL>|11993,11994

