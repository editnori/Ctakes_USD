 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|184,193|false|false|false|C1717415||Allergies
Event|Event|Allergies|184,193|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|184,193|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|196,218|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|204,208|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|204,208|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|204,218|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|209,218|false|false|false|||Reactions
Event|Event|Allergies|221,230|false|false|false|||Attending
Finding|Functional Concept|Allergies|221,230|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|260,275|false|false|false|||tachyarrhythmia
Finding|Finding|Chief Complaint|260,275|false|false|false|C0080203|Tachyarrhythmia|tachyarrhythmia
Finding|Classification|Chief Complaint|278,283|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|284,292|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|296,314|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|305,314|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|305,314|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|305,314|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|305,314|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|305,314|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|History of Present Illness|361,367|false|false|false|||smoker
Finding|Finding|History of Present Illness|361,367|false|false|false|C0337664;C3241966|Current Smoker;Smoker|smoker
Event|Event|History of Present Illness|373,376|false|false|false|||PMH
Finding|Finding|History of Present Illness|373,376|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|History of Present Illness|380,386|false|false|false|C0004096|Asthma|asthma
Event|Event|History of Present Illness|380,386|false|false|false|||asthma
Disorder|Disease or Syndrome|History of Present Illness|387,391|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|387,391|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|387,391|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|387,391|false|false|false|C1412502|ARCN1 gene|COPD
Drug|Organic Chemical|History of Present Illness|395,407|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|395,407|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|395,407|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|395,407|false|false|false|C0039773|Assay of theophylline|theophylline
Disorder|Disease or Syndrome|History of Present Illness|409,412|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|409,412|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|409,412|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|409,412|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|409,412|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|409,412|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|409,412|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|409,412|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|415,418|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|History of Present Illness|415,418|false|false|false|||HTN
Disorder|Disease or Syndrome|History of Present Illness|420,434|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|History of Present Illness|420,434|false|false|false|||hyperlipidemia
Finding|Finding|History of Present Illness|420,434|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Finding|Finding|History of Present Illness|440,448|false|false|false|C0741302|atypia morphology|atypical
Finding|Sign or Symptom|History of Present Illness|440,459|false|false|false|C0262384|Atypical chest pain|atypical chest pain
Anatomy|Body Location or Region|History of Present Illness|449,454|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|449,454|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|449,459|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|449,459|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|455,459|false|false|false|C2598155||pain
Event|Event|History of Present Illness|455,459|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|455,459|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|455,459|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|460,470|false|false|false|||presenting
Event|Event|History of Present Illness|477,484|false|false|false|||malaise
Finding|Sign or Symptom|History of Present Illness|477,484|false|false|false|C0231218|Malaise|malaise
Event|Event|History of Present Illness|489,492|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|489,492|false|false|false|C0013404|Dyspnea|SOB
Event|Event|History of Present Illness|503,510|false|false|false|||episode
Event|Event|History of Present Illness|514,528|false|false|false|||tachyarrythmia
Finding|Finding|History of Present Illness|529,536|false|false|false|C4534363|At home|at home
Event|Event|History of Present Illness|532,536|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|532,536|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|532,536|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|532,536|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|554,562|false|false|false|||resolved
Event|Event|History of Present Illness|568,575|false|false|false|||recalls
Event|Event|History of Present Illness|585,589|false|false|false|||took
Event|Event|History of Present Illness|605,615|false|false|false|||telehealth
Procedure|Health Care Activity|History of Present Illness|605,615|false|false|false|C0162648;C1328956|Telehealth;Telemedicine|telehealth
Drug|Hazardous or Poisonous Substance|History of Present Illness|616,623|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|History of Present Illness|616,623|false|false|false|C0728873|Monitor brand of insecticide|monitor
Event|Event|History of Present Illness|616,623|false|false|false|||monitor
Finding|Intellectual Product|History of Present Illness|625,629|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|636,642|false|false|false|||called
Event|Event|History of Present Illness|647,652|false|false|false|||asked
Event|Event|History of Present Illness|661,668|false|false|false|||recheck
Event|Event|History of Present Illness|680,688|false|false|false|||services
Event|Occupational Activity|History of Present Illness|680,688|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|History of Present Illness|680,688|false|false|false|C1704289|Clinical Service|services
Event|Event|History of Present Illness|698,706|false|false|false|||measured
Event|Event|History of Present Illness|743,746|false|false|false|||SOB
Finding|Sign or Symptom|History of Present Illness|743,746|true|false|false|C0013404|Dyspnea|SOB
Finding|Functional Concept|History of Present Illness|748,754|false|false|false|C0234621|Visual|visual
Event|Event|History of Present Illness|763,768|false|false|false|||palps
Finding|Conceptual Entity|History of Present Illness|763,768|false|false|false|C2945620|Palp - CHV concept|palps
Event|Event|History of Present Illness|776,782|false|false|false|||denies
Anatomy|Body Location or Region|History of Present Illness|794,797|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|abd
Disorder|Cell or Molecular Dysfunction|History of Present Illness|794,797|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|abd
Attribute|Clinical Attribute|History of Present Illness|798,802|false|false|false|C2598155||pain
Event|Event|History of Present Illness|798,802|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|798,802|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|798,802|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|804,810|false|false|false|||change
Finding|Functional Concept|History of Present Illness|804,810|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|804,810|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|History of Present Illness|804,813|false|false|false|C0392747|Changing|change in
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|814,819|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|823,830|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|823,830|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|History of Present Illness|823,830|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|823,830|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Disease or Syndrome|History of Present Illness|841,844|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|841,844|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|841,844|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|841,844|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|841,844|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|841,844|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|841,844|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|841,844|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|841,844|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|841,844|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|841,844|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|History of Present Illness|860,867|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|860,867|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|860,867|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|880,887|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|880,887|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|880,887|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|880,887|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|880,890|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|891,906|false|false|false|||tachyarrythmias
Finding|Body Substance|History of Present Illness|924,931|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|924,931|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|924,931|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|932,938|false|false|false|||denies
Event|Event|History of Present Illness|944,951|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|944,951|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|944,951|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|944,951|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Drug|Organic Chemical|History of Present Illness|969,981|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|969,981|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|969,981|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|969,981|false|false|false|C0039773|Assay of theophylline|theophylline
Finding|Finding|History of Present Illness|991,995|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|991,995|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|991,995|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Congenital Abnormality|History of Present Illness|1023,1026|false|true|false|C0026760|Multiple Epiphyseal Dysplasia|med
Finding|Gene or Genome|History of Present Illness|1023,1026|false|true|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Finding|Intellectual Product|History of Present Illness|1023,1026|false|true|false|C1413596;C1413597;C1419866;C1456376;C1549978;C4321267;C5781216|COL9A2 gene;COL9A3 gene;COMP gene;COMP wt Allele;Master of Education;SCN8A gene;SCN8A wt Allele|med
Event|Event|History of Present Illness|1027,1031|false|false|false|||list
Finding|Intellectual Product|History of Present Illness|1027,1031|false|true|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|History of Present Illness|1041,1047|false|false|false|||states
Event|Event|History of Present Illness|1059,1064|false|false|false|||taken
Disorder|Disease or Syndrome|History of Present Illness|1089,1092|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1089,1092|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|History of Present Illness|1089,1092|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1089,1092|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|History of Present Illness|1089,1092|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|History of Present Illness|1089,1092|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|History of Present Illness|1089,1092|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|History of Present Illness|1089,1092|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|History of Present Illness|1089,1092|false|false|false|||PCP
Finding|Gene or Genome|History of Present Illness|1089,1092|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|History of Present Illness|1089,1092|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|History of Present Illness|1094,1101|false|false|false|||concern
Finding|Idea or Concept|History of Present Illness|1094,1101|false|false|false|C2699424|Concern|concern
Drug|Organic Chemical|History of Present Illness|1114,1126|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|1114,1126|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|1114,1126|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|1114,1126|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|History of Present Illness|1134,1146|false|false|false|||contributing
Attribute|Clinical Attribute|History of Present Illness|1157,1163|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|History of Present Illness|1157,1163|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|History of Present Illness|1157,1163|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|History of Present Illness|1157,1163|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|History of Present Illness|1157,1168|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|History of Present Illness|1164,1168|false|false|false|C4318744|Test - temporal region|test
Event|Event|History of Present Illness|1164,1168|false|false|false|||test
Finding|Functional Concept|History of Present Illness|1164,1168|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|History of Present Illness|1164,1168|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|History of Present Illness|1164,1168|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|History of Present Illness|1164,1168|false|false|false|C0022885|Laboratory Procedures|test
Finding|Functional Concept|History of Present Illness|1174,1184|false|false|false|C0205343|Reversible|reversible
Event|Event|History of Present Illness|1185,1191|false|false|false|||lesion
Finding|Finding|History of Present Illness|1185,1191|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|History of Present Illness|1185,1191|false|false|false|C0221198;C1546698|Lesion|lesion
Event|Event|History of Present Illness|1198,1205|false|false|false|||treated
Event|Event|History of Present Illness|1271,1274|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|1271,1274|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|1292,1304|false|false|false|||unremarkable
Event|Event|History of Present Illness|1307,1315|false|false|false|||Transfer
Finding|Functional Concept|History of Present Illness|1307,1315|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|History of Present Illness|1307,1315|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|History of Present Illness|1307,1315|false|false|false|C4706767|Transfer (immobility management)|Transfer
Event|Event|History of Present Illness|1324,1326|false|false|false|||HR
Event|Event|History of Present Illness|1331,1333|false|false|false|||BP
Event|Event|History of Present Illness|1342,1344|false|false|false|||RR
Event|Event|History of Present Illness|1349,1352|false|false|false|||POx
Finding|Gene or Genome|History of Present Illness|1349,1352|false|false|false|C1418945|PRODH gene|POx
Anatomy|Anatomical Structure|History of Present Illness|1370,1375|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|1380,1392|false|false|false|||asymptomatic
Finding|Finding|History of Present Illness|1380,1392|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|History of Present Illness|1397,1402|false|false|false|||feels
Finding|Finding|History of Present Illness|1403,1407|false|false|false|C5575035|Well (answer to question)|well
Finding|Mental Process|History of Present Illness|1415,1420|false|false|false|C3887804|Feeling upset|upset
Finding|Idea or Concept|History of Present Illness|1448,1456|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|History of Present Illness|1463,1468|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|1463,1468|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Procedure|Laboratory Procedure|History of Present Illness|1472,1475|false|false|false|C5400981|Fibrinogen to Albumin Ratio Measurement|far
Finding|Idea or Concept|History of Present Illness|1481,1485|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|1481,1485|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Disorder|Disease or Syndrome|Past Medical History|1513,1519|false|false|false|C0004096|Asthma|ASTHMA
Event|Event|Past Medical History|1513,1519|false|false|false|||ASTHMA
Disorder|Disease or Syndrome|Past Medical History|1524,1536|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|1524,1536|false|false|false|||HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|1541,1555|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|1541,1555|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|1541,1555|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Finding|Sign or Symptom|Past Medical History|1560,1568|false|false|false|C0018681|Headache|HEADACHE
Disorder|Disease or Syndrome|Past Medical History|1573,1587|false|false|false|C0029408|Degenerative polyarthritis|OSTEOARTHRITIS
Event|Event|Past Medical History|1573,1587|false|false|false|||OSTEOARTHRITIS
Finding|Finding|Past Medical History|1592,1600|false|false|false|C0741302|atypia morphology|ATYPICAL
Finding|Sign or Symptom|Past Medical History|1592,1611|false|false|false|C0262384|Atypical chest pain|ATYPICAL CHEST PAIN
Anatomy|Body Location or Region|Past Medical History|1601,1606|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1601,1606|false|false|false|C0741025|Chest problem|CHEST
Attribute|Clinical Attribute|Past Medical History|1601,1611|false|false|false|C2926613||CHEST PAIN
Finding|Sign or Symptom|Past Medical History|1601,1611|false|false|false|C0008031|Chest Pain|CHEST PAIN
Attribute|Clinical Attribute|Past Medical History|1607,1611|false|true|false|C2598155||PAIN
Event|Event|Past Medical History|1607,1611|false|false|false|||PAIN
Finding|Functional Concept|Past Medical History|1607,1611|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Past Medical History|1607,1611|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Drug|Hazardous or Poisonous Substance|Past Medical History|1616,1623|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Past Medical History|1616,1623|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Past Medical History|1616,1623|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Past Medical History|1616,1623|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1616,1629|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1624,1629|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Past Medical History|1624,1629|false|false|false|||ABUSE
Event|Event|Past Medical History|1624,1629|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Past Medical History|1624,1629|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Finding|Past Medical History|1634,1642|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Idea or Concept|Past Medical History|1634,1642|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Finding|Past Medical History|1634,1648|false|false|false|C0742257|chest abnormal|ABNORMAL CHEST
Finding|Finding|Past Medical History|1634,1653|false|false|false|C0436503|Standard chest X-ray abnormal|ABNORMAL CHEST XRAY
Anatomy|Body Location or Region|Past Medical History|1643,1648|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|CHEST
Finding|Finding|Past Medical History|1643,1648|false|false|false|C0741025|Chest problem|CHEST
Procedure|Diagnostic Procedure|Past Medical History|1643,1653|false|false|false|C0039985|Plain chest X-ray|CHEST XRAY
Event|Event|Past Medical History|1649,1653|false|false|false|||XRAY
Phenomenon|Natural Phenomenon or Process|Past Medical History|1649,1653|false|false|false|C0043309|Roentgen Rays|XRAY
Procedure|Diagnostic Procedure|Past Medical History|1649,1653|false|false|false|C0043299|Diagnostic radiologic examination|XRAY
Disorder|Disease or Syndrome|Past Medical History|1658,1662|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|1658,1662|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|1658,1662|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|1658,1662|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Idea or Concept|Family Medical History|1704,1710|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|1717,1720|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Family Medical History|1717,1720|false|false|false|||HTN
Finding|Conceptual Entity|Family Medical History|1723,1729|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1723,1729|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|Family Medical History|1740,1747|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|1740,1747|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1740,1747|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|1755,1762|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|1755,1762|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|1755,1762|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Event|Event|Family Medical History|1772,1780|false|false|false|||Physical
Finding|Finding|Family Medical History|1772,1780|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|Family Medical History|1772,1780|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|Family Medical History|1772,1780|false|false|false|C0031809|Physical Examination|Physical
Procedure|Health Care Activity|Family Medical History|1786,1795|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|Family Medical History|1796,1799|false|false|false|||PEx
Finding|Gene or Genome|Family Medical History|1796,1799|false|false|false|C1418526;C5891011|PHEX gene;PHEX wt Allele|PEx
Disorder|Disease or Syndrome|Family Medical History|1844,1847|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|Family Medical History|1844,1847|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|Family Medical History|1844,1847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Family Medical History|1844,1847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|Family Medical History|1844,1847|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|Family Medical History|1844,1847|false|false|false|||NAD
Finding|Finding|Family Medical History|1844,1847|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|Family Medical History|1848,1853|false|false|false|C1512338|HEENT|HEENT
Event|Event|Family Medical History|1856,1862|false|false|false|||PERRLA
Finding|Finding|Family Medical History|1856,1862|false|false|false|C2143306|PERRLA|PERRLA
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1864,1867|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|Family Medical History|1864,1867|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|Family Medical History|1864,1867|false|false|false|||MMM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1872,1875|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Family Medical History|1872,1875|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|Family Medical History|1872,1875|false|false|false|||LAD
Finding|Gene or Genome|Family Medical History|1872,1875|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|Family Medical History|1880,1883|false|false|false|||JVD
Finding|Finding|Family Medical History|1880,1883|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Location or Region|Family Medical History|1885,1889|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Family Medical History|1885,1889|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Family Medical History|1885,1889|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|Family Medical History|1885,1896|false|false|false|C2230237|Supple neck|neck supple
Event|Event|Family Medical History|1890,1896|false|false|false|||supple
Finding|Functional Concept|Family Medical History|1890,1896|false|false|false|C0332254|Supple|supple
Event|Event|Family Medical History|1906,1909|false|false|false|||PMI
Finding|Finding|Family Medical History|1906,1909|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Finding|Gene or Genome|Family Medical History|1906,1909|false|false|false|C1417244;C1418674;C1823304;C5238618;C5780972|MPI gene;PMM2 gene;PMM2 wt Allele;Point of Maximum Impulse;TMEM11 gene|PMI
Phenomenon|Natural Phenomenon or Process|Family Medical History|1929,1934|false|false|false|C0282173|Space (Astronomy)|space
Disorder|Disease or Syndrome|Family Medical History|1939,1942|true|false|false|C0162770|Right Ventricular Hypertrophy|RVH
Event|Event|Family Medical History|1939,1942|false|false|false|||RVH
Event|Event|Family Medical History|1948,1950|false|false|false|||S1
Event|Event|Family Medical History|1954,1959|false|false|false|||heard
Event|Event|Family Medical History|1965,1972|false|false|false|||murmurs
Finding|Finding|Family Medical History|1965,1972|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|Family Medical History|1981,1985|false|false|false|||rubs
Finding|Finding|Family Medical History|1981,1985|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|Family Medical History|1987,1991|false|false|false|||Pulm
Procedure|Health Care Activity|Family Medical History|1987,1991|false|false|false|C1315068|Pulmonary ventilator management|Pulm
Finding|Gene or Genome|Family Medical History|2003,2006|false|false|false|C1417055|MBNL1 gene|exp
Event|Event|Family Medical History|2007,2015|false|false|false|||wheezing
Finding|Sign or Symptom|Family Medical History|2007,2015|false|false|false|C0043144|Wheezing|wheezing
Drug|Inorganic Chemical|Family Medical History|2029,2032|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Family Medical History|2029,2032|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Family Medical History|2029,2032|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Family Medical History|2029,2032|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Family Medical History|2029,2032|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Family Medical History|2029,2032|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Event|Event|Family Medical History|2033,2040|false|false|false|||movment
Anatomy|Body Location or Region|Family Medical History|2041,2044|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|Abd
Disorder|Cell or Molecular Dysfunction|Family Medical History|2041,2044|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|Abd
Disorder|Disease or Syndrome|Family Medical History|2046,2050|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|Family Medical History|2046,2050|false|false|false|||soft
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2070,2081|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|Family Medical History|2091,2096|true|false|false|C1717255||edema
Event|Event|Family Medical History|2091,2096|false|false|false|||edema
Finding|Pathologic Function|Family Medical History|2091,2096|true|false|false|C0013604|Edema|edema
Event|Event|Family Medical History|2098,2101|false|false|false|||DPs
Finding|Gene or Genome|Family Medical History|2098,2101|false|false|false|C1843919|PDSS1 gene|DPs
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2103,2106|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Enzyme|Family Medical History|2103,2106|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Organic Chemical|Family Medical History|2103,2106|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Drug|Pharmacologic Substance|Family Medical History|2103,2106|false|false|false|C0048719;C5958725|4-toluenesulfonamide;PTS protein, human|PTs
Event|Event|Family Medical History|2103,2106|false|false|false|||PTs
Finding|Gene or Genome|Family Medical History|2103,2106|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Finding|Intellectual Product|Family Medical History|2103,2106|false|false|false|C1419129;C2698747|PTS gene;Patient Tracking System|PTs
Anatomy|Body System|Family Medical History|2111,2115|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|Family Medical History|2111,2115|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|Family Medical History|2111,2115|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|Family Medical History|2111,2115|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|Family Medical History|2111,2115|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|Family Medical History|2120,2126|false|false|false|||rashes
Finding|Sign or Symptom|Family Medical History|2120,2126|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Event|Event|Family Medical History|2128,2137|false|false|false|||eccymoses
Event|Event|Family Medical History|2139,2146|false|false|false|||lesions
Finding|Finding|Family Medical History|2139,2146|true|false|false|C0221198|Lesion|lesions
Disorder|Mental or Behavioral Dysfunction|Family Medical History|2154,2159|false|false|false|C0004936;C1306597|Mental disorders;Psychiatric problem|Psych
Anatomy|Body System|Family Medical History|2161,2164|false|false|false|C3714787|Central Nervous System|CNs
Event|Event|Family Medical History|2172,2178|false|false|false|||intact
Finding|Finding|Family Medical History|2172,2178|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|Family Medical History|2184,2192|false|false|false|||strength
Finding|Idea or Concept|Family Medical History|2184,2192|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2196,2202|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|Family Medical History|2196,2202|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Event|Event|Family Medical History|2203,2209|false|false|false|||groups
Finding|Idea or Concept|Family Medical History|2203,2209|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Finding|Intellectual Product|Family Medical History|2203,2209|false|false|false|C0441833;C1552839|Groups;Table Rules - groups|groups
Event|Event|Family Medical History|2211,2217|false|false|false|||tested
Event|Event|Family Medical History|2219,2228|false|false|false|||sensation
Finding|Finding|Family Medical History|2219,2228|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Family Medical History|2219,2228|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Family Medical History|2219,2228|false|false|false|C2229507|sensory exam|sensation
Event|Event|Family Medical History|2229,2238|false|false|false|||symmetric
Finding|Conceptual Entity|Family Medical History|2229,2238|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|Family Medical History|2229,2238|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|Family Medical History|2242,2251|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Family Medical History|2242,2251|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Family Medical History|2242,2251|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Family Medical History|2242,2251|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|Family Medical History|2252,2255|false|false|false|||PEx
Finding|Gene or Genome|Family Medical History|2252,2255|false|false|false|C1418526;C5891011|PHEX gene;PHEX wt Allele|PEx
Event|Activity|Family Medical History|2292,2306|false|false|false|C1882932|Representation (action)|representative
Lab|Laboratory or Test Result|Family Medical History|2307,2311|false|false|false|C0587081|Laboratory test finding|labs
Anatomy|Cell Component|Family Medical History|2313,2316|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|Family Medical History|2313,2316|false|false|false|||CBC
Procedure|Laboratory Procedure|Family Medical History|2313,2316|false|false|false|C0009555|Complete Blood Count|CBC
Disorder|Disease or Syndrome|Family Medical History|2341,2346|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2341,2346|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2341,2346|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2347,2350|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2355,2358|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2355,2358|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2355,2358|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2364,2367|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2364,2367|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2364,2367|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2364,2367|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2373,2376|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2373,2376|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2383,2386|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|2383,2386|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|2383,2386|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2383,2386|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2383,2386|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2390,2393|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2390,2393|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|2390,2393|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|2390,2393|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2390,2393|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2390,2393|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|2399,2403|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|2399,2403|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|Family Medical History|2409,2412|false|false|false|||RDW
Procedure|Laboratory Procedure|Family Medical History|2419,2422|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2440,2445|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2440,2445|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2440,2445|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Family Medical History|2446,2449|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Family Medical History|2454,2457|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Family Medical History|2454,2457|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Family Medical History|2454,2457|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2463,2466|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Family Medical History|2463,2466|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Family Medical History|2463,2466|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Family Medical History|2463,2466|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Family Medical History|2472,2475|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2472,2475|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Family Medical History|2482,2485|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|Family Medical History|2482,2485|false|false|false|||MCV
Lab|Laboratory or Test Result|Family Medical History|2482,2485|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Family Medical History|2482,2485|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2482,2485|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Family Medical History|2489,2492|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Family Medical History|2489,2492|false|false|false|C0600370|methacholine|MCH
Event|Event|Family Medical History|2489,2492|false|false|false|||MCH
Finding|Gene or Genome|Family Medical History|2489,2492|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Family Medical History|2489,2492|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Family Medical History|2489,2492|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|Family Medical History|2498,2502|false|false|false|||MCHC
Procedure|Laboratory Procedure|Family Medical History|2498,2502|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|Family Medical History|2508,2511|false|false|false|||RDW
Procedure|Laboratory Procedure|Family Medical History|2518,2521|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Family Medical History|2539,2544|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2539,2544|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2539,2544|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|Family Medical History|2549,2552|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|Family Medical History|2549,2552|false|false|false|||PTT
Procedure|Laboratory Procedure|Family Medical History|2549,2552|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Event|Event|Family Medical History|2563,2567|false|false|false|||Chem
Finding|Functional Concept|Family Medical History|2563,2567|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|Family Medical History|2563,2567|false|false|false|C0201682|Chemical procedure|Chem
Disorder|Disease or Syndrome|Family Medical History|2582,2587|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2582,2587|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2582,2587|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|2582,2595|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|2582,2595|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|2582,2595|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|2588,2595|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|2588,2595|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|2588,2595|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|2588,2595|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|2588,2595|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|2588,2595|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|2641,2645|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|2641,2645|false|false|false|C0005367|Bicarbonates|HCO3
Event|Event|Family Medical History|2641,2645|false|false|false|||HCO3
Procedure|Laboratory Procedure|Family Medical History|2641,2645|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Family Medical History|2663,2668|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2663,2668|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2663,2668|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Family Medical History|2663,2676|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Family Medical History|2663,2676|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Family Medical History|2663,2676|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Family Medical History|2669,2676|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Family Medical History|2669,2676|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Family Medical History|2669,2676|false|false|false|C0017725|glucose|Glucose
Event|Event|Family Medical History|2669,2676|false|false|false|||Glucose
Lab|Laboratory or Test Result|Family Medical History|2669,2676|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Family Medical History|2669,2676|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Family Medical History|2721,2725|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Family Medical History|2721,2725|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Family Medical History|2721,2725|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Congenital Abnormality|Family Medical History|2730,2733|false|false|false|C0265493;C1963580|Cat eye syndrome;Congenital stenosis of esophagus|CEs
Disorder|Disease or Syndrome|Family Medical History|2730,2733|false|false|false|C0265493;C1963580|Cat eye syndrome;Congenital stenosis of esophagus|CEs
Event|Event|Family Medical History|2730,2733|false|false|false|||CEs
Finding|Intellectual Product|Family Medical History|2730,2733|false|false|false|C4318461|Combat Exposure Scale Questionnaire|CEs
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2730,2733|false|false|false|C3899490|Cranial Electrical Stimulation|CEs
Disorder|Disease or Syndrome|Family Medical History|2748,2753|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2748,2753|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2748,2753|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|Family Medical History|2781,2786|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2781,2786|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2781,2786|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2787,2792|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|2787,2792|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|2787,2792|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|2787,2792|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|Family Medical History|2822,2827|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2822,2827|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2822,2827|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2828,2833|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|Family Medical History|2828,2833|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|Family Medical History|2828,2833|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|Family Medical History|2828,2833|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|Family Medical History|2831,2835|false|false|false|C0602254|MB 3|MB-3
Disorder|Disease or Syndrome|Family Medical History|2851,2855|false|false|false|C5391534|multisystem inflammatory syndrome in children with COVID-19 infection|Misc
Event|Event|Family Medical History|2851,2855|false|false|false|||Misc
Disorder|Disease or Syndrome|Family Medical History|2870,2875|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|Family Medical History|2870,2875|false|false|false|||BLOOD
Finding|Body Substance|Family Medical History|2870,2875|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2887,2890|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|Family Medical History|2887,2890|false|false|false|C0023821|High Density Lipoproteins|HDL
Event|Event|Family Medical History|2887,2890|false|false|false|||HDL
Finding|Gene or Genome|Family Medical History|2887,2890|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|Family Medical History|2887,2890|false|false|false|C0392885|High density lipoprotein measurement|HDL
Event|Event|Hospital Course|2965,2971|false|false|false|||follow
Drug|Organic Chemical|Hospital Course|2975,2987|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|2975,2987|false|false|false|C0039771|theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|2975,2987|false|false|false|C0039773|Assay of theophylline|theophylline
Procedure|Laboratory Procedure|Hospital Course|2975,2993|false|false|false|C0039773|Assay of theophylline|theophylline level
Event|Event|Hospital Course|2988,2993|false|false|false|||level
Event|Event|Hospital Course|3003,3009|false|false|false|||smoker
Finding|Finding|Hospital Course|3003,3009|false|false|false|C0337664;C3241966|Current Smoker;Smoker|smoker
Event|Event|Hospital Course|3015,3018|false|false|false|||PMH
Finding|Finding|Hospital Course|3015,3018|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|Hospital Course|3022,3028|false|false|false|C0004096|Asthma|asthma
Event|Event|Hospital Course|3022,3028|false|false|false|||asthma
Disorder|Disease or Syndrome|Hospital Course|3029,3033|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|3029,3033|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|3029,3033|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|3029,3033|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|3034,3041|false|false|false|||managed
Drug|Organic Chemical|Hospital Course|3047,3059|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|3047,3059|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|3047,3059|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|3047,3059|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Hospital Course|3076,3088|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|3076,3088|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|3076,3088|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|3076,3088|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Hospital Course|3093,3105|false|false|false|||discontinued
Event|Event|Hospital Course|3118,3129|false|false|false|||tachycardia
Finding|Finding|Hospital Course|3118,3129|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Disorder|Disease or Syndrome|Hospital Course|3131,3134|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3131,3134|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|3131,3134|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|3131,3134|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|3131,3134|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|3131,3134|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|3131,3134|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3131,3134|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|3136,3139|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|3136,3139|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|3145,3159|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Hospital Course|3145,3159|false|false|false|||hyperlipidemia
Finding|Finding|Hospital Course|3145,3159|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|Hospital Course|3164,3173|false|false|false|||presented
Event|Event|Hospital Course|3180,3184|false|false|false|||home
Finding|Idea or Concept|Hospital Course|3180,3184|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|3180,3184|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|3180,3184|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|3190,3202|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|Hospital Course|3203,3217|false|false|false|||tachyarrythmia
Event|Event|Hospital Course|3230,3236|false|false|false|||ISSUES
Event|Event|Hospital Course|3242,3256|false|false|false|||Tachycarrhymia
Event|Event|Hospital Course|3260,3267|false|false|false|||context
Finding|Idea or Concept|Hospital Course|3260,3267|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|Hospital Course|3260,3267|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|Hospital Course|3260,3267|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Functional Concept|Hospital Course|3278,3287|false|false|false|C0205263|Induce (action)|inducible
Event|Event|Hospital Course|3288,3296|false|false|false|||ischemia
Finding|Pathologic Function|Hospital Course|3288,3296|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3288,3296|false|false|false|C4321499|Ischemia Procedure|ischemia
Event|Event|Hospital Course|3297,3301|false|false|false|||seen
Event|Event|Hospital Course|3306,3310|false|false|false|||ECHO
Procedure|Health Care Activity|Hospital Course|3306,3310|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3306,3310|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|Hospital Course|3311,3317|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|3311,3317|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|3311,3317|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|3311,3317|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|3311,3322|false|false|false|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Hospital Course|3318,3322|false|false|false|C4318744|Test - temporal region|test
Event|Event|Hospital Course|3318,3322|false|false|false|||test
Finding|Functional Concept|Hospital Course|3318,3322|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Hospital Course|3318,3322|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Hospital Course|3318,3322|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Hospital Course|3318,3322|false|false|false|C0022885|Laboratory Procedures|test
Finding|Finding|Hospital Course|3338,3342|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|3338,3342|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|3338,3342|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|3346,3355|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|3346,3355|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|3362,3370|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|3362,3370|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|3362,3370|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|3375,3383|false|false|false|||resolved
Disorder|Congenital Abnormality|Hospital Course|3388,3401|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Hospital Course|3388,3401|false|false|false|||abnormalities
Finding|Functional Concept|Hospital Course|3388,3401|true|false|false|C0000769|teratologic|abnormalities
Event|Event|Hospital Course|3407,3411|false|false|false|||seen
Event|Event|Hospital Course|3415,3422|false|false|false|||imaging
Finding|Finding|Hospital Course|3415,3422|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|3415,3422|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Event|Event|Hospital Course|3427,3431|false|false|false|||labs
Lab|Laboratory or Test Result|Hospital Course|3427,3431|false|false|false|C0587081|Laboratory test finding|labs
Finding|Gene or Genome|Hospital Course|3448,3451|false|false|false|C1418526;C5891011|PHEX gene;PHEX wt Allele|PEx
Event|Event|Hospital Course|3457,3467|false|false|false|||remarkable
Anatomy|Body Location or Region|Hospital Course|3487,3491|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3487,3491|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|3487,3491|false|false|false|C0024115|Lung diseases|lung
Event|Event|Hospital Course|3487,3491|false|false|false|||lung
Finding|Finding|Hospital Course|3487,3491|false|false|false|C0740941|Lung Problem|lung
Event|Event|Findings|3511,3516|false|false|false|||ruled
Finding|Classification|Findings|3529,3537|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Findings|3529,3537|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Findings|3529,3537|false|false|false|C5237010|Expression Negative|negative
Event|Event|Findings|3545,3548|false|false|false|||EKG
Finding|Intellectual Product|Findings|3545,3548|true|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|Findings|3545,3548|true|false|false|C1623258|Electrocardiography|EKG
Event|Event|Findings|3549,3556|false|false|false|||changes
Finding|Functional Concept|Findings|3549,3556|true|false|false|C0392747|Changing|changes
Anatomy|Body System|Findings|3560,3570|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Event|Findings|3575,3584|false|false|false|||consulted
Event|Event|Findings|3588,3596|false|false|false|||evaluate
Event|Event|Findings|3597,3601|false|false|false|||need
Finding|Functional Concept|Findings|3597,3601|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Findings|3597,3605|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|Findings|3606,3621|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Findings|3606,3621|false|false|false|C0007430|Catheterization|catheterization
Event|Event|Findings|3632,3644|false|false|false|||intervention
Procedure|Health Care Activity|Findings|3632,3644|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Findings|3632,3644|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Event|Event|Findings|3658,3662|false|false|false|||feel
Event|Event|Findings|3672,3678|false|false|false|||urgent
Finding|Intellectual Product|Findings|3672,3678|true|false|false|C1546403;C1546845;C1547230;C1561556|Admission Type - Urgent;Certification patient type - Urgent;Triage Code - Urgent;Visit Priority Code - Urgent|urgent
Event|Event|Findings|3680,3689|false|false|false|||inpatient
Finding|Idea or Concept|Findings|3680,3689|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Findings|3680,3689|false|false|false|C1555324|inpatient encounter|inpatient
Event|Occupational Activity|Findings|3690,3694|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Findings|3690,3697|false|false|false|C0750430|Work-up|work-up
Event|Event|Findings|3702,3711|false|false|false|||necessary
Finding|Idea or Concept|Findings|3731,3738|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Intellectual Product|Findings|3731,3738|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Mental Process|Findings|3731,3738|false|false|false|C0449255;C0542559;C4281677|Application Context;Context;contextual factors|context
Finding|Finding|Findings|3743,3755|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|Findings|3756,3767|false|false|false|||tachycardia
Finding|Finding|Findings|3756,3767|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|tachycardia
Event|Event|Findings|3801,3805|false|false|false|||ECHO
Procedure|Health Care Activity|Findings|3801,3805|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Findings|3801,3805|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Event|Event|Findings|3821,3830|false|false|false|||admission
Procedure|Health Care Activity|Findings|3821,3830|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Anatomy|Body System|Findings|3833,3843|false|false|false|C0007226|Cardiovascular system|Cardiology
Event|Event|Findings|3844,3855|false|false|false|||recommended
Event|Event|Findings|3856,3866|false|false|false|||restarting
Drug|Organic Chemical|Findings|3868,3880|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Findings|3868,3880|false|false|false|C0039771|theophylline|theophylline
Event|Event|Findings|3868,3880|false|false|false|||theophylline
Procedure|Laboratory Procedure|Findings|3868,3880|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Amino Acid, Peptide, or Protein|Findings|3888,3892|false|false|false|C5552605|FACT Complex|fact
Drug|Biologically Active Substance|Findings|3888,3892|false|false|false|C5552605|FACT Complex|fact
Event|Event|Findings|3888,3892|false|false|false|||fact
Finding|Gene or Genome|Findings|3888,3892|false|false|false|C1420522;C5551287|SSRP1 wt Allele;SUPT16H gene|fact
Event|Event|Findings|3898,3906|false|false|false|||received
Event|Event|Findings|3912,3919|false|false|false|||benefit
Anatomy|Body Part, Organ, or Organ Component|Findings|3926,3935|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Findings|3926,3935|false|false|false|C2707265||pulmonary
Finding|Finding|Findings|3926,3935|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Findings|3960,3969|false|false|false|||restarted
Drug|Organic Chemical|Findings|3973,3985|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Findings|3973,3985|false|false|false|C0039771|theophylline|theophylline
Event|Event|Findings|3973,3985|false|false|false|||theophylline
Procedure|Laboratory Procedure|Findings|3973,3985|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Findings|3993,3996|false|false|false|||TID
Event|Event|Findings|4012,4016|false|false|false|||dose
Event|Event|Findings|4026,4041|false|false|false|||discontinuation
Finding|Finding|Findings|4026,4041|false|false|false|C0457454;C1444662|Discontinuation (procedure);Discontinued|discontinuation
Finding|Functional Concept|Findings|4026,4041|false|false|false|C0457454;C1444662|Discontinuation (procedure);Discontinued|discontinuation
Drug|Hazardous or Poisonous Substance|Findings|4058,4065|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Immunologic Factor|Findings|4058,4065|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Organic Chemical|Findings|4058,4065|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Drug|Pharmacologic Substance|Findings|4058,4065|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|tobacco
Finding|Individual Behavior|Findings|4058,4075|false|false|false|C0600549|Tobacco Use Cessation|tobacco cessation
Event|Activity|Findings|4066,4075|false|false|false|C1880019|Cessation|cessation
Event|Event|Findings|4076,4085|false|false|false|||education
Finding|Classification|Findings|4076,4085|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Finding|Finding|Findings|4076,4085|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Procedure|Educational Activity|Findings|4076,4085|false|false|false|C0013621;C0039401|Education (procedure);Knowledge acquisition|education
Event|Event|Findings|4091,4100|false|false|false|||continued
Event|Event|Findings|4104,4108|false|false|false|||home
Finding|Idea or Concept|Findings|4104,4108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Findings|4104,4108|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Findings|4104,4108|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Findings|4110,4119|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Findings|4110,4119|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Findings|4110,4119|false|false|false|||diltiazem
Drug|Organic Chemical|Findings|4124,4131|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Findings|4124,4131|false|false|false|C0004057|aspirin|aspirin
Event|Event|Findings|4124,4131|false|false|false|||aspirin
Event|Event|Findings|4133,4137|false|false|false|||dose
Event|Event|Findings|4154,4163|false|false|false|||increased
Event|Event|Findings|4183,4189|false|false|false|||ruling
Procedure|Health Care Activity|Findings|4200,4209|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|Findings|4233,4240|false|false|false|||pending
Finding|Idea or Concept|Findings|4233,4240|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|Findings|4248,4252|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Findings|4248,4252|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Findings|4248,4252|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Findings|4256,4265|false|false|false|||discharge
Finding|Body Substance|Findings|4256,4265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Findings|4256,4265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Findings|4256,4265|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Findings|4256,4265|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Findings|4273,4279|false|false|false|C0004096|Asthma|Asthma
Event|Event|Findings|4273,4279|false|false|false|||Asthma
Disorder|Disease or Syndrome|Findings|4284,4288|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Findings|4284,4288|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Findings|4284,4288|false|false|false|||COPD
Finding|Gene or Genome|Findings|4284,4288|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Body Substance|Findings|4290,4297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Findings|4290,4297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Findings|4290,4297|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Findings|4302,4307|false|false|false|||given
Drug|Organic Chemical|Findings|4308,4317|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Findings|4308,4317|false|false|false|C0001927|albuterol|Albuterol
Event|Event|Findings|4308,4317|false|false|false|||Albuterol
Drug|Organic Chemical|Findings|4322,4333|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|Findings|4322,4333|false|false|false|C0027235|ipratropium|ipratropium
Event|Event|Findings|4322,4333|false|false|false|||ipratropium
Drug|Biomedical or Dental Material|Findings|4335,4339|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|Findings|4335,4339|false|false|false|||nebs
Event|Event|Findings|4353,4362|false|false|false|||continued
Finding|Idea or Concept|Findings|4370,4374|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Findings|4370,4374|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Findings|4370,4374|false|false|false|C1553498|home health encounter|home
Event|Event|Findings|4375,4380|false|false|false|||doses
Drug|Organic Chemical|Findings|4384,4395|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|4384,4395|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Findings|4384,4395|false|false|false|||fluticasone
Drug|Organic Chemical|Findings|4398,4409|false|false|false|C0298130|montelukast|montelukast
Drug|Pharmacologic Substance|Findings|4398,4409|false|false|false|C0298130|montelukast|montelukast
Event|Event|Findings|4398,4409|false|false|false|||montelukast
Drug|Organic Chemical|Findings|4411,4422|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|4411,4422|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Findings|4411,4422|false|false|false|||fluticasone
Event|Event|Findings|4423,4432|false|false|false|||salmetrol
Event|Event|Findings|4452,4455|false|false|false|||PRN
Finding|Gene or Genome|Findings|4452,4455|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body System|Findings|4465,4475|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Findings|4476,4483|false|false|false|||consult
Procedure|Health Care Activity|Findings|4476,4483|false|false|false|C0009818|Consultation|consult
Event|Event|Findings|4493,4502|false|false|false|||restarted
Drug|Organic Chemical|Findings|4510,4522|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Findings|4510,4522|false|false|false|C0039771|theophylline|theophylline
Event|Event|Findings|4510,4522|false|false|false|||theophylline
Procedure|Laboratory Procedure|Findings|4510,4522|false|false|false|C0039773|Assay of theophylline|theophylline
Event|Event|Findings|4533,4536|false|false|false|||TID
Event|Event|Findings|4543,4547|false|false|false|||pulm
Procedure|Health Care Activity|Findings|4543,4547|false|false|false|C1315068|Pulmonary ventilator management|pulm
Anatomy|Body System|Findings|4552,4562|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Findings|4563,4569|false|false|false|||follow
Finding|Functional Concept|Findings|4563,4569|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Findings|4563,4569|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Findings|4563,4572|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Findings|4563,4572|false|false|false|C1522577|follow-up|follow-up
Event|Event|Findings|4570,4572|false|false|false|||up
Drug|Hazardous or Poisonous Substance|Findings|4580,4587|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|Findings|4580,4587|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|Findings|4580,4587|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|Findings|4580,4587|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Disorder|Mental or Behavioral Dysfunction|Findings|4580,4593|false|false|false|C0040336|Tobacco Use Disorder|Tobacco abuse
Disorder|Mental or Behavioral Dysfunction|Findings|4588,4593|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Findings|4588,4593|false|false|false|||abuse
Event|Event|Findings|4588,4593|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Findings|4588,4593|false|false|false|C0562381|Victim of abuse (finding)|abuse
Event|Event|Findings|4599,4607|false|false|false|||declined
Drug|Hazardous or Poisonous Substance|Findings|4608,4616|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|Findings|4608,4616|false|false|false|C0028040|nicotine|nicotine
Drug|Clinical Drug|Findings|4608,4622|false|false|false|C0358855|Nicotine Transdermal Patch|nicotine patch
Drug|Biomedical or Dental Material|Findings|4617,4622|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Event|Event|Findings|4617,4622|false|false|false|||patch
Finding|Finding|Findings|4617,4622|false|false|false|C0332461|Plaque (lesion)|patch
Event|Event|Findings|4628,4637|false|false|false|||education
Finding|Classification|Findings|4628,4637|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Finding|Finding|Findings|4628,4637|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Procedure|Educational Activity|Findings|4628,4637|false|false|false|C0013621;C0039401|Education (procedure);Knowledge acquisition|education
Finding|Idea or Concept|Findings|4663,4669|false|false|false|C0018684|Health|health
Drug|Hazardous or Poisonous Substance|Findings|4663,4677|false|false|false|C0079483|health hazards|health hazards
Event|Event|Findings|4670,4677|false|false|false|||hazards
Event|Event|Findings|4681,4688|false|false|false|||smoking
Finding|Individual Behavior|Findings|4681,4688|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|Findings|4681,4688|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Body Substance|Findings|4700,4707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Findings|4700,4707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Findings|4700,4707|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Findings|4712,4721|false|false|false|||continued
Drug|Organic Chemical|Findings|4729,4740|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Findings|4729,4740|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Findings|4729,4740|false|false|false|||simvastatin
Drug|Biologically Active Substance|Findings|4759,4762|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Findings|4759,4762|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Findings|4759,4762|false|false|false|||LDL
Procedure|Laboratory Procedure|Findings|4759,4762|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Idea or Concept|Findings|4774,4778|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Findings|4774,4778|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|Findings|4790,4794|false|false|false|||dose
Event|Event|Findings|4799,4808|false|false|false|||increased
Finding|Finding|Findings|4826,4834|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|INACTIVE
Finding|Idea or Concept|Findings|4826,4834|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|INACTIVE
Event|Event|Findings|4835,4841|false|false|false|||ISSUES
Disorder|Disease or Syndrome|Findings|4847,4850|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Findings|4847,4850|false|false|false|||HTN
Finding|Idea or Concept|Findings|4852,4861|false|false|false|C0549178|Continuous|continued
Drug|Organic Chemical|Findings|4862,4872|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Findings|4862,4872|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|Findings|4862,4872|false|false|false|||isosorbide
Drug|Organic Chemical|Findings|4877,4896|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Findings|4877,4896|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Findings|4877,4896|false|false|false|||hydrochlorothiazide
Finding|Finding|Findings|4897,4904|false|false|false|C4534363|At home|at home
Event|Event|Findings|4900,4904|false|false|false|||home
Finding|Idea or Concept|Findings|4900,4904|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Findings|4900,4904|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Findings|4900,4904|false|false|false|C1553498|home health encounter|home
Event|Event|Findings|4906,4911|false|false|false|||doses
Event|Event|Findings|4917,4921|false|false|false|||Code
Event|Occupational Activity|Findings|4917,4921|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Findings|4917,4921|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Attribute|Clinical Attribute|Findings|4930,4941|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Findings|4930,4941|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Findings|4930,4941|false|false|false|||Medications
Finding|Intellectual Product|Findings|4930,4941|false|false|false|C4284232|Medications|Medications
Finding|Finding|Findings|4930,4954|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Findings|4945,4954|false|false|false|||Admission
Procedure|Health Care Activity|Findings|4945,4954|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|Findings|4957,4970|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Findings|4957,4970|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Findings|4957,4970|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Findings|4957,4970|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Findings|4978,4984|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Findings|4998,5004|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|5033,5039|false|false|false|||needed
Attribute|Clinical Attribute|Findings|5044,5048|false|false|false|C2598155||pain
Event|Event|Findings|5044,5048|false|false|false|||pain
Finding|Functional Concept|Findings|5044,5048|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Findings|5044,5048|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Findings|5053,5062|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Findings|5053,5062|false|false|false|C0001927|albuterol|albuterol
Event|Event|Findings|5053,5062|false|false|false|||albuterol
Drug|Organic Chemical|Findings|5053,5070|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Findings|5053,5070|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Findings|5063,5070|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Findings|5063,5070|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Findings|5063,5070|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Findings|5063,5070|false|false|false|||sulfate
Disorder|Disease or Syndrome|Findings|5088,5091|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Findings|5088,5091|false|false|false|||HFA
Procedure|Diagnostic Procedure|Findings|5088,5091|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Findings|5092,5099|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|Findings|5100,5107|false|false|false|||Inhaler
Finding|Functional Concept|Findings|5100,5107|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Finding|Functional Concept|Findings|5123,5133|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|5123,5133|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Drug|Organic Chemical|Findings|5154,5163|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Findings|5154,5163|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Findings|5154,5163|false|false|false|||diltiazem
Drug|Organic Chemical|Findings|5154,5167|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Findings|5154,5167|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Findings|5164,5167|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Findings|5164,5167|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Findings|5164,5167|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Findings|5164,5167|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Findings|5164,5167|false|false|false|||HCl
Anatomy|Body Part, Organ, or Organ Component|Findings|5175,5182|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5175,5182|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5175,5182|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|5175,5200|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Findings|5184,5192|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|5184,5192|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|5193,5200|false|false|false|||Release
Finding|Functional Concept|Findings|5193,5200|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5193,5200|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5193,5200|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Findings|5215,5222|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5215,5222|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5215,5222|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|5215,5240|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Findings|5224,5232|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|5224,5232|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|5233,5240|false|false|false|||Release
Finding|Functional Concept|Findings|5233,5240|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5233,5240|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5233,5240|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|5262,5273|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|5262,5273|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Findings|5262,5273|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|Findings|5291,5296|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Findings|5291,5296|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Findings|5291,5296|false|false|false|||Spray
Finding|Functional Concept|Findings|5291,5296|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Findings|5291,5308|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Findings|5298,5308|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Findings|5298,5308|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|Findings|5298,5308|false|false|false|||Suspension
Finding|Functional Concept|Findings|5298,5308|false|false|false|C1705537|Suspension (action)|Suspension
Drug|Biomedical or Dental Material|Findings|5323,5328|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Findings|5323,5328|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Findings|5323,5328|false|false|false|||Spray
Finding|Functional Concept|Findings|5323,5328|false|false|false|C4521772|Spray (administration method)|Spray
Anatomy|Body Part, Organ, or Organ Component|Findings|5329,5334|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Findings|5329,5334|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Findings|5329,5334|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Findings|5329,5334|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Findings|5329,5334|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Findings|5329,5334|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Findings|5335,5340|false|false|false|||DAILY
Drug|Organic Chemical|Findings|5353,5364|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|5353,5364|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|5353,5375|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Findings|5365,5375|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Findings|5365,5375|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|Findings|5365,5375|false|false|false|||salmeterol
Anatomy|Body Part, Organ, or Organ Component|Findings|5392,5396|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Findings|5392,5396|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Findings|5402,5408|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Findings|5409,5412|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Findings|5409,5412|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Findings|5409,5412|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Findings|5409,5412|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|5423,5427|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Findings|5423,5427|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Findings|5433,5439|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Findings|5440,5450|false|false|false|||Inhalation
Finding|Functional Concept|Findings|5440,5450|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|5440,5450|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Findings|5451,5454|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Findings|5451,5454|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Findings|5451,5454|false|false|false|C1530795|BID protein, human|BID
Event|Event|Findings|5451,5454|false|false|false|||BID
Finding|Gene or Genome|Findings|5451,5454|false|false|false|C1332410|BID gene|BID
Finding|Finding|Findings|5456,5463|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Findings|5458,5463|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Findings|5466,5469|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|5466,5469|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Findings|5475,5494|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Findings|5475,5494|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Findings|5475,5494|false|false|false|||hydrochlorothiazide
Anatomy|Body Part, Organ, or Organ Component|Findings|5503,5510|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5503,5510|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5503,5510|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Findings|5511,5514|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|5524,5531|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5524,5531|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5524,5531|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|Findings|5554,5564|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Findings|5554,5564|false|false|false|C0022251|isosorbide|isosorbide
Drug|Organic Chemical|Findings|5554,5576|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|Findings|5554,5576|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|Findings|5565,5576|false|false|false|||mononitrate
Drug|Biomedical or Dental Material|Findings|5583,5589|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Findings|5590,5598|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|5590,5598|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|5599,5606|false|false|false|||Release
Finding|Functional Concept|Findings|5599,5606|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5599,5606|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5599,5606|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Findings|5614,5617|false|false|false|||Sig
Drug|Biomedical or Dental Material|Findings|5627,5633|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Findings|5634,5642|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|5634,5642|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|5643,5650|false|false|false|||Release
Finding|Functional Concept|Findings|5643,5650|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5643,5650|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5643,5650|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|5678,5689|false|false|false|C0298130|montelukast|montelukast
Drug|Pharmacologic Substance|Findings|5678,5689|false|false|false|C0298130|montelukast|montelukast
Event|Event|Findings|5678,5689|false|false|false|||montelukast
Drug|Biomedical or Dental Material|Findings|5696,5702|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Findings|5716,5722|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|5716,5722|false|false|false|||Tablet
Drug|Organic Chemical|Findings|5745,5755|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Findings|5745,5755|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Findings|5745,5755|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Findings|5762,5769|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5762,5769|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5762,5769|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Findings|5771,5778|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Findings|5771,5786|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Findings|5779,5786|false|false|false|||Release
Finding|Functional Concept|Findings|5779,5786|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5779,5786|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5779,5786|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Findings|5793,5796|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|5807,5814|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5807,5814|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5807,5814|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Findings|5816,5823|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Findings|5816,5831|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Findings|5824,5831|false|false|false|||Release
Finding|Functional Concept|Findings|5824,5831|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|5824,5831|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|5824,5831|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|5859,5869|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|Findings|5859,5869|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|Findings|5859,5869|false|false|false|||tiotropium
Drug|Organic Chemical|Findings|5859,5877|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Pharmacologic Substance|Findings|5859,5877|false|false|false|C1306772|tiotropium bromide|tiotropium bromide
Drug|Inorganic Chemical|Findings|5870,5877|false|false|false|C0006222|Bromides|bromide
Event|Event|Findings|5870,5877|false|false|false|||bromide
Procedure|Laboratory Procedure|Findings|5870,5877|false|false|false|C0202341|Bromides measurement|bromide
Anatomy|Body Part, Organ, or Organ Component|Findings|5885,5892|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|5885,5892|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|5885,5892|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Findings|5896,5906|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|5896,5906|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Functional Concept|Findings|5907,5913|false|false|false|C1550509|Participation Type - device|Device
Disorder|Congenital Abnormality|Findings|5928,5931|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|Cap
Drug|Biomedical or Dental Material|Findings|5928,5931|false|false|false|C0006935|capsule (pharmacologic)|Cap
Event|Event|Findings|5928,5931|false|false|false|||Cap
Finding|Gene or Genome|Findings|5928,5931|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|Cap
Procedure|Therapeutic or Preventive Procedure|Findings|5928,5931|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|Cap
Finding|Functional Concept|Findings|5932,5942|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|5932,5942|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Findings|5943,5948|false|false|false|||DAILY
Drug|Biologically Active Substance|Findings|5961,5968|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Findings|5961,5968|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Findings|5961,5968|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Findings|5961,5968|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Findings|5961,5968|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Findings|5961,5968|false|false|false|||calcium
Finding|Physiologic Function|Findings|5961,5968|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Findings|5961,5968|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Findings|5961,5978|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Findings|5961,5978|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Findings|5969,5978|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Findings|5969,5978|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Findings|5969,5978|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Findings|5969,5978|false|false|false|||carbonate
Drug|Biomedical or Dental Material|Findings|5995,6001|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|5995,6001|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|5995,6011|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Findings|6012,6015|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Findings|6012,6015|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Findings|6012,6015|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Findings|6012,6015|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Findings|6026,6032|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6026,6032|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|6026,6042|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Organic Chemical|Findings|6064,6076|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Findings|6064,6076|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Findings|6064,6076|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Findings|6064,6087|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Findings|6081,6087|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6081,6087|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|6101,6107|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6101,6107|false|false|false|||Tablet
Drug|Organic Chemical|Findings|6130,6137|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Findings|6130,6137|false|false|false|C0004057|aspirin|aspirin
Event|Event|Findings|6130,6137|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Findings|6144,6150|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6151,6154|false|false|false|||Sig
Drug|Biomedical or Dental Material|Findings|6164,6170|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6164,6170|false|false|false|||Tablet
Event|Event|Findings|6171,6173|false|false|false|||PO
Finding|Intellectual Product|Findings|6174,6178|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Findings|6174,6184|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Findings|6181,6184|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|6181,6184|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Findings|6189,6200|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Findings|6189,6200|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Findings|6213,6222|false|false|false|||Discharge
Finding|Body Substance|Findings|6213,6222|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Findings|6213,6222|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Findings|6213,6222|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Findings|6213,6222|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Findings|6213,6234|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Findings|6223,6234|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Findings|6223,6234|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Findings|6223,6234|false|false|false|||Medications
Finding|Intellectual Product|Findings|6223,6234|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Findings|6239,6250|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Findings|6239,6250|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Findings|6239,6250|false|false|false|||simvastatin
Drug|Biomedical or Dental Material|Findings|6257,6263|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Findings|6277,6283|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6277,6283|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|6312,6318|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Findings|6323,6330|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Findings|6338,6357|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Findings|6338,6357|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Findings|6338,6357|false|false|false|||hydrochlorothiazide
Anatomy|Body Part, Organ, or Organ Component|Findings|6366,6373|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|6366,6373|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|6366,6373|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Event|Event|Findings|6374,6377|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|6387,6394|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|6387,6394|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|6387,6394|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Organic Chemical|Findings|6419,6430|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|6419,6430|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Findings|6419,6430|false|false|false|||fluticasone
Drug|Biomedical or Dental Material|Findings|6448,6453|false|false|false|C1154182|Spray Dosage Form|Spray
Event|Activity|Findings|6448,6453|false|false|false|C2003858|Spray (action)|Spray
Event|Event|Findings|6448,6453|false|false|false|||Spray
Finding|Functional Concept|Findings|6448,6453|false|false|false|C4521772|Spray (administration method)|Spray
Drug|Biomedical or Dental Material|Findings|6448,6465|false|false|false|C1710170|SPRAY, SUSPENSION|Spray, Suspension
Drug|Biomedical or Dental Material|Findings|6455,6465|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Drug|Substance|Findings|6455,6465|false|false|false|C0038960;C1382107|Suspension substance;Suspensions|Suspension
Event|Event|Findings|6455,6465|false|false|false|||Suspension
Finding|Functional Concept|Findings|6455,6465|false|false|false|C1705537|Suspension (action)|Suspension
Disorder|Mental or Behavioral Dysfunction|Findings|6476,6482|false|false|false|C0233601|Spraying behavior|Sprays
Drug|Biomedical or Dental Material|Findings|6476,6482|false|false|false|C1154182|Spray Dosage Form|Sprays
Event|Event|Findings|6476,6482|false|false|false|||Sprays
Anatomy|Body Part, Organ, or Organ Component|Findings|6483,6488|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Findings|6483,6488|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Findings|6483,6488|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Findings|6483,6488|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Findings|6483,6488|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Findings|6483,6488|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Event|Event|Findings|6489,6494|false|false|false|||DAILY
Event|Event|Findings|6506,6512|false|false|false|||needed
Event|Event|Findings|6517,6527|false|false|false|||congestion
Finding|Pathologic Function|Findings|6517,6527|false|false|false|C0700148|Congestion|congestion
Drug|Organic Chemical|Findings|6534,6544|false|false|false|C0022251|isosorbide|isosorbide
Drug|Pharmacologic Substance|Findings|6534,6544|false|false|false|C0022251|isosorbide|isosorbide
Event|Event|Findings|6534,6544|false|false|false|||isosorbide
Drug|Organic Chemical|Findings|6534,6556|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Drug|Pharmacologic Substance|Findings|6534,6556|false|false|false|C0064079|isosorbide mononitrate|isosorbide mononitrate
Event|Event|Findings|6545,6556|false|false|false|||mononitrate
Drug|Biomedical or Dental Material|Findings|6563,6569|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Findings|6570,6578|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|6570,6578|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|6579,6586|false|false|false|||Release
Finding|Functional Concept|Findings|6579,6586|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|6579,6586|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|6579,6586|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Findings|6594,6597|false|false|false|||Sig
Drug|Biomedical or Dental Material|Findings|6607,6613|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Finding|Findings|6614,6622|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|6614,6622|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|6623,6630|false|false|false|||Release
Finding|Functional Concept|Findings|6623,6630|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|6623,6630|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|6623,6630|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|6660,6671|false|false|false|C0298130|montelukast|montelukast
Drug|Pharmacologic Substance|Findings|6660,6671|false|false|false|C0298130|montelukast|montelukast
Event|Event|Findings|6660,6671|false|false|false|||montelukast
Drug|Biomedical or Dental Material|Findings|6678,6684|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Findings|6698,6704|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6698,6704|false|false|false|||Tablet
Drug|Organic Chemical|Findings|6729,6740|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Findings|6729,6740|false|false|false|C0082607|fluticasone|fluticasone
Event|Event|Findings|6729,6740|false|false|false|||fluticasone
Drug|Pharmacologic Substance|Findings|6729,6751|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Findings|6741,6751|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Findings|6741,6751|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|Findings|6741,6751|false|false|false|||salmeterol
Anatomy|Body Part, Organ, or Organ Component|Findings|6768,6772|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Findings|6768,6772|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Findings|6778,6784|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Findings|6785,6788|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Findings|6785,6788|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Findings|6785,6788|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Findings|6785,6788|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|6799,6803|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Findings|6799,6803|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Findings|6809,6815|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Findings|6816,6826|false|false|false|||Inhalation
Finding|Functional Concept|Findings|6816,6826|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|6816,6826|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Findings|6827,6830|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Findings|6827,6830|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Findings|6827,6830|false|false|false|C1530795|BID protein, human|BID
Event|Event|Findings|6827,6830|false|false|false|||BID
Finding|Gene or Genome|Findings|6827,6830|false|false|false|C1332410|BID gene|BID
Finding|Finding|Findings|6832,6839|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Findings|6834,6839|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Findings|6842,6845|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|6842,6845|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Findings|6853,6866|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Findings|6853,6866|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Findings|6853,6866|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Findings|6853,6866|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Pharmacologic Substance|Findings|6853,6874|false|false|false|C2351132|Acetaminophen / Codeine|acetaminophen-codeine
Drug|Organic Chemical|Findings|6867,6874|false|false|false|C0009214|codeine|codeine
Drug|Pharmacologic Substance|Findings|6867,6874|false|false|false|C0009214|codeine|codeine
Event|Event|Findings|6867,6874|false|false|false|||codeine
Drug|Biomedical or Dental Material|Findings|6885,6891|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6892,6895|false|false|false|||Sig
Drug|Biomedical or Dental Material|Findings|6905,6911|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|6940,6946|false|false|false|||needed
Attribute|Clinical Attribute|Findings|6951,6955|false|false|false|C2598155||pain
Event|Event|Findings|6951,6955|false|false|false|||pain
Finding|Functional Concept|Findings|6951,6955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Findings|6951,6955|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Findings|6962,6971|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Findings|6962,6971|false|false|false|C0001927|albuterol|albuterol
Event|Event|Findings|6962,6971|false|false|false|||albuterol
Drug|Organic Chemical|Findings|6962,6979|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Findings|6962,6979|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Findings|6972,6979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Findings|6972,6979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Findings|6972,6979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Findings|6972,6979|false|false|false|||sulfate
Disorder|Disease or Syndrome|Findings|6997,7000|false|false|false|C0015458|Facial Hemiatrophy|HFA
Event|Event|Findings|6997,7000|false|false|false|||HFA
Procedure|Diagnostic Procedure|Findings|6997,7000|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Biomedical or Dental Material|Findings|7001,7008|false|false|false|C1112870|Aerosol Dose Form|Aerosol
Event|Event|Findings|7009,7016|false|false|false|||Inhaler
Finding|Functional Concept|Findings|7009,7016|false|false|false|C4319647|Inhaler (unit of presentation)|Inhaler
Event|Event|Findings|7037,7047|false|false|false|||Inhalation
Finding|Functional Concept|Findings|7037,7047|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|7037,7047|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Findings|7067,7073|false|false|false|||needed
Event|Event|Findings|7078,7087|false|false|false|||shortness
Finding|Body Substance|Findings|7092,7098|false|false|false|C0225386|Breath|breath
Event|Event|Findings|7102,7110|false|false|false|||wheezing
Finding|Sign or Symptom|Findings|7102,7110|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|Findings|7117,7127|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Findings|7117,7127|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Findings|7117,7127|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Findings|7134,7141|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7134,7141|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7134,7141|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Findings|7143,7150|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Findings|7143,7158|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Findings|7151,7158|false|false|false|||Release
Finding|Functional Concept|Findings|7151,7158|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7151,7158|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7151,7158|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Findings|7165,7168|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|7179,7186|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7179,7186|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7179,7186|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Findings|7188,7195|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Findings|7188,7203|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Findings|7196,7203|false|false|false|||Release
Finding|Functional Concept|Findings|7196,7203|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7196,7203|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7196,7203|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|7234,7241|false|false|false|C0905678|Spiriva|Spiriva
Drug|Pharmacologic Substance|Findings|7234,7241|false|false|false|C0905678|Spiriva|Spiriva
Event|Event|Findings|7234,7241|false|false|false|||Spiriva
Anatomy|Body Part, Organ, or Organ Component|Findings|7265,7272|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7265,7272|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7265,7272|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Functional Concept|Findings|7276,7286|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|7276,7286|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Findings|7287,7293|false|false|false|||Device
Finding|Functional Concept|Findings|7287,7293|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Findings|7295,7298|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Findings|7308,7315|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Findings|7308,7315|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Findings|7308,7315|false|false|false|C0006935|capsule (pharmacologic)|capsule
Event|Event|Findings|7316,7326|false|false|false|||Inhalation
Finding|Functional Concept|Findings|7316,7326|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|7316,7326|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Intellectual Product|Findings|7327,7331|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Findings|7327,7337|false|false|false|C3537736|Once A Day|once a day
Event|Event|Findings|7334,7337|false|false|false|||day
Finding|Idea or Concept|Findings|7334,7337|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|7334,7337|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Findings|7345,7352|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Findings|7345,7352|false|false|false|C0004057|aspirin|aspirin
Event|Event|Findings|7345,7352|false|false|false|||aspirin
Drug|Biomedical or Dental Material|Findings|7359,7365|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7366,7369|false|false|false|||Sig
Drug|Biomedical or Dental Material|Findings|7379,7385|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7379,7385|false|false|false|||Tablet
Event|Event|Findings|7386,7388|false|false|false|||PO
Finding|Intellectual Product|Findings|7389,7393|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Pharmacologic Substance|Findings|7389,7399|false|false|false|C3537736|Once A Day|once a day
Finding|Idea or Concept|Findings|7396,7399|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|7396,7399|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biologically Active Substance|Findings|7407,7414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Findings|7407,7414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Findings|7407,7414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Findings|7407,7414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Findings|7407,7414|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Findings|7407,7414|false|false|false|||calcium
Finding|Physiologic Function|Findings|7407,7414|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Findings|7407,7414|false|false|false|C0201925|Calcium measurement|calcium
Drug|Inorganic Chemical|Findings|7407,7424|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Pharmacologic Substance|Findings|7407,7424|false|false|false|C0006681|calcium carbonate|calcium carbonate
Drug|Element, Ion, or Isotope|Findings|7415,7424|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Organic Chemical|Findings|7415,7424|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Drug|Pharmacologic Substance|Findings|7415,7424|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|carbonate
Event|Event|Findings|7415,7424|false|false|false|||carbonate
Drug|Biomedical or Dental Material|Findings|7441,7447|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7441,7447|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|7441,7457|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Anatomy|Body Part, Organ, or Organ Component|Findings|7458,7461|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Findings|7458,7461|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Findings|7458,7461|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Findings|7458,7461|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Biomedical or Dental Material|Findings|7472,7478|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7472,7478|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|7472,7488|false|false|false|C0304290|Chewable Tablet|Tablet, Chewable
Drug|Organic Chemical|Findings|7513,7522|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Findings|7513,7522|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Findings|7513,7522|false|false|false|||diltiazem
Drug|Organic Chemical|Findings|7513,7526|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Drug|Pharmacologic Substance|Findings|7513,7526|false|false|false|C0700579|diltiazem hydrochloride|diltiazem HCl
Disorder|Neoplastic Process|Findings|7523,7526|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|Findings|7523,7526|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|Findings|7523,7526|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|Findings|7523,7526|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|Findings|7523,7526|false|false|false|||HCl
Anatomy|Body Part, Organ, or Organ Component|Findings|7534,7541|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7534,7541|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7534,7541|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|7534,7559|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Findings|7543,7551|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|7543,7551|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|7552,7559|false|false|false|||Release
Finding|Functional Concept|Findings|7552,7559|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7552,7559|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7552,7559|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Findings|7574,7581|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7574,7581|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7574,7581|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|7574,7599|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Findings|7583,7591|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Findings|7583,7591|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Findings|7592,7599|false|false|false|||Release
Finding|Functional Concept|Findings|7592,7599|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7592,7599|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7592,7599|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Findings|7624,7636|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Findings|7624,7636|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Vitamin|Findings|7624,7636|false|false|false|C0301532|Multivitamin preparation|multivitamin
Drug|Pharmacologic Substance|Findings|7624,7647|false|false|false|C0978787|Multivitamin tablet|multivitamin     Tablet
Drug|Biomedical or Dental Material|Findings|7641,7647|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7641,7647|false|false|false|||Tablet
Drug|Biomedical or Dental Material|Findings|7661,7667|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Findings|7661,7667|false|false|false|||Tablet
Drug|Organic Chemical|Findings|7693,7705|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Findings|7693,7705|false|false|false|C0039771|theophylline|theophylline
Event|Event|Findings|7693,7705|false|false|false|||theophylline
Procedure|Laboratory Procedure|Findings|7693,7705|false|false|false|C0039773|Assay of theophylline|theophylline
Anatomy|Body Part, Organ, or Organ Component|Findings|7713,7720|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7713,7720|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7713,7720|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|7713,7739|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Findings|7722,7725|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|Findings|7722,7725|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Findings|7726,7733|false|false|false|||Release
Finding|Functional Concept|Findings|7726,7733|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7726,7733|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7726,7733|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Findings|7754,7761|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7754,7761|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7754,7761|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|7754,7780|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Findings|7763,7766|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Findings|7763,7766|false|false|false|||Ext
Finding|Gene or Genome|Findings|7763,7766|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Findings|7767,7774|false|false|false|||Release
Finding|Functional Concept|Findings|7767,7774|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7767,7774|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7767,7774|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Disease or Syndrome|Findings|7790,7795|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Findings|7798,7801|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Findings|7798,7801|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Anatomy|Body Part, Organ, or Organ Component|Findings|7812,7819|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Findings|7812,7819|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Findings|7812,7819|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Findings|7812,7838|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Findings|7821,7824|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Findings|7821,7824|false|false|false|||Ext
Finding|Gene or Genome|Findings|7821,7824|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Findings|7825,7832|false|false|false|||Release
Finding|Functional Concept|Findings|7825,7832|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Findings|7825,7832|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Findings|7825,7832|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Idea or Concept|Findings|7843,7850|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Findings|7859,7868|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Findings|7859,7868|false|false|false|C0001927|albuterol|albuterol
Event|Event|Findings|7859,7868|false|false|false|||albuterol
Drug|Organic Chemical|Findings|7859,7876|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Findings|7859,7876|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Findings|7869,7876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Findings|7869,7876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Findings|7869,7876|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Findings|7869,7876|false|false|false|||sulfate
Drug|Biomedical or Dental Material|Findings|7890,7898|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Drug|Substance|Findings|7890,7898|false|false|false|C0037633;C0525069;C1382100|Pharmaceutical Solutions;Solution Dosage Form;Solutions|Solution
Event|Event|Findings|7890,7898|false|false|false|||Solution
Finding|Conceptual Entity|Findings|7890,7898|false|false|false|C2699488|Resolution|Solution
Event|Event|Findings|7903,7915|false|false|false|||Nebulization
Procedure|Therapeutic or Preventive Procedure|Findings|7903,7915|false|false|false|C1659427|nebulization-mediated drug administration|Nebulization
Event|Event|Findings|7917,7920|false|false|false|||Sig
Event|Event|Findings|7930,7939|false|false|false|||treatment
Finding|Conceptual Entity|Findings|7930,7939|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Findings|7930,7939|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Findings|7930,7939|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Findings|7930,7939|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Event|Event|Findings|7940,7950|false|false|false|||Inhalation
Finding|Functional Concept|Findings|7940,7950|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Findings|7940,7950|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Event|Event|Findings|7970,7976|false|false|false|||needed
Event|Event|Findings|7982,7991|false|false|false|||shortness
Attribute|Clinical Attribute|Findings|7982,8001|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Findings|7982,8001|false|false|false|C0013404|Dyspnea|shortness of breath
Event|Event|Findings|7995,8001|false|false|false|||breath
Finding|Body Substance|Findings|7995,8001|false|false|false|C0225386|Breath|breath
Event|Event|Findings|8005,8013|false|false|false|||wheezing
Finding|Sign or Symptom|Findings|8005,8013|false|false|false|C0043144|Wheezing|wheezing
Finding|Idea or Concept|Findings|8046,8053|false|false|false|C0807726|refill|Refills
Event|Event|Findings|8061,8070|false|false|false|||Discharge
Finding|Body Substance|Findings|8061,8070|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Findings|8061,8070|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Findings|8061,8070|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Findings|8061,8070|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Findings|8061,8082|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Findings|8061,8082|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Findings|8071,8082|false|false|false|C2926604||Disposition
Event|Event|Findings|8071,8082|false|false|false|||Disposition
Procedure|Health Care Activity|Findings|8071,8082|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Findings|8084,8088|false|false|false|||Home
Finding|Idea or Concept|Findings|8084,8088|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Findings|8084,8088|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Findings|8084,8088|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Findings|8094,8101|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Findings|8094,8101|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Findings|8104,8112|false|false|false|||Facility
Finding|Intellectual Product|Findings|8104,8112|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Findings|8120,8129|false|false|false|||Discharge
Finding|Body Substance|Findings|8120,8129|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Findings|8120,8129|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Findings|8120,8129|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Findings|8120,8129|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Findings|8120,8139|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Findings|8130,8139|false|false|false|C0945731||Diagnosis
Event|Event|Findings|8130,8139|false|false|false|||Diagnosis
Finding|Classification|Findings|8130,8139|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Findings|8130,8139|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Findings|8130,8139|false|false|false|C0011900|Diagnosis|Diagnosis
Event|Event|Findings|8151,8166|false|false|false|||Tachyarrhythmia
Finding|Finding|Findings|8151,8166|false|false|false|C0080203|Tachyarrhythmia|Tachyarrhythmia
Disorder|Disease or Syndrome|Findings|8168,8182|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Findings|8168,8182|false|false|false|||Hyperlipidemia
Finding|Finding|Findings|8168,8182|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Disorder|Disease or Syndrome|Findings|8184,8190|false|false|false|C0004096|Asthma|Asthma
Event|Event|Findings|8184,8190|false|false|false|||Asthma
Disorder|Disease or Syndrome|Findings|8192,8196|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Findings|8192,8196|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Findings|8192,8196|false|false|false|||COPD
Finding|Gene or Genome|Findings|8192,8196|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Neoplastic Process|Findings|8198,8207|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|Findings|8198,8207|false|false|false|||Secondary
Finding|Functional Concept|Findings|8198,8207|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|Findings|8210,8222|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Findings|8210,8222|false|false|false|||Hypertension
Drug|Hazardous or Poisonous Substance|Findings|8225,8232|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Immunologic Factor|Findings|8225,8232|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Organic Chemical|Findings|8225,8232|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Drug|Pharmacologic Substance|Findings|8225,8232|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|Tobacco
Attribute|Clinical Attribute|Findings|8225,8236|false|false|false|C4522050||Tobacco Use
Finding|Finding|Findings|8225,8236|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco Use
Finding|Individual Behavior|Findings|8225,8236|false|false|false|C0040335;C0543414;C0841002;C3853727|Encounter due to tobacco use;History of tobacco use;Tobacco use;Tobacco user|Tobacco Use
Event|Event|Findings|8233,8236|false|false|false|||Use
Finding|Functional Concept|Findings|8233,8236|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Finding|Intellectual Product|Findings|8233,8236|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|Use
Finding|Mental Process|Discharge Condition|8263,8269|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|8263,8276|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|8263,8276|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|8270,8276|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|8270,8276|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8278,8283|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|8278,8283|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|8288,8296|false|false|false|||coherent
Finding|Finding|Discharge Condition|8288,8296|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|8298,8303|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|8298,8320|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|8298,8320|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|8307,8320|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|8307,8320|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|8307,8320|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|8322,8327|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|8322,8327|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|8322,8327|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|8322,8327|false|false|false|||Alert
Finding|Finding|Discharge Condition|8322,8327|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|8322,8327|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|8322,8327|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|8332,8343|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|8332,8343|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|8345,8353|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|8345,8353|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|8345,8353|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|8354,8360|false|false|false|C5889824||Status
Event|Event|Discharge Condition|8354,8360|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|8354,8360|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|8362,8372|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|8362,8372|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|8362,8372|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|8362,8372|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|8362,8372|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|8375,8386|false|false|false|||Independent
Finding|Finding|Discharge Condition|8375,8386|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|8375,8386|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|8435,8447|false|false|false|||hospitalized
Event|Event|Discharge Instructions|8469,8475|false|false|false|||nurses
Event|Event|Discharge Instructions|8481,8490|false|false|false|||concerned
Finding|Finding|Discharge Instructions|8501,8520|false|false|false|C4020868|Elevated heart rate|elevated heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8510,8515|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8510,8515|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8510,8515|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|8510,8520|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|8510,8520|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|8510,8520|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|8516,8520|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|8516,8520|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|8516,8520|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|Discharge Instructions|8533,8537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|8533,8537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|8533,8537|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|8542,8546|false|false|false|||came
Event|Event|Discharge Instructions|8555,8563|false|false|false|||hospital
Finding|Idea or Concept|Discharge Instructions|8555,8563|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|Discharge Instructions|8570,8589|false|false|false|C4020868|Elevated heart rate|elevated heart rate
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8579,8584|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8579,8584|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8579,8584|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|Discharge Instructions|8579,8589|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|Discharge Instructions|8579,8589|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|Discharge Instructions|8579,8589|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|Discharge Instructions|8585,8589|false|false|false|C0871208|Rating (action)|rate
Event|Event|Discharge Instructions|8585,8589|false|false|false|||rate
Finding|Idea or Concept|Discharge Instructions|8585,8589|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|Discharge Instructions|8594,8602|false|false|false|||resolved
Event|Event|Discharge Instructions|8629,8637|false|false|false|||admitted
Event|Event|Discharge Instructions|8641,8647|false|false|false|||ensure
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8658,8663|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|8658,8663|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|8658,8663|false|false|false|C0795691|HEART PROBLEM|heart
Event|Event|Discharge Instructions|8671,8679|false|false|false|||suffered
Disorder|Injury or Poisoning|Discharge Instructions|8685,8691|false|false|false|C0010957|Tissue damage|damage
Event|Event|Discharge Instructions|8685,8691|false|false|false|||damage
Finding|Functional Concept|Discharge Instructions|8685,8691|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Finding|Gene or Genome|Discharge Instructions|8685,8691|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Event|Event|Discharge Instructions|8700,8703|false|false|false|||see
Event|Event|Discharge Instructions|8708,8717|false|false|false|||inpatient
Finding|Idea or Concept|Discharge Instructions|8708,8717|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Discharge Instructions|8708,8717|false|false|false|C1555324|inpatient encounter|inpatient
Lab|Laboratory or Test Result|Discharge Instructions|8738,8742|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|Discharge Instructions|8749,8761|false|false|false|||unremarkable
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8769,8776|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Discharge Instructions|8769,8776|false|false|false|C1314974|Cardiac attachment|cardiac
Event|Event|Discharge Instructions|8797,8800|false|false|false|||saw
Event|Event|Discharge Instructions|8824,8833|false|false|false|||recommend
Event|Event|Discharge Instructions|8837,8849|false|false|false|||intervention
Procedure|Health Care Activity|Discharge Instructions|8837,8849|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|8837,8849|true|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Finding|Discharge Instructions|8858,8862|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|8858,8862|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|8858,8862|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|8878,8884|false|false|false|||follow
Finding|Classification|Discharge Instructions|8918,8928|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|8918,8928|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Attribute|Clinical Attribute|Discharge Instructions|8939,8948|false|false|false|C5885990||breathing
Finding|Finding|Discharge Instructions|8939,8948|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|8939,8948|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|8939,8948|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|8939,8948|false|false|false|C1160636|respiratory system process|breathing
Event|Event|Discharge Instructions|8949,8955|false|false|false|||issues
Disorder|Disease or Syndrome|Discharge Instructions|8962,8966|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|8962,8966|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|8962,8966|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Anatomy|Body Location or Region|Discharge Instructions|8993,8997|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|8993,8997|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|8993,8997|false|false|false|C0024115|Lung diseases|lung
Event|Event|Discharge Instructions|8993,8997|false|false|false|||lung
Finding|Finding|Discharge Instructions|8993,8997|false|false|false|C0740941|Lung Problem|lung
Event|Event|Discharge Instructions|8999,9005|false|false|false|||health
Finding|Idea or Concept|Discharge Instructions|8999,9005|false|false|false|C0018684|Health|health
Event|Event|Discharge Instructions|9012,9016|false|false|false|||quit
Event|Event|Discharge Instructions|9017,9024|false|false|false|||smoking
Event|Event|Discharge Instructions|9033,9042|false|false|false|||encourage
Event|Event|Discharge Instructions|9072,9079|false|false|false|||changes
Finding|Functional Concept|Discharge Instructions|9072,9079|false|false|false|C0392747|Changing|changes
Event|Event|Discharge Instructions|9085,9089|false|false|false|||made
Attribute|Clinical Attribute|Discharge Instructions|9098,9109|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|9098,9109|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|9098,9109|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|9098,9109|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|9112,9120|false|false|false|||INCREASE
Finding|Functional Concept|Discharge Instructions|9112,9120|false|false|false|C0442805|Increase|INCREASE
Drug|Organic Chemical|Discharge Instructions|9126,9137|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Discharge Instructions|9126,9137|false|false|false|C0074554|simvastatin|simvastatin
Event|Event|Discharge Instructions|9126,9137|false|false|false|||simvastatin
Event|Activity|Discharge Instructions|9155,9160|false|false|false|C1705178|Order (action)|order
Finding|Classification|Discharge Instructions|9155,9160|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Idea or Concept|Discharge Instructions|9155,9160|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Intellectual Product|Discharge Instructions|9155,9160|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|9155,9160|false|false|false|C1373200|Order [PK]|order
Drug|Biologically Active Substance|Discharge Instructions|9176,9187|false|false|false|C0008377|cholesterol|cholesterol
Drug|Organic Chemical|Discharge Instructions|9176,9187|false|false|false|C0008377|cholesterol|cholesterol
Event|Event|Discharge Instructions|9176,9187|false|false|false|||cholesterol
Procedure|Laboratory Procedure|Discharge Instructions|9176,9187|false|false|false|C0201950|Cholesterol measurement|cholesterol
Event|Event|Discharge Instructions|9191,9195|false|false|false|||goal
Finding|Idea or Concept|Discharge Instructions|9191,9195|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Discharge Instructions|9191,9195|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|Discharge Instructions|9200,9211|false|false|false|||recommended
Drug|Organic Chemical|Discharge Instructions|9242,9254|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Discharge Instructions|9242,9254|false|false|false|C0039771|theophylline|theophylline
Event|Event|Discharge Instructions|9242,9254|false|false|false|||theophylline
Procedure|Laboratory Procedure|Discharge Instructions|9242,9254|false|false|false|C0039773|Assay of theophylline|theophylline
Disorder|Disease or Syndrome|Discharge Instructions|9267,9272|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Discharge Instructions|9275,9278|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|9275,9278|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|9296,9302|false|false|false|||giving
Attribute|Clinical Attribute|Discharge Instructions|9309,9321|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Discharge Instructions|9309,9321|false|false|false|||prescription
Finding|Intellectual Product|Discharge Instructions|9309,9321|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Discharge Instructions|9309,9321|false|false|false|C0033080|Prescription (procedure)|prescription
Drug|Organic Chemical|Discharge Instructions|9326,9335|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Discharge Instructions|9326,9335|false|false|false|C0001927|albuterol|albuterol
Event|Event|Discharge Instructions|9326,9335|false|false|false|||albuterol
Drug|Pharmacologic Substance|Discharge Instructions|9337,9347|false|false|false|C2064916|nebulizers (medication)|nebulizers
Event|Event|Discharge Instructions|9337,9347|false|false|false|||nebulizers
Event|Event|Discharge Instructions|9351,9354|false|false|false|||use
Event|Event|Discharge Instructions|9371,9378|false|false|false|||inhaler
Finding|Functional Concept|Discharge Instructions|9371,9378|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Event|Event|Discharge Instructions|9385,9391|false|false|false|||needed
Event|Event|Discharge Instructions|9399,9406|false|false|false|||refills
Attribute|Clinical Attribute|Discharge Instructions|9444,9453|false|false|false|C0804815||physician
Event|Event|Discharge Instructions|9477,9484|false|false|false|||discuss
Drug|Organic Chemical|Discharge Instructions|9490,9502|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Discharge Instructions|9490,9502|false|false|false|C0039771|theophylline|theophylline
Event|Event|Discharge Instructions|9490,9502|false|false|false|||theophylline
Procedure|Laboratory Procedure|Discharge Instructions|9490,9502|false|false|false|C0039773|Assay of theophylline|theophylline
Attribute|Clinical Attribute|Discharge Instructions|9490,9507|false|false|true|C0366665||theophylline dose
Event|Event|Discharge Instructions|9503,9507|false|false|false|||dose
Attribute|Clinical Attribute|Discharge Instructions|9512,9521|false|false|true|C5885990||breathing
Event|Event|Discharge Instructions|9512,9521|false|false|false|||breathing
Finding|Finding|Discharge Instructions|9512,9521|false|false|true|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|9512,9521|false|false|true|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|9512,9521|false|false|true|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|9512,9521|false|false|true|C1160636|respiratory system process|breathing
Attribute|Clinical Attribute|Discharge Instructions|9522,9528|false|false|false|C5889824||status
Event|Event|Discharge Instructions|9522,9528|false|false|false|||status
Finding|Idea or Concept|Discharge Instructions|9522,9528|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Discharge Instructions|9548,9556|false|false|false|||provider
Finding|Functional Concept|Discharge Instructions|9548,9556|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|Discharge Instructions|9548,9556|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Procedure|Health Care Activity|Discharge Instructions|9604,9612|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9613,9625|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|9613,9625|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|9613,9625|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

