 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|164,173|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|164,173|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|185,194|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|SIMPLE_SEGMENT|222,231|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|240,255|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|246,255|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|246,255|false|false|false|C5441521|Complaint (finding)|Complaint
Finding|Sign or Symptom|SIMPLE_SEGMENT|257,264|false|false|false|C0039070|Syncope|Syncope
Finding|Classification|SIMPLE_SEGMENT|267,272|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|273,281|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|273,281|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|285,303|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|294,303|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|294,303|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|294,303|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|294,303|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|312,319|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|312,322|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|312,338|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|312,338|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|323,330|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|323,330|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|323,338|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|331,338|false|false|false|C0221423|Illness (finding)|Illness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|369,383|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|395,398|false|false|false|C0020538|Hypertensive disease|HTN
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|401,404|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Finding|Functional Concept|SIMPLE_SEGMENT|423,431|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|423,431|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|423,431|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Intellectual Product|SIMPLE_SEGMENT|545,554|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|545,554|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Intellectual Product|SIMPLE_SEGMENT|550,554|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|550,554|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|SIMPLE_SEGMENT|556,567|false|false|false|C0220870|Lightheadedness|lightheaded
Finding|Sign or Symptom|SIMPLE_SEGMENT|573,581|false|false|false|C0027497|Nausea|nauseous
Finding|Sign or Symptom|SIMPLE_SEGMENT|602,619|false|false|false|C0751534|Syncopal Episode|syncopal episodes
Finding|Intellectual Product|SIMPLE_SEGMENT|644,651|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|644,651|false|false|false|C0700287|Reporting|reports
Finding|Idea or Concept|SIMPLE_SEGMENT|679,685|false|false|false|C0018684|Health|health
Finding|Idea or Concept|SIMPLE_SEGMENT|686,694|false|false|false|C1546466|Problems - What subject filter|problems
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|713,716|false|false|false|C0600500|Peptide Nucleic Acids|PNA
Finding|Sign or Symptom|SIMPLE_SEGMENT|729,739|false|false|false|C0019079|Hemoptysis|hemoptysis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|756,763|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|759,763|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|772,775|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|799,812|false|true|false|C0521530|Lung consolidation|consolidation
Finding|Finding|SIMPLE_SEGMENT|829,836|false|false|false|C3845930|Copious|copious
Finding|Body Substance|SIMPLE_SEGMENT|844,854|false|false|false|C0036537|Bodily secretions|secretions
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|855,858|false|false|false|C4281590|Structure of middle lobe of right lung|RML
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|859,866|false|false|false|C0225740;C0228475;C1561517|Lingula;Lingula of cerebellum;Lingula of left lung|lingula
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|867,870|false|false|false|C1261074|Structure of right upper lobe of lung|RUL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|881,886|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|881,886|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|914,921|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|917,921|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Intellectual Product|SIMPLE_SEGMENT|970,974|false|false|false|C1720594|Then - dosing instruction fragment|then
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|996,1008|false|false|false|C0752295|Confusional Arousals|unresponsive
Finding|Finding|SIMPLE_SEGMENT|996,1008|false|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Finding|Functional Concept|SIMPLE_SEGMENT|996,1008|false|false|false|C0205269;C0237284|Unresponsive to Treatment;unresponsive behavior|unresponsive
Finding|Sign or Symptom|SIMPLE_SEGMENT|1042,1050|true|false|false|C0240805|Prodrome|prodrome
Finding|Finding|SIMPLE_SEGMENT|1055,1067|false|false|false|C0030252|Palpitations|palpitations
Finding|Finding|SIMPLE_SEGMENT|1082,1095|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|SIMPLE_SEGMENT|1082,1095|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1113,1122|false|false|false|C0009676|Confusion|confusion
Finding|Finding|SIMPLE_SEGMENT|1113,1122|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Sign or Symptom|SIMPLE_SEGMENT|1138,1145|true|false|false|C0036572|Seizures|seizure
Event|Activity|SIMPLE_SEGMENT|1151,1159|false|false|false|C0441655|Activities|activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|1151,1159|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|SIMPLE_SEGMENT|1151,1159|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1183,1188|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1192,1199|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1192,1199|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1192,1199|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Organism Function|SIMPLE_SEGMENT|1219,1227|true|false|false|C0015264|Exertion|exertion
Finding|Finding|SIMPLE_SEGMENT|1272,1284|true|false|false|C0030252|Palpitations|palpitations
Finding|Sign or Symptom|SIMPLE_SEGMENT|1286,1289|true|false|false|C0013404|Dyspnea|SOB
Finding|Body Substance|SIMPLE_SEGMENT|1433,1439|false|false|false|C0225378|Upper respiratory tract mucus|phlegm
Finding|Finding|SIMPLE_SEGMENT|1475,1479|false|false|false|C5575035|Well (answer to question)|well
Finding|Sign or Symptom|SIMPLE_SEGMENT|1490,1496|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1497,1503|false|false|false|C0085593|Chills|chills
Procedure|Health Care Activity|SIMPLE_SEGMENT|1514,1518|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1514,1518|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Gene or Genome|SIMPLE_SEGMENT|1536,1539|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Idea or Concept|SIMPLE_SEGMENT|1554,1561|false|false|false|C1555582|Initial (abbreviation)|initial
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|1597,1601|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|SIMPLE_SEGMENT|1620,1623|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1654,1657|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1654,1657|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Anatomy|Cell|SIMPLE_SEGMENT|1691,1694|false|false|false|C0023516|Leukocytes|WBC
Finding|Functional Concept|SIMPLE_SEGMENT|1712,1720|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1712,1720|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1712,1720|false|false|false|C4706767|Transfer (immobility management)|transfer
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1766,1774|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1775,1780|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Sign or Symptom|SIMPLE_SEGMENT|1818,1823|false|false|false|C0012833|Dizziness|dizzy
Finding|Sign or Symptom|SIMPLE_SEGMENT|1827,1838|false|false|false|C0220870|Lightheadedness|lightheaded
Finding|Finding|SIMPLE_SEGMENT|1851,1856|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1851,1856|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1858,1864|false|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1866,1872|true|false|false|C2707266||vision
Finding|Organism Function|SIMPLE_SEGMENT|1866,1872|true|false|false|C0042789|Vision|vision
Finding|Functional Concept|SIMPLE_SEGMENT|1874,1881|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1883,1902|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|1883,1902|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|1896,1902|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1904,1909|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1904,1909|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1904,1914|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1904,1914|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1910,1914|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1910,1914|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1910,1914|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1910,1925|false|false|false|C0000737|Abdominal Pain|pain, abdominal
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1916,1925|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1916,1930|false|true|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1926,1930|false|true|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1926,1930|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1926,1930|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1933,1939|false|false|false|C4255480||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1933,1939|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1941,1949|false|false|false|C0042963|Vomiting|vomiting
Finding|Finding|SIMPLE_SEGMENT|1951,1959|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1951,1959|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1961,1973|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1975,1980|false|false|false|C0018932|Hematochezia|BRBPR
Finding|Pathologic Function|SIMPLE_SEGMENT|1982,1988|false|false|false|C0025222|Melena|melena
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1991,2003|false|false|false|C0018932|Hematochezia|hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|1991,2003|false|false|false|C1321898|Blood in stool|hematochezia
Finding|Sign or Symptom|SIMPLE_SEGMENT|2005,2012|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2014,2023|false|false|false|C0018965|Hematuria|hematuria
Finding|Functional Concept|SIMPLE_SEGMENT|2042,2046|false|false|false|C0745777|Lost|lost
Finding|Gene or Genome|SIMPLE_SEGMENT|2101,2106|true|false|false|C1424898|RXFP2 gene|great
Finding|Organism Function|SIMPLE_SEGMENT|2107,2115|false|false|false|C0003618|Desire for food|appetite
Finding|Idea or Concept|SIMPLE_SEGMENT|2129,2134|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|2129,2134|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Finding|SIMPLE_SEGMENT|2138,2158|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|2143,2150|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2143,2150|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2143,2150|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2143,2150|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2143,2158|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2151,2158|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2151,2158|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2151,2158|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2160,2163|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2164,2178|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Finding|Gene or Genome|SIMPLE_SEGMENT|2188,2191|false|false|false|C1417026|MAPK8IP3 gene|Syd
Finding|Functional Concept|SIMPLE_SEGMENT|2195,2201|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2195,2209|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2202,2209|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2202,2209|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2202,2209|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2215,2221|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2215,2221|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2215,2221|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2215,2221|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2215,2229|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2222,2229|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2222,2229|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2222,2229|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2236,2243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2236,2243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2236,2243|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2236,2246|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|2236,2259|false|false|false|C0455527||history of hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2247,2259|false|false|false|C0020538|Hypertensive disease|hypertension
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2263,2273|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|SIMPLE_SEGMENT|2263,2273|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|SIMPLE_SEGMENT|2263,2273|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|SIMPLE_SEGMENT|2267,2273|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2267,2273|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2267,2273|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2267,2273|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2285,2291|false|false|false|C4255046||report
Finding|Intellectual Product|SIMPLE_SEGMENT|2285,2291|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|SIMPLE_SEGMENT|2285,2291|false|false|false|C0700287|Reporting|report
Finding|Conceptual Entity|SIMPLE_SEGMENT|2302,2308|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Idea or Concept|SIMPLE_SEGMENT|2302,2308|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|father
Finding|Classification|SIMPLE_SEGMENT|2311,2317|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2311,2317|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2311,2317|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2311,2317|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2324,2331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2324,2331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2324,2331|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2324,2334|false|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2344,2351|false|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|SIMPLE_SEGMENT|2384,2391|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2384,2391|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2384,2391|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2384,2394|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2395,2402|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2395,2402|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2395,2402|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|SIMPLE_SEGMENT|2395,2402|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2395,2402|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2395,2409|false|false|false|C0024623;C0699791|Malignant neoplasm of stomach;Stomach Carcinoma|stomach cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2403,2409|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|2431,2438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2431,2438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2431,2438|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2431,2441|false|false|false|C0262926|Medical History|history of
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2442,2448|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2442,2448|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2442,2448|false|false|false|C1950455|Throat Homeopathic Medication|throat
Finding|Body Substance|SIMPLE_SEGMENT|2442,2448|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|SIMPLE_SEGMENT|2442,2448|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2442,2455|false|false|false|C0740339|Throat cancer|throat cancer
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2449,2455|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|2473,2480|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2473,2480|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2473,2480|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2473,2483|true|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2485,2490|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2485,2490|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2485,2490|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|SIMPLE_SEGMENT|2485,2490|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2485,2498|false|false|false|C0007102|Malignant tumor of colon|colon cancers
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2491,2498|false|false|false|C0006826|Malignant Neoplasms|cancers
Finding|Conceptual Entity|SIMPLE_SEGMENT|2500,2506|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|2500,2506|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2511,2517|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|SIMPLE_SEGMENT|2511,2517|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Classification|SIMPLE_SEGMENT|2522,2528|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2522,2528|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2522,2528|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2522,2528|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2537,2543|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2551,2556|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2551,2556|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|2551,2556|false|false|false|C0795691|HEART PROBLEM|heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2551,2562|false|false|false|C0018826;C1305961|Heart Valves|heart valve
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2557,2562|false|false|false|C1186983|Anatomical valve|valve
Finding|Intellectual Product|SIMPLE_SEGMENT|2580,2584|true|false|false|C4724437|SURE Test|sure
Finding|Finding|SIMPLE_SEGMENT|2600,2608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2600,2608|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2600,2608|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2600,2613|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2600,2613|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2609,2613|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2609,2613|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2615,2624|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|SIMPLE_SEGMENT|2625,2629|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2625,2629|false|false|false|C0582103|Medical Examination|EXAM
Finding|Gene or Genome|SIMPLE_SEGMENT|2637,2641|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2637,2641|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Classification|SIMPLE_SEGMENT|2687,2694|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2687,2694|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2721,2724|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2721,2724|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2721,2724|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2721,2724|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2721,2724|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|2721,2724|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Finding|Finding|SIMPLE_SEGMENT|2726,2737|false|false|false|C5546696|Feeling comfortable|comfortable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2751,2756|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|2766,2771|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|SIMPLE_SEGMENT|2787,2796|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2798,2801|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2798,2801|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Idea or Concept|SIMPLE_SEGMENT|2806,2811|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2812,2816|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2812,2816|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2812,2816|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|SIMPLE_SEGMENT|2819,2825|false|false|false|C0332254|Supple|supple
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2830,2841|true|false|false|C0018021|Goiter|thyromegaly
Finding|Finding|SIMPLE_SEGMENT|2846,2849|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2851,2858|false|false|false|C0007272|Carotid Arteries|carotid
Finding|Finding|SIMPLE_SEGMENT|2851,2865|false|false|false|C0007280|Carotid bruit|carotid bruits
Finding|Finding|SIMPLE_SEGMENT|2859,2865|false|false|false|C0006318|Bruit|bruits
Finding|Finding|SIMPLE_SEGMENT|2867,2873|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|2867,2873|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2885,2891|false|false|false|C0037709||sounds
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2897,2903|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2897,2917|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|SIMPLE_SEGMENT|2904,2917|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|2904,2917|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|2904,2917|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2919,2924|false|false|false|C0024109|Lung|LUNGS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2927,2930|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|2927,2930|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2927,2930|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Idea or Concept|SIMPLE_SEGMENT|2950,2954|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|2955,2958|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2955,2958|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|2955,2958|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|2955,2958|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|2955,2958|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|2955,2958|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2955,2967|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|2959,2967|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2969,2973|false|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2969,2973|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Finding|Functional Concept|SIMPLE_SEGMENT|2975,2984|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2989,3005|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|2989,3009|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2999,3005|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|2999,3005|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|SIMPLE_SEGMENT|3006,3009|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3006,3009|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3010,3015|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3010,3015|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|3010,3015|false|false|false|C0795691|HEART PROBLEM|HEART
Finding|Finding|SIMPLE_SEGMENT|3026,3045|false|false|false|C0232259|Mid-systolic murmur|mid-systolic murmur
Finding|Finding|SIMPLE_SEGMENT|3039,3045|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3057,3060|false|false|false|C0175200|lateral longitudinal stria|LLS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3057,3060|false|false|false|C4085873|LUSCAN-LUMISH SYNDROME|LLS
Finding|Gene or Genome|SIMPLE_SEGMENT|3057,3060|false|false|false|C2348110|SETD2 wt Allele|LLS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3061,3067|false|false|false|C1522411|Anatomic Border|border
Finding|Idea or Concept|SIMPLE_SEGMENT|3061,3067|false|false|false|C1552830|Table Frame - border|border
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3082,3088|false|false|false|C0004454|Axilla|axilla
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3099,3106|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3099,3106|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3099,3106|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3115,3119|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Gene or Genome|SIMPLE_SEGMENT|3140,3143|true|false|false|C1537594|LRRC4B gene|HSM
Finding|Finding|SIMPLE_SEGMENT|3157,3165|false|false|false|C0427198|Protective muscle spasm|guarding
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3166,3177|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3198,3215|false|false|false|C0232139|Peripheral pulse|peripheral pulses
Drug|Food|SIMPLE_SEGMENT|3209,3215|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3209,3215|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3209,3215|false|false|false|C0034107|Pulse taking|pulses
Finding|Gene or Genome|SIMPLE_SEGMENT|3226,3229|false|false|false|C1843919|PDSS1 gene|DPs
Finding|Finding|SIMPLE_SEGMENT|3239,3244|false|false|false|C0234422|Awake (finding)|awake
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3253,3259|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|3253,3259|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3253,3268|false|false|false|C4050373||muscle strength
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3253,3268|false|false|false|C0517349|Muscle Strength|muscle strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3260,3268|false|false|false|C0808080|Strength (attribute)|strength
Finding|Body Substance|SIMPLE_SEGMENT|3280,3289|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3280,3289|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3280,3289|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3280,3289|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|SIMPLE_SEGMENT|3290,3294|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|3290,3294|false|false|false|C0582103|Medical Examination|EXAM
Finding|Finding|SIMPLE_SEGMENT|3296,3305|false|false|false|C0442739||Unchanged
Finding|Gene or Genome|SIMPLE_SEGMENT|3353,3357|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3353,3357|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3403,3408|false|false|false|C0024109|Lung|LUNGS
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3411,3414|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|SIMPLE_SEGMENT|3411,3414|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3411,3414|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Finding|Idea or Concept|SIMPLE_SEGMENT|3434,3438|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3439,3442|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3439,3442|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|SIMPLE_SEGMENT|3439,3442|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|SIMPLE_SEGMENT|3439,3442|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|SIMPLE_SEGMENT|3439,3442|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|SIMPLE_SEGMENT|3439,3442|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3439,3451|false|false|false|C0001868|Air Movements|air movement
Finding|Organism Function|SIMPLE_SEGMENT|3443,3451|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3453,3457|false|false|false|C0231832|Respiratory rate|resp
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3453,3457|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|resp
Finding|Functional Concept|SIMPLE_SEGMENT|3459,3468|false|false|false|C2983702|Unlabored|unlabored
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3473,3489|true|false|false|C0158784|Accessory skeletal muscle|accessory muscle
Finding|Finding|SIMPLE_SEGMENT|3473,3493|true|false|false|C1821466|Use of accessory muscles|accessory muscle use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3483,3489|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Anatomy|Tissue|SIMPLE_SEGMENT|3483,3489|false|false|false|C0026845;C4083049|Muscle (organ);Muscle Tissue|muscle
Finding|Functional Concept|SIMPLE_SEGMENT|3490,3493|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3490,3493|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3494,3499|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3494,3499|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|SIMPLE_SEGMENT|3494,3499|false|false|false|C0795691|HEART PROBLEM|HEART
Finding|Finding|SIMPLE_SEGMENT|3510,3529|false|false|false|C0232259|Mid-systolic murmur|mid-systolic murmur
Finding|Finding|SIMPLE_SEGMENT|3523,3529|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3545,3551|false|false|false|C1522411|Anatomic Border|border
Finding|Idea or Concept|SIMPLE_SEGMENT|3545,3551|false|false|false|C1552830|Table Frame - border|border
Procedure|Health Care Activity|SIMPLE_SEGMENT|3603,3612|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3613,3617|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3631,3636|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3631,3636|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3637,3640|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3648,3651|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3648,3651|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3648,3651|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3658,3661|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3658,3661|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3658,3661|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3658,3661|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3668,3671|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3668,3671|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3679,3682|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3679,3682|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3679,3682|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3679,3682|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3686,3689|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3686,3689|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3686,3689|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3686,3689|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3686,3689|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3696,3700|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3715,3718|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3735,3740|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3735,3740|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3753,3759|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|3766,3771|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3766,3771|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3766,3771|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3777,3780|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3777,3780|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3806,3811|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3806,3811|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3812,3815|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3832,3837|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3832,3837|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|3832,3845|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3832,3845|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3832,3845|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3838,3845|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|3838,3845|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3838,3845|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3838,3845|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3838,3845|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|3891,3895|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3891,3895|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3891,3895|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3920,3925|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3920,3925|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3952,3957|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3952,3957|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3974,3983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3974,3983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3974,3983|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3974,3983|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3984,3988|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4002,4007|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4002,4007|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4008,4011|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4016,4019|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4016,4019|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4016,4019|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4026,4029|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4026,4029|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4026,4029|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4026,4029|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4036,4039|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4036,4039|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4047,4050|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4047,4050|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4047,4050|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4047,4050|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4054,4057|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4054,4057|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4054,4057|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4054,4057|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4054,4057|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4064,4068|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4083,4086|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4103,4108|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4103,4108|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4109,4112|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4129,4134|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4129,4134|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4129,4142|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4129,4142|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4129,4142|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4135,4142|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4135,4142|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4135,4142|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4135,4142|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4135,4142|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4187,4191|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4187,4191|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4187,4191|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4216,4221|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4216,4221|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4216,4229|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4222,4229|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4222,4229|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4222,4229|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4222,4229|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|4222,4229|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|4222,4229|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4222,4229|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4262,4267|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4262,4267|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4262,4272|false|false|false|C0853169|Blood iron measurement|BLOOD Iron
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4268,4272|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4268,4272|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4268,4272|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4268,4272|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4288,4293|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4288,4293|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4349,4352|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4349,4352|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|4349,4352|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4349,4352|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|4349,4352|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Finding|Functional Concept|SIMPLE_SEGMENT|4359,4371|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|4359,4371|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4359,4371|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4377,4382|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|SIMPLE_SEGMENT|4377,4382|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Finding|Idea or Concept|SIMPLE_SEGMENT|4387,4394|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|Pending
Finding|Body Substance|SIMPLE_SEGMENT|4399,4404|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|4399,4404|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|4399,4404|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Idea or Concept|SIMPLE_SEGMENT|4409,4416|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Finding|SIMPLE_SEGMENT|4419,4426|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4419,4426|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Finding|Intellectual Product|SIMPLE_SEGMENT|4432,4437|false|false|false|C3463807|Video Media|Video
Finding|Functional Concept|SIMPLE_SEGMENT|4438,4445|false|false|false|C1706486;C4521686|Swallow (administration method);Swallow - dosing instruction imperative|swallow
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4438,4451|false|false|false|C3888792|Swallow study|swallow study
Finding|Intellectual Product|SIMPLE_SEGMENT|4446,4451|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|4446,4451|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Finding|SIMPLE_SEGMENT|4457,4463|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|4457,4463|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4464,4474|false|true|false|C1720922|Respiratory Aspiration|aspiration
Finding|Finding|SIMPLE_SEGMENT|4464,4474|false|true|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4464,4474|false|true|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|4464,4474|false|true|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4464,4474|false|true|false|C0349707||aspiration
Finding|Idea or Concept|SIMPLE_SEGMENT|4477,4492|false|false|false|C0034866|Recommendation|RECOMMENDATIONS
Drug|Food|SIMPLE_SEGMENT|4500,4504|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|4500,4504|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|4500,4504|false|false|false|C0012159|Diet therapy|diet
Drug|Substance|SIMPLE_SEGMENT|4513,4520|false|false|false|C0302908|Liquid substance|liquids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4525,4529|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4530,4536|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Drug|Substance|SIMPLE_SEGMENT|4530,4536|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4541,4551|false|false|false|C1720922|Respiratory Aspiration|Aspiration
Finding|Finding|SIMPLE_SEGMENT|4541,4551|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|Aspiration
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|4541,4551|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|Aspiration
Finding|Pathologic Function|SIMPLE_SEGMENT|4541,4551|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|Aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4541,4551|false|false|false|C0349707||Aspiration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4541,4563|false|false|false|C0150138|Aspiration precautions|Aspiration precautions
Finding|Conceptual Entity|SIMPLE_SEGMENT|4552,4563|false|false|false|C1882442|Precaution|precautions
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4584,4590|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Drug|Substance|SIMPLE_SEGMENT|4584,4590|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4591,4595|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Functional Concept|SIMPLE_SEGMENT|4610,4613|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|4610,4613|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4614,4620|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Drug|Substance|SIMPLE_SEGMENT|4614,4620|false|false|false|C0302908;C1697794|Liquid Dosage Form;Liquid substance|liquid
Finding|Finding|SIMPLE_SEGMENT|4614,4620|false|false|false|C1304698|Liquid (finding)|liquid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4614,4620|false|false|false|C0301571|Liquid diet|liquid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4621,4625|false|false|false|C1883550|Wash Dosage Form|wash
Event|Activity|SIMPLE_SEGMENT|4621,4625|false|false|false|C0441648|Wash (cleansing action)|wash
Finding|Functional Concept|SIMPLE_SEGMENT|4621,4625|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Finding|Gene or Genome|SIMPLE_SEGMENT|4621,4625|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Finding|Intellectual Product|SIMPLE_SEGMENT|4621,4625|false|false|false|C1547959;C1549545;C2240171;C5779845|WASHC1 gene;Wash - Administration Method;Wash - Specimen Source Codes;Wash - dosing instruction imperative|wash
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4621,4625|false|false|false|C2699154|Cell Wash|wash
Finding|Idea or Concept|SIMPLE_SEGMENT|4629,4634|false|false|false|C1550016|Remote control command - Clear|clear
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4636,4642|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Drug|Substance|SIMPLE_SEGMENT|4636,4642|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|solids
Finding|Functional Concept|SIMPLE_SEGMENT|4657,4666|false|false|false|C0332270;C1552848|Alternating;alternate - HtmlLinkType|alternate
Finding|Idea or Concept|SIMPLE_SEGMENT|4657,4666|false|false|false|C0332270;C1552848|Alternating;alternate - HtmlLinkType|alternate
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|4667,4672|false|false|false|C0005658|bite injury|bites
Finding|Cell Function|SIMPLE_SEGMENT|4677,4681|false|false|false|C3157027;C4255036|Sips;stress-induced premature senescence|sips
Finding|Finding|SIMPLE_SEGMENT|4677,4681|false|false|false|C3157027;C4255036|Sips;stress-induced premature senescence|sips
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4685,4689|false|false|false|C3280240|MICROCEPHALY, EPILEPSY, AND DIABETES SYNDROME 1|Meds
Finding|Intellectual Product|SIMPLE_SEGMENT|4685,4689|false|false|false|C4284232|Medications|Meds
Finding|Functional Concept|SIMPLE_SEGMENT|4696,4706|false|false|false|C1883711|With Water|with water
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4701,4706|false|false|false|C0043047;C1550678|Water Specimen;water|water
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4701,4706|false|false|false|C0043047;C1550678|Water Specimen;water|water
Finding|Intellectual Product|SIMPLE_SEGMENT|4701,4706|false|false|false|C1547961|Water - Specimen Source Codes|water
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4701,4706|false|false|false|C0020311|Hydrotherapy|water
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|4719,4723|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4719,4723|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|4719,4723|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|4719,4723|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Procedure|Health Care Activity|SIMPLE_SEGMENT|4719,4728|false|false|false|C1272386;C2599893|Mouth care management;Oral care|oral care
Event|Activity|SIMPLE_SEGMENT|4724,4728|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|4724,4728|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|4724,4728|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4740,4751|false|false|false|C2707262||nutritional
Drug|Food|SIMPLE_SEGMENT|4740,4763|false|true|false|C0242295|Dietary Supplements|nutritional supplements
Finding|Finding|SIMPLE_SEGMENT|4764,4771|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|4767,4771|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4767,4771|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4767,4771|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4778,4785|false|false|false|C0684224|Report (document)|reports
Procedure|Health Care Activity|SIMPLE_SEGMENT|4778,4785|false|false|false|C0700287|Reporting|reports
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4797,4803|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|4797,4803|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|4797,4803|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|4797,4803|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|4797,4808|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|4797,4808|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|SIMPLE_SEGMENT|4804,4808|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Intellectual Product|SIMPLE_SEGMENT|4812,4817|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|4818,4826|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4818,4833|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|4818,4833|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Mental Process|SIMPLE_SEGMENT|4848,4856|false|false|false|C2987187|Pleasant|pleasant
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4870,4876|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4870,4890|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|SIMPLE_SEGMENT|4877,4890|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|4877,4890|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|4877,4890|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4893,4907|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4923,4926|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Functional Concept|SIMPLE_SEGMENT|4945,4953|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|4945,4953|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|4945,4953|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Sign or Symptom|SIMPLE_SEGMENT|4972,4988|false|false|false|C0751534|Syncopal Episode|syncopal episode
Procedure|Health Care Activity|SIMPLE_SEGMENT|5005,5014|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|SIMPLE_SEGMENT|5025,5047|false|false|false|C0578150|Hemodynamically stable|hemodynamically stable
Finding|Intellectual Product|SIMPLE_SEGMENT|5041,5047|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|SIMPLE_SEGMENT|5072,5084|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Finding|SIMPLE_SEGMENT|5085,5091|false|false|false|C0034359|Pyuria|pyuria
Drug|Organic Chemical|SIMPLE_SEGMENT|5093,5098|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5093,5098|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|5093,5098|false|false|false|C0010200|Coughing|cough
Anatomy|Cell|SIMPLE_SEGMENT|5106,5109|false|false|false|C0023516|Leukocytes|WBC
Finding|Sign or Symptom|SIMPLE_SEGMENT|5139,5146|false|false|false|C0039070|Syncope|Syncope
Finding|Sign or Symptom|SIMPLE_SEGMENT|5153,5169|false|false|false|C0751534|Syncopal Episode|syncopal episode
Finding|Functional Concept|SIMPLE_SEGMENT|5188,5197|false|false|false|C1519959|Vasovagal|vasovagal
Finding|Sign or Symptom|SIMPLE_SEGMENT|5199,5206|false|false|false|C0039070|Syncope|syncope
Finding|Finding|SIMPLE_SEGMENT|5208,5214|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5208,5214|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Mental Process|SIMPLE_SEGMENT|5222,5229|false|false|false|C0542559|contextual factors|setting
Finding|Finding|SIMPLE_SEGMENT|5237,5249|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Finding|Finding|SIMPLE_SEGMENT|5250,5256|false|false|false|C0034359|Pyuria|pyuria
Finding|Classification|SIMPLE_SEGMENT|5301,5309|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|5301,5309|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5301,5309|false|false|false|C5237010|Expression Negative|negative
Finding|Intellectual Product|SIMPLE_SEGMENT|5317,5320|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5317,5320|false|false|false|C1623258|Electrocardiography|EKG
Finding|Finding|SIMPLE_SEGMENT|5337,5346|false|false|false|C0442739||unchanged
Finding|Intellectual Product|SIMPLE_SEGMENT|5387,5393|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Substance|SIMPLE_SEGMENT|5407,5413|false|false|false|C0302908|Liquid substance|fluids
Finding|Body Substance|SIMPLE_SEGMENT|5407,5413|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5407,5413|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Organic Chemical|SIMPLE_SEGMENT|5418,5425|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5418,5425|false|false|false|C0591139|Bactrim|bactrim
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5454,5460|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5454,5474|true|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|SIMPLE_SEGMENT|5461,5474|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|SIMPLE_SEGMENT|5461,5474|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|SIMPLE_SEGMENT|5461,5474|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Procedure|Health Care Activity|SIMPLE_SEGMENT|5479,5483|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5479,5483|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Finding|Classification|SIMPLE_SEGMENT|5534,5544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5534,5544|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5545,5550|false|false|false|C1874451|Basis|basis
Finding|Functional Concept|SIMPLE_SEGMENT|5545,5550|false|false|false|C1527178|Basis - conceptual entity|basis
Finding|Finding|SIMPLE_SEGMENT|5555,5561|false|false|false|C0034359|Pyuria|Pyuria
Anatomy|Cell|SIMPLE_SEGMENT|5574,5577|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5590,5598|false|false|false|C0014894|Esterases|esterase
Drug|Enzyme|SIMPLE_SEGMENT|5590,5598|false|false|false|C0014894|Esterases|esterase
Procedure|Health Care Activity|SIMPLE_SEGMENT|5608,5617|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Functional Concept|SIMPLE_SEGMENT|5640,5648|true|false|false|C1510439|bacteria aspects|bacteria
Finding|Sign or Symptom|SIMPLE_SEGMENT|5664,5671|false|false|false|C0085624|Burning sensation|burning
Finding|Sign or Symptom|SIMPLE_SEGMENT|5672,5679|false|false|false|C0013428|Dysuria|dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|5692,5708|false|false|false|C0751534|Syncopal Episode|syncopal episode
Finding|Mental Process|SIMPLE_SEGMENT|5716,5723|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5729,5732|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5729,5732|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5729,5732|false|false|false|C0077906|urinastatin|UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|5729,5732|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Finding|Conceptual Entity|SIMPLE_SEGMENT|5734,5743|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|5734,5743|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5734,5743|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5734,5743|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Organic Chemical|SIMPLE_SEGMENT|5750,5757|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5750,5757|false|false|false|C0591139|Bactrim|bactrim
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5821,5833|false|false|false|C0023518|Leukocytosis|Leukocytosis
Finding|Finding|SIMPLE_SEGMENT|5821,5833|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Anatomy|Cell|SIMPLE_SEGMENT|5839,5842|false|false|false|C0023516|Leukocytes|WBC
Finding|Finding|SIMPLE_SEGMENT|5854,5860|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5854,5860|false|true|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Mental Process|SIMPLE_SEGMENT|5868,5875|false|true|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5884,5887|false|false|false|C0042029|Urinary tract infection|UTI
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5884,5887|false|false|false|C0077906|urinastatin|UTI
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5884,5887|false|false|false|C0077906|urinastatin|UTI
Finding|Gene or Genome|SIMPLE_SEGMENT|5884,5887|false|false|false|C1412376;C5780748|AMBP gene;AMBP wt Allele|UTI
Drug|Organic Chemical|SIMPLE_SEGMENT|5913,5920|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5913,5920|false|false|false|C0591139|Bactrim|bactrim
Finding|Idea or Concept|SIMPLE_SEGMENT|5924,5929|false|false|false|C1552828|Table Frame - above|above
Finding|Finding|SIMPLE_SEGMENT|5934,5942|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|INACTIVE
Finding|Idea or Concept|SIMPLE_SEGMENT|5934,5942|false|false|false|C1547420;C1608263;C1608264;C3244313;C3834263;C3890554|Certificate Status - Inactive;Edit Status - Inactive;Immunization Registry Status - Inactive;Inactive - answer to question;Inactive Healthcare Coverage;Physical Inactivity|INACTIVE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5954,5960|false|false|false|C0002871|Anemia|Anemia
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5962,5965|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5962,5965|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5998,6006|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|5998,6006|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6020,6024|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6020,6024|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6020,6024|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6020,6024|false|false|false|C0337439|Iron measurement|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6020,6032|false|false|false|C2079295|iron studies|Iron studies
Procedure|Research Activity|SIMPLE_SEGMENT|6025,6032|false|false|false|C0947630|Scientific Study|studies
Finding|Gene or Genome|SIMPLE_SEGMENT|6034,6037|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Drug|Organic Chemical|SIMPLE_SEGMENT|6043,6049|false|false|false|C0178638|folate|Folate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6043,6049|false|false|false|C0178638|folate|Folate
Drug|Vitamin|SIMPLE_SEGMENT|6043,6049|false|false|false|C0178638|folate|Folate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6043,6049|false|false|false|C0523631|Folic acid measurement|Folate
Finding|Finding|SIMPLE_SEGMENT|6055,6075|false|false|false|C0442816||within normal limits
Finding|Functional Concept|SIMPLE_SEGMENT|6069,6075|false|false|false|C0439801|Limited (extensiveness)|limits
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6080,6083|false|false|false|C0020538|Hypertensive disease|HTN
Finding|Idea or Concept|SIMPLE_SEGMENT|6089,6093|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6089,6093|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6089,6093|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6094,6104|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6094,6104|false|false|false|C0065374|lisinopril|lisinopril
Finding|Mental Process|SIMPLE_SEGMENT|6144,6151|false|false|false|C0542559|contextual factors|setting
Finding|Sign or Symptom|SIMPLE_SEGMENT|6159,6166|false|false|false|C0039070|Syncope|syncope
Event|Activity|SIMPLE_SEGMENT|6170,6175|false|false|false|C1705178|Order (action)|order
Finding|Classification|SIMPLE_SEGMENT|6170,6175|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Idea or Concept|SIMPLE_SEGMENT|6170,6175|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Intellectual Product|SIMPLE_SEGMENT|6170,6175|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|6170,6175|false|false|false|C1373200|Order [PK]|order
Finding|Finding|SIMPLE_SEGMENT|6208,6215|false|false|false|C4036057|Too low|too low
Finding|Finding|SIMPLE_SEGMENT|6212,6215|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|6212,6215|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6220,6234|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Finding|Idea or Concept|SIMPLE_SEGMENT|6246,6250|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|6246,6250|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6246,6250|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6251,6263|false|false|false|C0040165|levothyroxine|levothyroxin
Drug|Hormone|SIMPLE_SEGMENT|6251,6263|false|false|false|C0040165|levothyroxine|levothyroxin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6251,6263|false|false|false|C0040165|levothyroxine|levothyroxin
Event|Activity|SIMPLE_SEGMENT|6282,6286|false|false|false|C1947933|care activity|CARE
Finding|Finding|SIMPLE_SEGMENT|6282,6286|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Finding|Intellectual Product|SIMPLE_SEGMENT|6282,6286|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|CARE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6294,6298|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6294,6298|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6294,6298|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6294,6298|false|false|false|C0337439|Iron measurement|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6294,6306|false|false|false|C2079295|iron studies|Iron studies
Procedure|Research Activity|SIMPLE_SEGMENT|6299,6306|false|false|false|C0947630|Scientific Study|studies
Finding|Gene or Genome|SIMPLE_SEGMENT|6312,6315|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Drug|Organic Chemical|SIMPLE_SEGMENT|6326,6332|false|false|false|C0178638|folate|Folate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6326,6332|false|false|false|C0178638|folate|Folate
Drug|Vitamin|SIMPLE_SEGMENT|6326,6332|false|false|false|C0178638|folate|Folate
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6326,6332|false|false|false|C0523631|Folic acid measurement|Folate
Procedure|Health Care Activity|SIMPLE_SEGMENT|6355,6359|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6355,6359|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|Echo
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6372,6383|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6372,6383|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6372,6383|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|6372,6396|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6387,6396|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6398,6408|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6398,6408|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6422,6435|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6422,6435|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6422,6435|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6422,6435|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Finding|Body Substance|SIMPLE_SEGMENT|6453,6462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6453,6462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6453,6462|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6453,6462|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6453,6474|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6463,6474|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6463,6474|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6463,6474|false|false|false|C4284232|Medications|Medications
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6479,6492|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|SIMPLE_SEGMENT|6479,6492|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|SIMPLE_SEGMENT|6479,6492|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6479,6492|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6500,6506|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6520,6526|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6551,6561|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6551,6561|false|false|false|C0065374|lisinopril|lisinopril
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6568,6574|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6588,6594|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6622,6628|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6633,6640|false|false|false|C0807726|refill|Refills
Drug|Antibiotic|SIMPLE_SEGMENT|6648,6664|false|false|false|C0038689|sulfamethoxazole|sulfamethoxazole
Drug|Organic Chemical|SIMPLE_SEGMENT|6648,6664|false|false|false|C0038689|sulfamethoxazole|sulfamethoxazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6648,6677|false|false|false|C0041044|Trimethoprim-Sulfamethoxazole Combination|sulfamethoxazole-trimethoprim
Drug|Antibiotic|SIMPLE_SEGMENT|6665,6677|false|false|false|C0041041|trimethoprim|trimethoprim
Drug|Organic Chemical|SIMPLE_SEGMENT|6665,6677|false|false|false|C0041041|trimethoprim|trimethoprim
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6689,6695|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6710,6716|false|false|false|C0039225|Tablet Dosage Form|Tablet
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6720,6723|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6720,6723|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6720,6723|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6720,6723|false|false|false|C1332410|BID gene|BID
Finding|Finding|SIMPLE_SEGMENT|6725,6732|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6727,6732|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|SIMPLE_SEGMENT|6735,6738|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|6735,6738|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6760,6766|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6771,6778|false|false|false|C0807726|refill|Refills
Drug|Food|SIMPLE_SEGMENT|6786,6790|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Drug|Organic Chemical|SIMPLE_SEGMENT|6786,6790|false|false|false|C3257082;C4521129|Fish (substance);Fish extract|Fish
Finding|Gene or Genome|SIMPLE_SEGMENT|6786,6790|false|false|false|C1822711;C3274826|SH3PXD2A gene;SH3PXD2A wt Allele|Fish
Procedure|Molecular Biology Research Technique|SIMPLE_SEGMENT|6786,6790|false|false|false|C0162789|Fluorescent in Situ Hybridization|Fish
Drug|Organic Chemical|SIMPLE_SEGMENT|6786,6794|false|false|false|C0016157|fish oils|Fish Oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6786,6794|false|false|false|C0016157|fish oils|Fish Oil
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6791,6794|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Food|SIMPLE_SEGMENT|6791,6794|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Organic Chemical|SIMPLE_SEGMENT|6791,6794|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6791,6794|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|Oil
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6796,6800|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6796,6800|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|6796,6800|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|6796,6800|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6804,6811|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6804,6811|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6804,6811|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6804,6811|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|SIMPLE_SEGMENT|6804,6811|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|6804,6811|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6804,6811|false|false|false|C0201925|Calcium measurement|calcium
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6813,6817|false|false|false|C0226896|Oral cavity|Oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6813,6817|false|false|false|C1272919|Oral Dosage Form|Oral
Finding|Finding|SIMPLE_SEGMENT|6813,6817|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Functional Concept|SIMPLE_SEGMENT|6813,6817|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|Oral
Finding|Body Substance|SIMPLE_SEGMENT|6821,6830|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6821,6830|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6821,6830|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6821,6830|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6821,6842|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6821,6842|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6831,6842|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6831,6842|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|6844,6848|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6844,6848|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6844,6848|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|SIMPLE_SEGMENT|6851,6860|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6851,6860|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6851,6860|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6851,6860|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6851,6870|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6861,6870|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6861,6870|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6861,6870|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6861,6870|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6872,6889|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6880,6889|false|false|false|C0945731||diagnosis
Finding|Classification|SIMPLE_SEGMENT|6880,6889|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6880,6889|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6880,6889|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Sign or Symptom|SIMPLE_SEGMENT|6891,6898|false|false|false|C0039070|Syncope|Syncope
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6900,6909|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6900,6909|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6910,6919|false|false|false|C0011900|Diagnosis|diagnoses
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6921,6935|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6936,6948|false|false|false|C0020538|Hypertensive disease|Hypertension
Finding|Body Substance|SIMPLE_SEGMENT|6952,6961|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6952,6961|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6952,6961|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6952,6961|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6962,6971|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6962,6971|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6962,6971|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|6973,6979|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6973,6986|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|6973,6986|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6980,6986|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6980,6986|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|6988,6993|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|6998,7006|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7008,7030|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7008,7030|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7017,7030|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|7017,7030|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7032,7037|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|7032,7037|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7032,7037|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|7032,7037|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7032,7037|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|7032,7037|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7042,7053|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|7055,7063|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7055,7063|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|7055,7063|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7064,7070|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7064,7070|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|7072,7082|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|7072,7082|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|7072,7082|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|7072,7082|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|7085,7096|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|7085,7096|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|7101,7110|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7101,7110|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7101,7110|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7101,7110|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7101,7123|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7101,7123|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|7101,7123|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7111,7123|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7111,7123|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|7125,7129|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|SIMPLE_SEGMENT|7149,7157|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|7149,7157|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|7168,7172|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|7168,7172|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7168,7172|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Sign or Symptom|SIMPLE_SEGMENT|7248,7256|false|false|false|C0039070|Syncope|fainting
Finding|Idea or Concept|SIMPLE_SEGMENT|7304,7312|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7304,7315|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7318,7325|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7318,7331|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|7318,7331|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7318,7341|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7326,7331|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7332,7341|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|7332,7341|false|false|false|C3714514|Infection|infection
Drug|Antibiotic|SIMPLE_SEGMENT|7368,7378|false|false|false|C0003232|Antibiotics|antibiotic
Drug|Organic Chemical|SIMPLE_SEGMENT|7386,7393|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7386,7393|false|false|false|C0591139|Bactrim|Bactrim
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7401,7406|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|7401,7406|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7401,7412|false|false|false|C0039985|Plain chest X-ray|chest x-ray
Finding|Functional Concept|SIMPLE_SEGMENT|7407,7412|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|SIMPLE_SEGMENT|7407,7412|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7407,7412|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7407,7412|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Finding|Idea or Concept|SIMPLE_SEGMENT|7427,7435|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|SIMPLE_SEGMENT|7449,7457|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7449,7460|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7463,7472|true|false|false|C0032285|Pneumonia|pneumonia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7494,7499|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7494,7499|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|7494,7499|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7494,7506|false|false|false|C0232187|Cardiac rhythm type|heart rhythm
Finding|Finding|SIMPLE_SEGMENT|7500,7506|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|7500,7506|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|7538,7551|true|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|7538,7551|true|false|false|C0000769|teratologic|abnormalities
Finding|Intellectual Product|SIMPLE_SEGMENT|7560,7577|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|electrocardiogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7560,7577|false|false|false|C1623258|Electrocardiography|electrocardiogram
Finding|Functional Concept|SIMPLE_SEGMENT|7595,7602|true|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7610,7615|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|7610,7615|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|7617,7625|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|7617,7625|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|7617,7625|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|7617,7625|false|false|false|C0033095||pressure
Finding|Intellectual Product|SIMPLE_SEGMENT|7635,7641|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|SIMPLE_SEGMENT|7661,7671|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7661,7671|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7661,7671|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7680,7685|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7680,7685|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|7680,7685|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Idea or Concept|SIMPLE_SEGMENT|7698,7708|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|SIMPLE_SEGMENT|7698,7708|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7710,7724|false|false|false|C0013516|Echocardiography|echocardiogram
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7781,7790|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7781,7790|false|false|false|C0012634|Disease|condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|7781,7790|false|false|false|C1705253|Logical Condition|condition
Finding|Idea or Concept|SIMPLE_SEGMENT|7833,7837|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7833,7837|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7833,7837|false|false|false|C1553498|home health encounter|home
Finding|Functional Concept|SIMPLE_SEGMENT|7854,7861|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7880,7891|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7880,7891|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7880,7891|false|false|false|C4284232|Medications|medications
Finding|Finding|SIMPLE_SEGMENT|7894,7897|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|NEW
Finding|Idea or Concept|SIMPLE_SEGMENT|7894,7897|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|NEW
Drug|Organic Chemical|SIMPLE_SEGMENT|7901,7908|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7901,7908|false|false|false|C0591139|Bactrim|Bactrim
Event|Activity|SIMPLE_SEGMENT|7909,7915|false|false|false|C1705764|Doubling|double
Finding|Functional Concept|SIMPLE_SEGMENT|7909,7915|false|false|false|C0205173|Double (qualifier value)|double
Finding|Idea or Concept|SIMPLE_SEGMENT|7916,7924|false|false|false|C0808080|Strength (attribute)|strength
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7925,7928|false|false|false|C0039225|Tablet Dosage Form|tab
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|7932,7935|false|false|false|C0039225|Tablet Dosage Form|tab
Finding|Functional Concept|SIMPLE_SEGMENT|7936,7944|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7939,7944|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|7939,7944|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7984,7991|false|false|false|C0042027|Urinary tract|urinary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7984,7997|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Anatomy|Body System|SIMPLE_SEGMENT|7984,7997|false|false|false|C0042027;C1508753|Urinary system;Urinary tract|urinary tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7984,8007|false|false|false|C0042029|Urinary tract infection|urinary tract infection
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7992,7997|false|false|false|C1185740|Tract|tract
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7998,8007|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|SIMPLE_SEGMENT|7998,8007|false|false|false|C3714514|Infection|infection
Finding|Finding|SIMPLE_SEGMENT|8021,8030|false|false|false|C0392756;C0442797|Decreasing;Reduced|DECREASED
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8031,8041|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8031,8041|false|false|false|C0065374|lisinopril|Lisinopril
Finding|Functional Concept|SIMPLE_SEGMENT|8050,8058|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|8053,8058|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|8053,8058|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Functional Concept|SIMPLE_SEGMENT|8083,8089|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|8083,8089|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|SIMPLE_SEGMENT|8083,8092|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|SIMPLE_SEGMENT|8083,8092|false|false|false|C1522577|follow-up|follow-up
Event|Activity|SIMPLE_SEGMENT|8093,8105|false|false|false|C0003629|Appointments|appointments
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8165,8179|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Intellectual Product|SIMPLE_SEGMENT|8221,8226|false|false|false|C3463807|Video Media|video
Finding|Functional Concept|SIMPLE_SEGMENT|8227,8234|false|false|false|C1706486;C4521686|Swallow (administration method);Swallow - dosing instruction imperative|swallow
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8227,8240|false|false|false|C3888792|Swallow study|swallow study
Finding|Intellectual Product|SIMPLE_SEGMENT|8235,8240|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|SIMPLE_SEGMENT|8235,8240|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Finding|Idea or Concept|SIMPLE_SEGMENT|8260,8268|false|false|false|C3887511|Evidence|evidence
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|8339,8351|false|false|false|C0184625||regular diet
Drug|Food|SIMPLE_SEGMENT|8347,8351|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Finding|Functional Concept|SIMPLE_SEGMENT|8347,8351|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|8347,8351|false|false|false|C0012159|Diet therapy|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|8355,8363|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8364,8376|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8364,8376|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

