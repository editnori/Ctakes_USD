 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|40,49|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|40,49|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|40,54|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|74,83|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|74,83|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|74,83|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|74,88|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|106,111|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|130,133|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|130,133|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|141,148|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|141,148|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|150,158|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|161,170|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|161,170|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|161,170|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Body Substance|SIMPLE_SEGMENT|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|173,180|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|181,189|false|false|false|||recorded
Attribute|Clinical Attribute|SIMPLE_SEGMENT|209,218|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|209,218|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|209,218|true|false|false|C0020517|Hypersensitivity|Allergies
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|222,227|false|false|false|C0013227|Pharmaceutical Preparations|Drugs
Event|Event|SIMPLE_SEGMENT|222,227|false|false|false|||Drugs
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|222,227|false|false|false|C3687832|Drugs - dental services|Drugs
Event|Event|SIMPLE_SEGMENT|230,239|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|230,239|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|248,263|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|254,263|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|254,263|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|254,263|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|265,274|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|SIMPLE_SEGMENT|265,285|false|false|false|C0000731|Abdomen distended|Abdominal distention
Event|Event|SIMPLE_SEGMENT|275,285|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|275,285|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|275,285|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|286,290|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|286,290|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|286,290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|286,290|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|286,300|false|false|false|C3499958|Pain and Fever|pain and fever
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|286,300|false|false|false|C3499958|Pain and Fever|pain and fever
Event|Event|SIMPLE_SEGMENT|295,300|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|295,300|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|295,300|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Classification|SIMPLE_SEGMENT|303,308|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|309,317|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|309,317|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|321,339|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|330,339|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|330,339|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|330,339|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|330,339|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|330,339|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|341,353|false|false|false|||Paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|341,353|false|false|false|C0034115|Paracentesis|Paracentesis
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|359,369|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|SIMPLE_SEGMENT|359,369|false|false|false|||diagnostic
Finding|Functional Concept|SIMPLE_SEGMENT|359,369|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|SIMPLE_SEGMENT|359,369|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|359,369|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Drug|Organic Chemical|SIMPLE_SEGMENT|380,391|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|380,391|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|SIMPLE_SEGMENT|380,391|false|false|false|||therapeutic
Finding|Functional Concept|SIMPLE_SEGMENT|380,391|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|SIMPLE_SEGMENT|380,391|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|380,391|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|SIMPLE_SEGMENT|396,403|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|396,403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|396,403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|396,403|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|396,406|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|396,422|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|396,422|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|407,414|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|407,414|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|407,422|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|415,422|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|442,451|false|false|false|||diagnosed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|452,471|false|false|false|C0019187|Hepatitis, Alcoholic|alcoholic hepatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|462,471|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|SIMPLE_SEGMENT|462,471|false|false|false|||hepatitis
Event|Event|SIMPLE_SEGMENT|473,483|false|false|false|||persistent
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|485,492|false|false|false|C0003962|Ascites|ascites
Event|Event|SIMPLE_SEGMENT|485,492|false|false|false|||ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|485,492|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|SIMPLE_SEGMENT|509,515|false|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|509,515|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|520,532|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|520,532|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|520,532|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Event|Event|SIMPLE_SEGMENT|550,559|false|false|false|||atributed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|567,576|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|SIMPLE_SEGMENT|567,576|false|false|false|||hepatitis
Event|Event|SIMPLE_SEGMENT|581,590|false|false|false|||presented
Finding|Idea or Concept|SIMPLE_SEGMENT|610,619|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Anatomy|Body Location or Region|SIMPLE_SEGMENT|620,629|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|620,640|false|false|false|C0000731|Abdomen distended|abdominal distention
Event|Event|SIMPLE_SEGMENT|630,640|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|630,640|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|630,640|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|642,646|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|642,646|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|642,646|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Pathologic Function|SIMPLE_SEGMENT|652,668|false|false|false|C0476474|Persistent fever|persistent fever
Event|Event|SIMPLE_SEGMENT|663,668|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|663,668|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|663,668|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|675,681|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|682,688|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|682,688|true|false|false|C0085593|Chills|chills
Finding|Intellectual Product|SIMPLE_SEGMENT|697,708|false|false|false|C4084908|Have Sweats|have sweats
Event|Event|SIMPLE_SEGMENT|702,708|false|false|false|||sweats
Finding|Body Substance|SIMPLE_SEGMENT|702,708|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|SIMPLE_SEGMENT|702,708|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Event|Event|SIMPLE_SEGMENT|728,737|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|728,737|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|748,753|false|false|false|||tried
Event|Event|SIMPLE_SEGMENT|769,778|false|false|false|||compliant
Finding|Individual Behavior|SIMPLE_SEGMENT|769,778|false|false|false|C1321605|Compliance behavior|compliant
Finding|Finding|SIMPLE_SEGMENT|788,791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|788,791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Drug|Food|SIMPLE_SEGMENT|799,803|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|SIMPLE_SEGMENT|799,803|false|false|false|||diet
Finding|Functional Concept|SIMPLE_SEGMENT|799,803|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|799,803|false|false|false|C0012159|Diet therapy|diet
Drug|Substance|SIMPLE_SEGMENT|809,814|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|809,814|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|809,826|false|false|false|C0204700|Fluid restriction|fluid restriction
Event|Event|SIMPLE_SEGMENT|815,826|false|false|false|||restriction
Finding|Functional Concept|SIMPLE_SEGMENT|815,826|false|false|false|C0443288|Restricted|restriction
Event|Event|SIMPLE_SEGMENT|832,838|false|false|false|||denies
Finding|Finding|SIMPLE_SEGMENT|843,852|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Finding|Functional Concept|SIMPLE_SEGMENT|843,852|false|false|false|C0442805;C5236002|Increase;Increased (finding)|increased
Drug|Substance|SIMPLE_SEGMENT|853,858|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|853,858|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|853,858|true|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Biologically Active Substance|SIMPLE_SEGMENT|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|862,868|true|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|862,868|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|862,868|true|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|862,868|true|false|false|C0337443|Sodium measurement|sodium
Event|Event|SIMPLE_SEGMENT|870,876|false|false|false|||intake
Finding|Functional Concept|SIMPLE_SEGMENT|870,876|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|SIMPLE_SEGMENT|870,876|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|SIMPLE_SEGMENT|882,889|false|false|false|||reports
Event|Event|SIMPLE_SEGMENT|890,898|false|false|false|||sobriety
Finding|Individual Behavior|SIMPLE_SEGMENT|890,898|false|false|false|C0680686|sobriety|sobriety
Drug|Organic Chemical|SIMPLE_SEGMENT|904,911|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|904,911|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Event|Event|SIMPLE_SEGMENT|904,911|false|false|false|||alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|904,911|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Event|Event|SIMPLE_SEGMENT|939,946|false|false|false|||febrile
Finding|Sign or Symptom|SIMPLE_SEGMENT|939,946|false|false|false|C0015967|Fever|febrile
Event|Event|SIMPLE_SEGMENT|951,957|false|false|false|||tender
Event|Event|SIMPLE_SEGMENT|961,970|false|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|961,970|false|false|false|C0030247|Palpation|palpation
Event|Event|SIMPLE_SEGMENT|983,991|false|false|false|||referred
Finding|Idea or Concept|SIMPLE_SEGMENT|1020,1027|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|SIMPLE_SEGMENT|1028,1033|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1028,1039|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|1028,1039|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|SIMPLE_SEGMENT|1034,1039|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|1034,1039|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1034,1039|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|1080,1084|false|false|false|||temp
Finding|Gene or Genome|SIMPLE_SEGMENT|1080,1084|false|false|false|C1823816|C1orf210 gene|temp
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1080,1084|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|temp
Event|Event|SIMPLE_SEGMENT|1085,1094|false|false|false|||increased
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1112,1117|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|1112,1117|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|1112,1117|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1112,1117|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|1112,1117|false|false|false|C0034107|Pulse taking|pulse
Event|Event|SIMPLE_SEGMENT|1118,1122|false|false|false|||came
Drug|Organic Chemical|SIMPLE_SEGMENT|1146,1152|false|false|false|C0699194|Ativan|Ativan
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1146,1152|false|false|false|C0699194|Ativan|Ativan
Drug|Organic Chemical|SIMPLE_SEGMENT|1167,1175|false|false|false|C0026549|morphine|morphine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1167,1175|false|false|false|C0026549|morphine|morphine
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1191,1195|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1191,1195|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1191,1195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1191,1195|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|1197,1204|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1197,1204|false|false|false|C0699142|Tylenol|tylenol
Event|Event|SIMPLE_SEGMENT|1197,1204|false|false|false|||tylenol
Event|Event|SIMPLE_SEGMENT|1220,1225|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|1220,1225|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|1220,1225|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Drug|Organic Chemical|SIMPLE_SEGMENT|1227,1238|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1227,1238|false|false|false|C0061851|ondansetron|ondansetron
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1253,1259|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|1253,1259|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1253,1259|false|false|false|C0027497|Nausea|nausea
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1292,1299|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|1292,1299|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|1292,1299|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1317,1327|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|SIMPLE_SEGMENT|1317,1327|false|false|false|||diagnostic
Finding|Functional Concept|SIMPLE_SEGMENT|1317,1327|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|SIMPLE_SEGMENT|1317,1327|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1317,1327|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Event|Event|SIMPLE_SEGMENT|1329,1341|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1329,1341|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|SIMPLE_SEGMENT|1350,1357|false|false|false|||samples
Event|Event|SIMPLE_SEGMENT|1373,1377|false|false|false|||lost
Event|Event|SIMPLE_SEGMENT|1388,1395|false|false|false|||treated
Drug|Antibiotic|SIMPLE_SEGMENT|1401,1412|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|1401,1412|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|1401,1412|false|false|false|||ceftriaxone
Event|Event|SIMPLE_SEGMENT|1419,1421|false|false|false|||x1
Finding|Finding|SIMPLE_SEGMENT|1426,1434|false|false|false|C0332149|Possible|possible
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1435,1438|false|true|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1435,1438|false|true|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1435,1438|false|true|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|1435,1438|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|1435,1438|false|true|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1435,1438|false|true|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|SIMPLE_SEGMENT|1449,1457|false|false|false|||admitted
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1461,1469|false|false|false|C0013227|Pharmaceutical Preparations|Medicine
Event|Event|SIMPLE_SEGMENT|1482,1492|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|1482,1492|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|1482,1492|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|1512,1519|false|false|false|||samples
Event|Event|SIMPLE_SEGMENT|1525,1530|false|false|false|||found
Event|Event|SIMPLE_SEGMENT|1541,1548|false|false|false|||arrived
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1556,1561|false|false|false|C3714591|Floor (anatomic)|floor
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|1576,1581|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1586,1590|false|false|false|C2713234||mood
Event|Event|SIMPLE_SEGMENT|1586,1590|false|false|false|||mood
Finding|Conceptual Entity|SIMPLE_SEGMENT|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Finding|SIMPLE_SEGMENT|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Finding|Mental Process|SIMPLE_SEGMENT|1586,1590|false|false|false|C0026516;C3889585;C5444612|Mood (attribute);Mood (psychological function);mood (physical finding)|mood
Event|Event|SIMPLE_SEGMENT|1594,1600|false|false|false|||labile
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1612,1617|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|1618,1625|false|false|false|||tearful
Finding|Finding|SIMPLE_SEGMENT|1618,1625|false|false|false|C0424109|Weepiness|tearful
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1634,1639|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|SIMPLE_SEGMENT|1634,1639|false|false|false|||times
Event|Event|SIMPLE_SEGMENT|1640,1648|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|1640,1648|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|1659,1663|false|false|false|||seem
Event|Event|SIMPLE_SEGMENT|1664,1677|false|false|false|||uncomfortable
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|1690,1698|true|false|false|C0009676|Confusion|confused
Event|Event|SIMPLE_SEGMENT|1690,1698|false|false|false|||confused
Finding|Finding|SIMPLE_SEGMENT|1690,1698|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Finding|Intellectual Product|SIMPLE_SEGMENT|1690,1698|true|false|false|C0683369;C1547301|Clouded consciousness;Precaution Code - Confused|confused
Event|Event|SIMPLE_SEGMENT|1713,1728|false|false|false|||encephalopathic
Event|Event|SIMPLE_SEGMENT|1734,1740|false|false|false|||denies
Drug|Organic Chemical|SIMPLE_SEGMENT|1741,1746|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1741,1746|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|1741,1746|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|1741,1746|true|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|1748,1755|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|1748,1755|true|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|1758,1766|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1758,1766|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1758,1766|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1771,1775|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|SIMPLE_SEGMENT|1771,1775|false|false|false|||rash
Finding|Pathologic Function|SIMPLE_SEGMENT|1771,1775|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|SIMPLE_SEGMENT|1771,1775|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Finding|SIMPLE_SEGMENT|1794,1803|false|false|false|C0392756;C0442797|Decreasing;Reduced|decreased
Event|Event|SIMPLE_SEGMENT|1804,1807|false|false|false|||UOP
Event|Event|SIMPLE_SEGMENT|1836,1842|false|false|false|||Review
Finding|Idea or Concept|SIMPLE_SEGMENT|1836,1842|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Intellectual Product|SIMPLE_SEGMENT|1836,1842|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|Review
Finding|Functional Concept|SIMPLE_SEGMENT|1836,1845|false|false|false|C0699752|Review of|Review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1836,1853|false|false|false|C0488564;C0488565||Review of Systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|1836,1853|false|false|false|C0489633|Review of systems (procedure)|Review of Systems
Event|Event|SIMPLE_SEGMENT|1846,1853|false|false|false|||Systems
Finding|Functional Concept|SIMPLE_SEGMENT|1846,1853|false|false|false|C0449913|System|Systems
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1865,1868|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|SIMPLE_SEGMENT|1865,1868|false|false|false|||HPI
Finding|Finding|SIMPLE_SEGMENT|1865,1868|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|SIMPLE_SEGMENT|1865,1868|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|SIMPLE_SEGMENT|1875,1881|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|1882,1888|false|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1882,1888|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1890,1896|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|1897,1905|false|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|1897,1905|true|false|false|C0018681|Headache|headache
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|1907,1912|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|1907,1912|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|SIMPLE_SEGMENT|1907,1912|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1907,1912|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Event|Event|SIMPLE_SEGMENT|1913,1923|false|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|1913,1923|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1913,1923|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|1925,1935|false|false|false|||rhinorrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1925,1935|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Event|Event|SIMPLE_SEGMENT|1940,1950|false|false|false|||congestion
Finding|Pathologic Function|SIMPLE_SEGMENT|1940,1950|false|false|false|C0700148|Congestion|congestion
Event|Event|SIMPLE_SEGMENT|1952,1958|false|false|false|||Denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1959,1964|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1959,1964|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1959,1969|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1959,1969|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1965,1969|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1965,1969|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1965,1969|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1965,1969|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1973,1982|false|false|false|||tightness
Event|Event|SIMPLE_SEGMENT|1984,1996|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|1984,1996|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|1999,2005|false|false|false|||Denies
Drug|Organic Chemical|SIMPLE_SEGMENT|2006,2011|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2006,2011|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2006,2011|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2006,2011|false|false|false|C0010200|Coughing|cough
Event|Event|SIMPLE_SEGMENT|2013,2022|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2013,2032|true|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|2013,2032|true|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|2026,2032|false|false|false|C0225386|Breath|breath
Event|Event|SIMPLE_SEGMENT|2037,2044|false|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2037,2044|true|false|false|C0043144|Wheezing|wheezes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2053,2059|false|false|false|C4255480||nausea
Event|Event|SIMPLE_SEGMENT|2053,2059|false|false|false|||nausea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2053,2059|false|false|false|C0027497|Nausea|nausea
Event|Event|SIMPLE_SEGMENT|2062,2070|false|false|false|||vomiting
Finding|Sign or Symptom|SIMPLE_SEGMENT|2062,2070|false|false|false|C0042963|Vomiting|vomiting
Event|Event|SIMPLE_SEGMENT|2072,2080|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|2072,2080|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|2072,2080|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|SIMPLE_SEGMENT|2082,2094|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|2082,2094|false|false|false|C0009806|Constipation|constipation
Event|Event|SIMPLE_SEGMENT|2106,2112|false|false|false|||change
Finding|Functional Concept|SIMPLE_SEGMENT|2106,2112|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2106,2112|true|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|SIMPLE_SEGMENT|2106,2115|true|false|false|C0392747|Changing|change in
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2116,2121|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2126,2133|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2126,2133|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Event|Event|SIMPLE_SEGMENT|2126,2133|false|false|false|||bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2126,2133|false|false|false|C0872388|Procedures on bladder|bladder
Event|Event|SIMPLE_SEGMENT|2134,2140|false|false|false|||habits
Finding|Finding|SIMPLE_SEGMENT|2134,2140|false|false|false|C0018464;C2242848|Behaviorial Habits;habits (history)|habits
Finding|Individual Behavior|SIMPLE_SEGMENT|2134,2140|false|false|false|C0018464;C2242848|Behaviorial Habits;habits (history)|habits
Event|Event|SIMPLE_SEGMENT|2145,2152|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|2145,2152|true|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|2154,2160|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2161,2172|false|false|false|||arthralgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2161,2172|true|false|false|C0003862|Arthralgia|arthralgias
Event|Event|SIMPLE_SEGMENT|2176,2184|false|false|false|||myalgias
Finding|Sign or Symptom|SIMPLE_SEGMENT|2176,2184|true|false|false|C0231528|Myalgia|myalgias
Event|Event|SIMPLE_SEGMENT|2187,2193|false|false|false|||Denies
Event|Event|SIMPLE_SEGMENT|2194,2200|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2194,2200|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Anatomy|Body System|SIMPLE_SEGMENT|2204,2208|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2204,2208|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2204,2208|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|2204,2208|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2204,2208|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|SIMPLE_SEGMENT|2204,2218|true|false|false|C0150077;C4048181|Broken skin;Impaired skin integrity|skin breakdown
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2209,2218|false|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Event|Event|SIMPLE_SEGMENT|2209,2218|false|false|false|||breakdown
Finding|Organism Function|SIMPLE_SEGMENT|2209,2218|false|false|false|C0699900|Catabolism|breakdown
Event|Event|SIMPLE_SEGMENT|2223,2231|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|2223,2231|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2223,2231|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2232,2240|true|false|false|C0030554|Paresthesia|tingling
Event|Event|SIMPLE_SEGMENT|2232,2240|false|false|false|||tingling
Finding|Sign or Symptom|SIMPLE_SEGMENT|2232,2240|true|false|false|C2242996|Has tingling sensation|tingling
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2245,2256|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|2261,2269|false|false|false|||feelings
Finding|Intellectual Product|SIMPLE_SEGMENT|2261,2269|true|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|SIMPLE_SEGMENT|2261,2269|true|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2273,2283|true|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|SIMPLE_SEGMENT|2273,2283|false|false|false|||depression
Finding|Functional Concept|SIMPLE_SEGMENT|2273,2283|true|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|2273,2283|true|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2287,2294|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|2287,2294|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|2287,2294|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|SIMPLE_SEGMENT|2296,2305|false|false|false|C5425799|All other|All other
Event|Event|SIMPLE_SEGMENT|2307,2313|false|false|false|||review
Finding|Idea or Concept|SIMPLE_SEGMENT|2307,2313|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Intellectual Product|SIMPLE_SEGMENT|2307,2313|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|review
Finding|Functional Concept|SIMPLE_SEGMENT|2307,2316|false|false|false|C0699752|Review of|review of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2307,2324|false|false|false|C0488564;C0488565||review of systems
Procedure|Health Care Activity|SIMPLE_SEGMENT|2307,2324|false|false|false|C0489633|Review of systems (procedure)|review of systems
Event|Event|SIMPLE_SEGMENT|2317,2324|false|false|false|||systems
Finding|Functional Concept|SIMPLE_SEGMENT|2317,2324|false|false|false|C0449913|System|systems
Event|Event|SIMPLE_SEGMENT|2325,2333|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|2325,2333|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|2325,2333|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2325,2333|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|SIMPLE_SEGMENT|2340,2360|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|2345,2352|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|2345,2352|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|2345,2352|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|2345,2352|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2345,2352|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|2345,2360|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2353,2360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2353,2360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2353,2360|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Drug|Organic Chemical|SIMPLE_SEGMENT|2364,2371|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2364,2371|false|false|false|C0001962;C0001975|Alcohols;ethanol|Alcohol
Finding|Intellectual Product|SIMPLE_SEGMENT|2364,2371|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|Alcohol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2364,2377|false|false|false|C0085762|Alcohol abuse|Alcohol abuse
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2372,2377|false|false|false|C0013146|Drug abuse|abuse
Event|Event|SIMPLE_SEGMENT|2372,2377|false|false|false|||abuse
Event|Event|SIMPLE_SEGMENT|2372,2377|false|false|false|C1546935|Abuse|abuse
Finding|Finding|SIMPLE_SEGMENT|2372,2377|false|false|false|C0562381|Victim of abuse (finding)|abuse
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2382,2401|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2392,2401|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|SIMPLE_SEGMENT|2392,2401|false|false|false|||hepatitis
Finding|Pathologic Function|SIMPLE_SEGMENT|2408,2424|false|false|false|C0476474|Persistent fever|persistent fever
Event|Event|SIMPLE_SEGMENT|2419,2424|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|2419,2424|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|2419,2424|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2429,2441|false|false|false|C0023518|Leukocytosis|leukocytosis
Event|Event|SIMPLE_SEGMENT|2429,2441|false|false|false|||leukocytosis
Finding|Finding|SIMPLE_SEGMENT|2429,2441|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2444,2451|false|false|false|C0003962|Ascites|Ascites
Event|Event|SIMPLE_SEGMENT|2444,2451|false|false|false|||Ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|2444,2451|false|false|false|C5441966|Peritoneal Effusion|Ascites
Event|Event|SIMPLE_SEGMENT|2455,2462|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|2455,2462|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|2455,2462|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|SIMPLE_SEGMENT|2455,2472|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2463,2472|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2468,2472|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|2468,2472|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|2468,2472|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|2468,2472|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|SIMPLE_SEGMENT|2476,2482|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2476,2490|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|2483,2490|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2483,2490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2483,2490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2483,2490|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2496,2502|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2496,2502|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2496,2502|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2496,2502|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2496,2510|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|2503,2510|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2503,2510|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2503,2510|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2503,2510|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Idea or Concept|SIMPLE_SEGMENT|2514,2520|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2526,2532|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|2526,2532|false|false|false|||cancer
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2534,2537|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2534,2537|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|2534,2537|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|SIMPLE_SEGMENT|2534,2537|false|false|false|||age
Finding|Classification|SIMPLE_SEGMENT|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2549,2555|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|SIMPLE_SEGMENT|2549,2563|true|false|false|C0241889|Family Medical History|family history
Finding|Finding|SIMPLE_SEGMENT|2549,2566|true|false|false|C0241889|Family Medical History|family history of
Event|Event|SIMPLE_SEGMENT|2556,2563|false|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|2556,2563|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|2556,2566|true|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|2556,2580|true|false|false|C0455550||history of liver disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2567,2572|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2567,2572|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2567,2572|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|2567,2572|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Finding|Finding|SIMPLE_SEGMENT|2567,2572|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|2567,2572|true|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2567,2580|true|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2573,2580|true|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|2573,2580|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|2594,2603|false|false|false|||relatives
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2609,2619|false|false|false|C0001973|Alcoholic Intoxication, Chronic|alcoholism
Event|Event|SIMPLE_SEGMENT|2609,2619|false|false|false|||alcoholism
Event|Event|SIMPLE_SEGMENT|2624,2632|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2624,2632|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2624,2632|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2624,2632|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2624,2637|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2624,2637|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2633,2637|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2633,2637|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2633,2637|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2639,2647|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|2639,2647|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2639,2647|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2639,2647|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2639,2652|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2639,2652|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|2648,2652|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2648,2652|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2648,2652|false|false|false|C0582103|Medical Examination|Exam
Event|Event|SIMPLE_SEGMENT|2656,2665|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|2656,2665|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Event|Event|SIMPLE_SEGMENT|2669,2672|false|false|false|||GEN
Finding|Classification|SIMPLE_SEGMENT|2669,2672|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Finding|Gene or Genome|SIMPLE_SEGMENT|2669,2672|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|GEN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2674,2677|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2674,2677|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2674,2677|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2674,2677|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2674,2677|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2679,2692|false|false|false|C0233472|Labile affect|labile affect
Event|Event|SIMPLE_SEGMENT|2686,2692|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|2686,2692|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|2686,2692|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|2701,2709|false|false|false|||pleasant
Finding|Mental Process|SIMPLE_SEGMENT|2701,2709|false|false|false|C2987187|Pleasant|pleasant
Event|Event|SIMPLE_SEGMENT|2714,2721|false|false|false|||tearful
Finding|Finding|SIMPLE_SEGMENT|2714,2721|false|false|false|C0424109|Weepiness|tearful
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2760,2765|false|false|false|C1512338|HEENT|HEENT
Event|Event|SIMPLE_SEGMENT|2781,2788|false|false|false|||lesions
Finding|Finding|SIMPLE_SEGMENT|2781,2788|true|false|false|C0221198|Lesion|lesions
Finding|Intellectual Product|SIMPLE_SEGMENT|2790,2794|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2795,2802|false|false|false|C0036410|Sclera|scleral
Finding|Finding|SIMPLE_SEGMENT|2795,2810|false|false|false|C0240962|Scleral icterus|scleral icterus
Event|Event|SIMPLE_SEGMENT|2803,2810|false|false|false|||icterus
Finding|Sign or Symptom|SIMPLE_SEGMENT|2803,2810|false|false|false|C0022346|Icterus|icterus
Event|Event|SIMPLE_SEGMENT|2831,2834|false|false|false|||MRG
Finding|Gene or Genome|SIMPLE_SEGMENT|2831,2834|true|false|false|C1422304|MAS1L gene|MRG
Event|Event|SIMPLE_SEGMENT|2837,2841|false|false|false|||PULM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2837,2841|false|false|false|C1315068|Pulmonary ventilator management|PULM
Event|Event|SIMPLE_SEGMENT|2853,2861|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2853,2861|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|2862,2863|false|false|false|||R
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2870,2873|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2870,2873|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|SIMPLE_SEGMENT|2870,2873|false|false|false|||ABD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2880,2884|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2886,2895|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|2886,2895|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|2907,2913|false|false|false|||tender
Finding|Intellectual Product|SIMPLE_SEGMENT|2919,2923|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|2924,2931|false|false|false|||rebound
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2942,2952|false|false|false|C1275670|Collateral branch of vessel|collateral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2953,2958|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2953,2958|false|false|false|C0398102|Procedure on vein|veins
Finding|Intellectual Product|SIMPLE_SEGMENT|2965,2969|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|SIMPLE_SEGMENT|2970,2979|false|false|false|||angiomata
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2982,2987|false|false|false|C0015385|Limb structure|LIMBS
Finding|Functional Concept|SIMPLE_SEGMENT|2989,2994|false|false|false|C1883002|Sequence Chromatogram|Trace
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2999,3004|false|false|false|C1717255||edema
Event|Event|SIMPLE_SEGMENT|2999,3004|false|false|false|||edema
Finding|Pathologic Function|SIMPLE_SEGMENT|2999,3004|false|false|false|C0013604|Edema|edema
Event|Event|SIMPLE_SEGMENT|3009,3016|false|false|false|||tremors
Finding|Sign or Symptom|SIMPLE_SEGMENT|3009,3016|true|false|false|C0040822|Tremor|tremors
Event|Event|SIMPLE_SEGMENT|3020,3029|false|false|false|||asterixis
Finding|Sign or Symptom|SIMPLE_SEGMENT|3020,3029|true|false|false|C0232766|Asterixis|asterixis
Anatomy|Body System|SIMPLE_SEGMENT|3032,3036|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3032,3036|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Event|Event|SIMPLE_SEGMENT|3032,3036|false|false|false|||SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3032,3036|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Event|Event|SIMPLE_SEGMENT|3041,3047|false|false|false|||rashes
Finding|Sign or Symptom|SIMPLE_SEGMENT|3041,3047|true|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Anatomy|Body System|SIMPLE_SEGMENT|3051,3055|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3051,3055|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3051,3055|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|SIMPLE_SEGMENT|3051,3055|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|3051,3055|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Finding|SIMPLE_SEGMENT|3051,3065|true|false|false|C0150077;C4048181|Broken skin;Impaired skin integrity|skin breakdown
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3056,3065|true|false|false|C1265875|Disintegration (morphologic abnormality)|breakdown
Event|Event|SIMPLE_SEGMENT|3056,3065|false|false|false|||breakdown
Finding|Organism Function|SIMPLE_SEGMENT|3056,3065|true|false|false|C0699900|Catabolism|breakdown
Event|Event|SIMPLE_SEGMENT|3077,3087|false|false|false|||ecchymoses
Finding|Pathologic Function|SIMPLE_SEGMENT|3077,3087|true|false|false|C0013491|Ecchymosis|ecchymoses
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3092,3100|false|false|false|C0033119|Puncture wound|puncture
Event|Event|SIMPLE_SEGMENT|3092,3100|false|false|false|||puncture
Procedure|Health Care Activity|SIMPLE_SEGMENT|3092,3100|false|false|false|C0034117|Puncture procedure|puncture
Finding|Pathologic Function|SIMPLE_SEGMENT|3132,3146|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|SIMPLE_SEGMENT|3141,3146|false|false|false|||drift
Event|Event|SIMPLE_SEGMENT|3148,3156|false|false|false|||reflexes
Finding|Finding|SIMPLE_SEGMENT|3148,3156|true|false|false|C0034929;C0596002|Observation of reflex;Reflex action|reflexes
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3148,3156|true|false|false|C0034929;C0596002|Observation of reflex;Reflex action|reflexes
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3148,3156|true|false|false|C0436145|Examination of reflexes|reflexes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3182,3187|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3182,3187|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3182,3199|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3188,3199|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|3223,3227|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3223,3227|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3230,3235|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|3230,3235|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|3230,3235|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Anatomy|Cell|SIMPLE_SEGMENT|3241,3244|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3251,3254|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3251,3254|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3251,3254|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3261,3264|false|false|false|C0019046|Hemoglobin|HGB
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3261,3264|false|false|false|C0019046|Hemoglobin|HGB
Event|Event|SIMPLE_SEGMENT|3261,3264|false|false|false|||HGB
Finding|Gene or Genome|SIMPLE_SEGMENT|3261,3264|false|false|false|C1424337|CYGB gene|HGB
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3261,3264|false|false|false|C0019029|Hemoglobin concentration|HGB
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3271,3274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3271,3274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Disorder|Virus|SIMPLE_SEGMENT|3281,3284|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3281,3284|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3281,3284|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3281,3284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3281,3284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3290,3293|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3290,3293|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3290,3293|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3290,3293|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3290,3293|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3290,3293|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3301,3305|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3301,3305|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3320,3323|false|false|false|C0201617|Primed lymphocyte test|PLT
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3338,3341|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|3338,3341|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3338,3341|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3352,3359|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|SIMPLE_SEGMENT|3352,3359|false|false|false|||ALBUMIN
Finding|Gene or Genome|SIMPLE_SEGMENT|3352,3359|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|SIMPLE_SEGMENT|3352,3359|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3352,3359|false|false|false|C0201838|Albumin measurement|ALBUMIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3365,3368|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3365,3368|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|SIMPLE_SEGMENT|3365,3368|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|SIMPLE_SEGMENT|3365,3368|false|false|false|||ALT
Finding|Gene or Genome|SIMPLE_SEGMENT|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|SIMPLE_SEGMENT|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|SIMPLE_SEGMENT|3365,3368|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3365,3368|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3369,3373|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Drug|Enzyme|SIMPLE_SEGMENT|3369,3373|false|false|false|C0376147|SGPT - Glutamate pyruvate transaminase|SGPT
Event|Event|SIMPLE_SEGMENT|3369,3373|false|false|false|||SGPT
Finding|Gene or Genome|SIMPLE_SEGMENT|3369,3373|false|false|false|C1415274|GPT gene|SGPT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3369,3373|false|false|false|C0036828|Serum Alanine Transaminase Test|SGPT
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3378,3381|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3378,3381|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|SIMPLE_SEGMENT|3378,3381|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|SIMPLE_SEGMENT|3378,3381|false|false|false|||AST
Finding|Gene or Genome|SIMPLE_SEGMENT|3378,3381|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3382,3386|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Drug|Enzyme|SIMPLE_SEGMENT|3382,3386|false|false|false|C0242192|SGOT - Glutamate oxaloacetate transaminase|SGOT
Event|Event|SIMPLE_SEGMENT|3382,3386|false|false|false|||SGOT
Finding|Gene or Genome|SIMPLE_SEGMENT|3382,3386|false|false|false|C1415181|GOT1 gene|SGOT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3382,3386|false|false|false|C0201899|Aspartate aminotransferase measurement|SGOT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3393,3396|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|SIMPLE_SEGMENT|3393,3396|false|false|false|C1663627|ALK protein, human|ALK
Event|Event|SIMPLE_SEGMENT|3393,3396|false|false|false|||ALK
Finding|Gene or Genome|SIMPLE_SEGMENT|3393,3396|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|SIMPLE_SEGMENT|3393,3396|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3393,3401|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|SIMPLE_SEGMENT|3393,3401|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3393,3401|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Event|Event|SIMPLE_SEGMENT|3397,3401|false|false|false|||PHOS
Event|Event|SIMPLE_SEGMENT|3412,3416|false|false|false|||BILI
Finding|Body Substance|SIMPLE_SEGMENT|3422,3435|false|false|false|C5441965|Ascitic Fluid|Ascitic Fluid
Drug|Substance|SIMPLE_SEGMENT|3430,3435|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|SIMPLE_SEGMENT|3430,3435|false|false|false|||Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3430,3435|false|false|false|C1546638|Fluid Specimen Code|Fluid
Anatomy|Cell|SIMPLE_SEGMENT|3443,3446|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3451,3454|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3451,3454|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3451,3454|false|false|false|C0014792|Erythrocytes|RBC
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3459,3464|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|POLYS
Finding|Body Substance|SIMPLE_SEGMENT|3469,3475|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|3480,3485|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3488,3491|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|3488,3491|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|3488,3491|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Event|Event|SIMPLE_SEGMENT|3524,3527|false|false|false|||TOT
Finding|Gene or Genome|SIMPLE_SEGMENT|3528,3532|false|false|false|C1420218|SLC6A7 gene|PROT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3540,3543|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Drug|Enzyme|SIMPLE_SEGMENT|3540,3543|false|false|false|C0022917|Lactate Dehydrogenase|LDH
Event|Event|SIMPLE_SEGMENT|3540,3543|false|false|false|||LDH
Finding|Finding|SIMPLE_SEGMENT|3540,3543|false|false|false|C0851148|Lifetime Drinking History|LDH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3540,3543|false|false|false|C0202113|Lactate dehydrogenase measurement|LDH
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3548,3555|false|false|false|C0001924;C5966160|Albumin;Albumins|ALBUMIN
Event|Event|SIMPLE_SEGMENT|3548,3555|false|false|false|||ALBUMIN
Finding|Gene or Genome|SIMPLE_SEGMENT|3548,3555|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Finding|Physiologic Function|SIMPLE_SEGMENT|3548,3555|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|ALBUMIN
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3548,3555|false|false|false|C0201838|Albumin measurement|ALBUMIN
Finding|Body Substance|SIMPLE_SEGMENT|3562,3575|false|false|false|C5441965|Ascitic Fluid|Ascitic Fluid
Drug|Substance|SIMPLE_SEGMENT|3570,3575|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Event|Event|SIMPLE_SEGMENT|3570,3575|false|false|false|||Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|3570,3575|false|false|false|C1546638|Fluid Specimen Code|Fluid
Anatomy|Cell|SIMPLE_SEGMENT|3581,3584|false|false|false|C0023516|Leukocytes|WBC
Finding|Gene or Genome|SIMPLE_SEGMENT|3590,3593|false|false|false|C1428294;C3812663|NACC2 gene;NACC2 wt Allele|RBB
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3599,3604|false|false|false|C0032400;C0071360|5'-Inosinic acid, 2'-deoxy-2'-fluoro-, homopolymer;Poly A|POLYS
Finding|Body Substance|SIMPLE_SEGMENT|3609,3615|false|false|false|C0024202|Lymph|LYMPHS
Drug|Antibiotic|SIMPLE_SEGMENT|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|3620,3625|false|true|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3629,3632|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Event|Event|SIMPLE_SEGMENT|3629,3632|false|false|false|||EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|3629,3632|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3654,3659|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Event|Event|SIMPLE_SEGMENT|3654,3659|false|false|false|||Blood
Finding|Body Substance|SIMPLE_SEGMENT|3654,3659|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Anatomy|Cell|SIMPLE_SEGMENT|3665,3668|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|3674,3677|false|false|false|||HCT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3674,3677|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3674,3677|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Event|Event|SIMPLE_SEGMENT|3685,3694|false|false|false|||RADIOLOGY
Finding|Finding|SIMPLE_SEGMENT|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Idea or Concept|SIMPLE_SEGMENT|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Finding|Intellectual Product|SIMPLE_SEGMENT|3685,3694|false|false|false|C1405978;C1548000;C1548429|Encounter due to radiological examination;Radiology Section ID;radiology referral type|RADIOLOGY
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3685,3694|false|false|false|C0043299;C0807679;C1962945|Diagnostic radiologic examination;Radiographic imaging procedure;Radiology studies|RADIOLOGY
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3696,3708|false|false|false|C5452879|Lumbo-sacral|Lumbo-sacral
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3702,3708|false|false|false|C0036033;C0036037|Bone structure of sacrum;Sacral Region|sacral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3702,3708|false|false|false|C0036033;C0036037|Bone structure of sacrum;Sacral Region|sacral
Event|Event|SIMPLE_SEGMENT|3713,3719|false|false|false|||Normal
Event|Event|SIMPLE_SEGMENT|3724,3732|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|3724,3732|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|3724,3735|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3736,3749|true|false|false|C0029443|Osteomyelitis|osteomyelitis
Event|Event|SIMPLE_SEGMENT|3736,3749|false|false|false|||osteomyelitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3750,3759|false|false|false|C0549207|Bone structure of spine|vertebral
Event|Event|SIMPLE_SEGMENT|3761,3772|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|3761,3772|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3761,3772|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|3761,3772|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3761,3772|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|3761,3781|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3773,3781|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|3773,3781|false|false|false|||fracture
Finding|Intellectual Product|SIMPLE_SEGMENT|3786,3791|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|3792,3800|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3792,3807|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|3792,3807|false|false|false|C0489547|Hospital course|Hospital Course
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3810,3819|false|false|false|C0000726|Abdomen|Abdominal
Finding|Finding|SIMPLE_SEGMENT|3810,3830|false|false|false|C0000731|Abdomen distended|Abdominal distention
Event|Event|SIMPLE_SEGMENT|3820,3830|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|3820,3830|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|3820,3830|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3831,3835|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3831,3835|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3831,3835|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3831,3835|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3845,3852|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|3872,3879|false|false|false|||concern
Finding|Idea or Concept|SIMPLE_SEGMENT|3872,3879|false|false|false|C2699424|Concern|concern
Event|Event|SIMPLE_SEGMENT|3884,3895|false|false|false|||spontaneous
Finding|Functional Concept|SIMPLE_SEGMENT|3884,3895|false|false|false|C0205359|Spontaneous|spontaneous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3897,3918|false|false|false|C0275550;C0341503|Acute bacterial peritonitis;Bacterial peritonitis|bacterial peritonitis
Event|Event|SIMPLE_SEGMENT|3907,3918|false|false|false|||peritonitis
Finding|Pathologic Function|SIMPLE_SEGMENT|3907,3918|false|false|false|C0031154|Peritonitis|peritonitis
Drug|Antibiotic|SIMPLE_SEGMENT|3924,3935|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|SIMPLE_SEGMENT|3924,3935|false|false|false|C0007561|ceftriaxone|ceftriaxone
Event|Event|SIMPLE_SEGMENT|3924,3935|false|false|false|||ceftriaxone
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|3947,3957|false|false|false|C0358514|Diagnostic agents|diagnostic
Event|Event|SIMPLE_SEGMENT|3947,3957|false|false|false|||diagnostic
Finding|Functional Concept|SIMPLE_SEGMENT|3947,3957|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Finding|Intellectual Product|SIMPLE_SEGMENT|3947,3957|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3947,3957|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|diagnostic
Event|Event|SIMPLE_SEGMENT|3959,3971|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3959,3971|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Body Substance|SIMPLE_SEGMENT|3998,4011|false|false|false|C5441965|Ascitic Fluid|Ascitic fluid
Drug|Substance|SIMPLE_SEGMENT|4006,4011|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4006,4011|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|4012,4020|false|false|false|||analysis
Finding|Functional Concept|SIMPLE_SEGMENT|4012,4020|false|false|false|C1524024|analysis aspect|analysis
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4012,4020|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Procedure|Research Activity|SIMPLE_SEGMENT|4012,4020|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Finding|Functional Concept|SIMPLE_SEGMENT|4038,4049|false|false|false|C0205359|Spontaneous|Spontaneous
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4038,4071|false|false|false|C0275551;C2062979|Primary bacterial peritonitis;acute spontaneous bacterial peritonitis|Spontaneous bacterial peritonitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4050,4071|false|false|false|C0275550;C0341503|Acute bacterial peritonitis;Bacterial peritonitis|bacterial peritonitis
Event|Event|SIMPLE_SEGMENT|4060,4071|false|false|false|||peritonitis
Finding|Pathologic Function|SIMPLE_SEGMENT|4060,4071|false|false|false|C0031154|Peritonitis|peritonitis
Event|Event|SIMPLE_SEGMENT|4076,4081|false|false|false|||ruled
Event|Event|SIMPLE_SEGMENT|4087,4092|false|false|false|||given
Drug|Substance|SIMPLE_SEGMENT|4102,4107|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4102,4107|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Cell|SIMPLE_SEGMENT|4108,4112|false|false|false|C0007634|Cells|cell
Finding|Gene or Genome|SIMPLE_SEGMENT|4108,4112|false|false|false|C1413336;C1413337|CEL gene;CELP gene|cell
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4108,4118|false|false|false|C0007584|Cell Count|cell count
Event|Event|SIMPLE_SEGMENT|4113,4118|false|false|false|||count
Event|Event|SIMPLE_SEGMENT|4119,4125|false|false|false|||showed
Anatomy|Cell|SIMPLE_SEGMENT|4134,4137|false|false|false|C0023516|Leukocytes|WBC
Drug|Antibiotic|SIMPLE_SEGMENT|4139,4150|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|SIMPLE_SEGMENT|4139,4150|false|false|false|||antibiotics
Event|Event|SIMPLE_SEGMENT|4157,4169|false|false|false|||discontinued
Finding|Mental Process|SIMPLE_SEGMENT|4178,4185|false|false|false|C0542559|contextual factors|setting
Finding|Gene or Genome|SIMPLE_SEGMENT|4204,4209|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|4210,4216|false|false|false|||volume
Finding|Intellectual Product|SIMPLE_SEGMENT|4210,4216|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|4218,4230|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4218,4230|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Substance|SIMPLE_SEGMENT|4265,4271|false|false|false|C0302908|Liquid substance|fluids
Event|Event|SIMPLE_SEGMENT|4265,4271|false|false|false|||fluids
Finding|Body Substance|SIMPLE_SEGMENT|4265,4271|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4265,4271|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|SIMPLE_SEGMENT|4273,4280|false|false|false|||removed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4292,4301|false|false|false|C0945766||procedure
Event|Event|SIMPLE_SEGMENT|4292,4301|false|false|false|||procedure
Event|Occupational Activity|SIMPLE_SEGMENT|4292,4301|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|SIMPLE_SEGMENT|4292,4301|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4292,4301|false|false|false|C0184661|Interventional procedure|procedure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4307,4314|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4307,4314|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|4307,4314|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|SIMPLE_SEGMENT|4324,4333|false|false|false|||distended
Finding|Finding|SIMPLE_SEGMENT|4324,4333|false|false|false|C0700124|Dilated|distended
Event|Event|SIMPLE_SEGMENT|4344,4351|false|false|false|||painful
Finding|Sign or Symptom|SIMPLE_SEGMENT|4344,4351|false|false|false|C0030193|Pain|painful
Drug|Substance|SIMPLE_SEGMENT|4354,4359|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|4354,4359|false|false|false|C1546638|Fluid Specimen Code|Fluid
Event|Event|SIMPLE_SEGMENT|4360,4368|false|false|false|||analysis
Finding|Functional Concept|SIMPLE_SEGMENT|4360,4368|false|false|false|C1524024|analysis aspect|analysis
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4360,4368|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Procedure|Research Activity|SIMPLE_SEGMENT|4360,4368|false|false|false|C0002778;C0936012|Analysis;Analysis of substances|analysis
Event|Event|SIMPLE_SEGMENT|4383,4389|false|false|false|||reveal
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4390,4393|true|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4390,4393|true|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4390,4393|true|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|SIMPLE_SEGMENT|4390,4393|false|false|false|||SBP
Finding|Gene or Genome|SIMPLE_SEGMENT|4390,4393|true|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4390,4393|true|false|false|C1306620|Systolic blood pressure measurement|SBP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4400,4419|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4410,4419|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|SIMPLE_SEGMENT|4410,4419|false|false|false|||hepatitis
Finding|Body Substance|SIMPLE_SEGMENT|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4421,4428|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|4431,4436|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|4431,4436|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|4431,4436|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|4431,4436|false|false|false|C0872387|Procedures on liver|liver
Event|Activity|SIMPLE_SEGMENT|4437,4446|false|false|false|C1883254|Synthesis|synthetic
Event|Event|SIMPLE_SEGMENT|4447,4455|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|4447,4455|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|4460,4469|false|false|false|||monitored
Event|Event|SIMPLE_SEGMENT|4477,4489|false|false|false|||hospitalized
Event|Event|SIMPLE_SEGMENT|4499,4509|false|false|false|||maintained
Finding|Idea or Concept|SIMPLE_SEGMENT|4517,4521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|4517,4521|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|4517,4521|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|4522,4529|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|4522,4529|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4522,4529|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Organic Chemical|SIMPLE_SEGMENT|4534,4543|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4534,4543|false|false|false|C0022957|lactulose|lactulose
Event|Event|SIMPLE_SEGMENT|4534,4543|false|false|false|||lactulose
Finding|Body Substance|SIMPLE_SEGMENT|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|4564,4569|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4564,4580|false|false|false|C0200354|Urine Specimen Collection|urine collection
Event|Event|SIMPLE_SEGMENT|4570,4580|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|4570,4580|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4585,4591|false|false|false|C0009968|copper|copper
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4585,4591|false|false|false|C0009968|copper|copper
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4585,4591|false|false|false|C0009968|copper|copper
Event|Event|SIMPLE_SEGMENT|4585,4591|false|false|false|||copper
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4585,4591|false|false|false|C0373587|Copper measurement|copper
Event|Event|SIMPLE_SEGMENT|4596,4604|false|false|false|||evaluate
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4613,4620|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|4613,4620|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4626,4638|false|false|false|C0023518|Leukocytosis|Leukocytosis
Event|Event|SIMPLE_SEGMENT|4626,4638|false|false|false|||Leukocytosis
Finding|Finding|SIMPLE_SEGMENT|4626,4638|false|false|false|C0750426|Blood leukocyte number above reference range|Leukocytosis
Finding|Intellectual Product|SIMPLE_SEGMENT|4643,4647|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|4643,4653|false|false|false|C0239574|Low grade fever|mild fever
Event|Event|SIMPLE_SEGMENT|4648,4653|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|4648,4653|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|4648,4653|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|4665,4676|false|false|false|||temparature
Event|Event|SIMPLE_SEGMENT|4689,4701|false|false|false|||presentation
Finding|Idea or Concept|SIMPLE_SEGMENT|4689,4701|false|false|false|C0449450|Presentation|presentation
Event|Event|SIMPLE_SEGMENT|4726,4731|false|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|4726,4731|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|4726,4731|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|4735,4743|false|false|false|||symptoms
Finding|Functional Concept|SIMPLE_SEGMENT|4735,4743|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|4735,4743|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4751,4760|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|4751,4760|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|4751,4760|true|false|false|C3714514|Infection|infection
Finding|Body Substance|SIMPLE_SEGMENT|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Functional Concept|SIMPLE_SEGMENT|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Finding|Intellectual Product|SIMPLE_SEGMENT|4763,4768|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|Urine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4763,4776|false|false|false|C0430404|Urine culture|Urine culture
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4769,4776|false|false|false|C1706355|Culture Dose Form|culture
Event|Event|SIMPLE_SEGMENT|4769,4776|false|false|false|||culture
Finding|Functional Concept|SIMPLE_SEGMENT|4769,4776|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|SIMPLE_SEGMENT|4769,4776|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4769,4776|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Event|Event|SIMPLE_SEGMENT|4777,4783|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|4800,4810|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4800,4810|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|4800,4815|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|4816,4829|false|false|false|||contamination
Finding|Idea or Concept|SIMPLE_SEGMENT|4816,4829|false|false|false|C2349974|Contamination|contamination
Phenomenon|Human-caused Phenomenon or Process|SIMPLE_SEGMENT|4816,4829|false|false|false|C0259846|adulteration|contamination
Event|Activity|SIMPLE_SEGMENT|4837,4844|false|false|false|C1706079||arrival
Event|Event|SIMPLE_SEGMENT|4837,4844|false|false|false|||arrival
Finding|Functional Concept|SIMPLE_SEGMENT|4837,4844|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|4853,4858|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|SIMPLE_SEGMENT|4863,4874|false|false|false|||temperature
Procedure|Health Care Activity|SIMPLE_SEGMENT|4863,4874|false|false|false|C0886414|Body temperature measurement|temperature
Event|Event|SIMPLE_SEGMENT|4879,4885|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|4879,4885|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|4887,4894|false|false|false|||ranging
Anatomy|Cell|SIMPLE_SEGMENT|4917,4920|false|false|false|C0023516|Leukocytes|WBC
Event|Event|SIMPLE_SEGMENT|4921,4928|false|false|false|||trended
Event|Event|SIMPLE_SEGMENT|4949,4964|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|4949,4964|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Finding|SIMPLE_SEGMENT|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|4984,4988|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|4992,5001|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4992,5001|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4992,5001|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|5010,5021|false|false|false|||Tachycardia
Finding|Finding|SIMPLE_SEGMENT|5010,5021|false|false|false|C0039231;C3827868|Tachycardia;Tachycardia by ECG Finding|Tachycardia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5027,5032|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5027,5032|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|5027,5032|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5027,5037|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|5027,5037|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|5027,5037|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|5033,5037|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|5033,5037|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|5033,5037|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|5042,5050|false|false|false|||elevated
Event|Event|SIMPLE_SEGMENT|5062,5066|false|false|false|||120s
Event|Event|SIMPLE_SEGMENT|5083,5098|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|5083,5098|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Idea or Concept|SIMPLE_SEGMENT|5108,5112|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|SIMPLE_SEGMENT|5113,5124|false|false|false|||oxygenation
Finding|Cell Function|SIMPLE_SEGMENT|5113,5124|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|5113,5124|false|false|false|C0231940;C0282636|Alveolar ventilation function;Cell Respiration|oxygenation
Event|Event|SIMPLE_SEGMENT|5136,5146|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|5136,5146|true|false|false|C5441521|Complaint (finding)|complaints
Event|Event|SIMPLE_SEGMENT|5151,5154|false|false|false|||SOB
Finding|Sign or Symptom|SIMPLE_SEGMENT|5151,5154|false|false|false|C0013404|Dyspnea|SOB
Event|Event|SIMPLE_SEGMENT|5156,5163|false|false|false|||dyspnea
Finding|Finding|SIMPLE_SEGMENT|5156,5163|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|5156,5163|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5165,5170|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|5165,5170|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5165,5175|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5165,5175|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5171,5175|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5171,5175|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5171,5175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5171,5175|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5177,5189|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|5177,5189|false|false|false|C0030252|Palpitations|palpitations
Finding|Idea or Concept|SIMPLE_SEGMENT|5195,5206|false|false|false|C0750501|most likely|most likely
Finding|Finding|SIMPLE_SEGMENT|5200,5206|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5200,5206|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|SIMPLE_SEGMENT|5208,5216|false|false|false|||etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|5208,5216|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|SIMPLE_SEGMENT|5208,5216|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5228,5232|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5228,5232|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5228,5232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5228,5232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5234,5241|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|SIMPLE_SEGMENT|5234,5241|false|false|false|||anxiety
Finding|Sign or Symptom|SIMPLE_SEGMENT|5234,5241|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Finding|SIMPLE_SEGMENT|5251,5254|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|SIMPLE_SEGMENT|5251,5254|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|SIMPLE_SEGMENT|5255,5268|false|false|false|||intravascular
Finding|Functional Concept|SIMPLE_SEGMENT|5255,5268|false|false|false|C2960476|Intravascular Route of Administration|intravascular
Event|Event|SIMPLE_SEGMENT|5270,5276|false|false|false|||volume
Finding|Intellectual Product|SIMPLE_SEGMENT|5270,5276|false|false|false|C1705102|Volume (publication)|volume
Event|Event|SIMPLE_SEGMENT|5287,5298|false|false|false|||tachycardic
Event|Event|SIMPLE_SEGMENT|5316,5325|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5316,5325|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5316,5325|false|false|false|C0030685|Patient Discharge|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5332,5341|false|false|false|C0004604|Back Pain|Back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5337,5341|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5337,5341|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5337,5341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5337,5341|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5343,5360|false|false|false|C0223603|Lumbosacral spine|Lumbosacral spine
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5355,5360|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|SIMPLE_SEGMENT|5355,5360|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|SIMPLE_SEGMENT|5355,5360|false|false|false|C0150920|Spine Problem|spine
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5361,5365|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Drug|Substance|SIMPLE_SEGMENT|5361,5365|false|false|false|C1561572;C1704608|Film Dosage Form;film - layer|film
Event|Event|SIMPLE_SEGMENT|5361,5365|false|false|false|||film
Finding|Intellectual Product|SIMPLE_SEGMENT|5361,5365|false|false|false|C4019020||film
Event|Event|SIMPLE_SEGMENT|5366,5374|false|false|false|||revealed
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5378,5400|true|false|false|C4021790|Abnormality of the skeletal system|skeletal abnormalities
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|5387,5400|true|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|SIMPLE_SEGMENT|5387,5400|false|false|false|||abnormalities
Finding|Functional Concept|SIMPLE_SEGMENT|5387,5400|true|false|false|C0000769|teratologic|abnormalities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5403,5412|false|false|false|C0549207|Bone structure of spine|vertebral
Finding|Pathologic Function|SIMPLE_SEGMENT|5403,5424|false|false|false|C0262431|Compression fracture of vertebral column|vertebral compression
Finding|Pathologic Function|SIMPLE_SEGMENT|5403,5433|false|false|false|C0262431|Compression fracture of vertebral column|vertebral compression fracture
Event|Event|SIMPLE_SEGMENT|5413,5424|false|false|false|||compression
Finding|Functional Concept|SIMPLE_SEGMENT|5413,5424|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5413,5424|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|SIMPLE_SEGMENT|5413,5424|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5413,5424|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Finding|Pathologic Function|SIMPLE_SEGMENT|5413,5433|false|false|false|C0521169|Compression fracture|compression fracture
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5425,5433|false|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|5425,5433|false|false|false|||fracture
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5438,5451|false|false|false|C0029443|Osteomyelitis|osteomyelitis
Event|Event|SIMPLE_SEGMENT|5438,5451|false|false|false|||osteomyelitis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5459,5463|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5459,5463|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5459,5463|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5459,5463|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5469,5476|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|5469,5476|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|5469,5476|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Finding|SIMPLE_SEGMENT|5481,5485|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|5486,5496|false|false|false|||controlled
Event|Event|SIMPLE_SEGMENT|5512,5527|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|5512,5527|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Organic Chemical|SIMPLE_SEGMENT|5534,5543|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5534,5543|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|SIMPLE_SEGMENT|5534,5543|false|false|false|||oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5534,5543|false|false|false|C0524222|Oxycodone measurement|oxycodone
Finding|Gene or Genome|SIMPLE_SEGMENT|5552,5555|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5556,5560|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5556,5560|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5556,5560|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5556,5560|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|5563,5574|false|false|false|||Recommended
Event|Event|SIMPLE_SEGMENT|5575,5581|false|false|false|||follow
Finding|Intellectual Product|SIMPLE_SEGMENT|5595,5607|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|5595,5607|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5595,5616|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|SIMPLE_SEGMENT|5595,5616|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|SIMPLE_SEGMENT|5603,5607|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|5603,5607|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|5603,5607|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|5603,5607|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|SIMPLE_SEGMENT|5608,5616|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|SIMPLE_SEGMENT|5608,5616|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Event|SIMPLE_SEGMENT|5620,5627|false|false|false|||address
Event|Event|SIMPLE_SEGMENT|5628,5638|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|5628,5638|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|5628,5638|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|5646,5653|false|false|false|||chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|5646,5653|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|5646,5653|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5655,5659|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5655,5659|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5655,5659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5655,5659|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Food|SIMPLE_SEGMENT|5665,5669|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|Diet
Event|Event|SIMPLE_SEGMENT|5665,5669|false|false|false|||Diet
Finding|Functional Concept|SIMPLE_SEGMENT|5665,5669|false|false|false|C1549512|diet - supply|Diet
Procedure|Health Care Activity|SIMPLE_SEGMENT|5665,5669|false|false|false|C0012159|Diet therapy|Diet
Finding|Finding|SIMPLE_SEGMENT|5671,5674|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Intellectual Product|SIMPLE_SEGMENT|5671,5674|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|Low
Finding|Finding|SIMPLE_SEGMENT|5671,5681|false|false|false|C0860871|Sodium decreased|Low sodium
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5671,5681|false|false|false|C0012169|Low sodium diet|Low sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5675,5681|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|SIMPLE_SEGMENT|5675,5681|false|false|false|||sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|5675,5681|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5675,5681|false|false|false|C0337443|Sodium measurement|sodium
Finding|Idea or Concept|SIMPLE_SEGMENT|5686,5689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5686,5689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Substance|SIMPLE_SEGMENT|5692,5697|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|5692,5697|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5692,5709|false|false|false|C0204700|Fluid restriction|fluid restriction
Event|Event|SIMPLE_SEGMENT|5698,5709|false|false|false|||restriction
Finding|Functional Concept|SIMPLE_SEGMENT|5698,5709|false|false|false|C0443288|Restricted|restriction
Finding|Idea or Concept|SIMPLE_SEGMENT|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|SIMPLE_SEGMENT|5718,5721|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|SIMPLE_SEGMENT|5726,5730|false|false|false|||Code
Event|Occupational Activity|SIMPLE_SEGMENT|5726,5730|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|SIMPLE_SEGMENT|5726,5730|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5740,5751|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5740,5751|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5740,5751|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5740,5751|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|5740,5764|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|5755,5764|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5755,5764|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Organic Chemical|SIMPLE_SEGMENT|5768,5781|false|false|false|C0002600|amitriptyline|AMITRIPTYLINE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5768,5781|false|false|false|C0002600|amitriptyline|AMITRIPTYLINE
Drug|Organic Chemical|SIMPLE_SEGMENT|5800,5809|false|false|false|C0030049|oxycodone|OXYCODONE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5800,5809|false|false|false|C0030049|oxycodone|OXYCODONE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5800,5809|false|false|false|C0524222|Oxycodone measurement|OXYCODONE
Finding|Gene or Genome|SIMPLE_SEGMENT|5824,5827|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5828,5832|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|5828,5832|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|5828,5832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|5828,5832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|SIMPLE_SEGMENT|5837,5845|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Event|Event|SIMPLE_SEGMENT|5837,5845|false|false|false|||Thiamine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5837,5845|false|false|false|C0373727|Thiamine measurement|Thiamine
Event|Event|SIMPLE_SEGMENT|5852,5854|false|false|false|||PO
Drug|Organic Chemical|SIMPLE_SEGMENT|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Drug|Vitamin|SIMPLE_SEGMENT|5865,5875|false|false|false|C0016410|folic acid|Folic acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5865,5875|false|false|false|C0523631|Folic acid measurement|Folic acid
Event|Event|SIMPLE_SEGMENT|5871,5875|false|false|false|||acid
Event|Event|SIMPLE_SEGMENT|5893,5896|false|false|false|||MVI
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5893,5896|false|false|false|C5417720|MVI Regimen|MVI
Event|Event|SIMPLE_SEGMENT|5910,5919|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|5910,5919|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|5910,5919|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|5910,5931|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5920,5931|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5920,5931|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|5920,5931|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5920,5931|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Drug|Vitamin|SIMPLE_SEGMENT|5936,5944|false|false|false|C0039840;C3714802|Thiamine Drug Class;thiamine|Thiamine
Event|Event|SIMPLE_SEGMENT|5936,5944|false|false|false|||Thiamine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5936,5944|false|false|false|C0373727|Thiamine measurement|Thiamine
Drug|Organic Chemical|SIMPLE_SEGMENT|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Drug|Vitamin|SIMPLE_SEGMENT|5936,5948|false|false|false|C0770309|thiamine hydrochloride|Thiamine HCl
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5945,5948|false|false|false|C0023443|Hairy Cell Leukemia|HCl
Drug|Immunologic Factor|SIMPLE_SEGMENT|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5945,5948|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|HCl
Event|Event|SIMPLE_SEGMENT|5945,5948|false|false|false|||HCl
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5956,5962|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5976,5982|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|5976,5982|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Drug|Vitamin|SIMPLE_SEGMENT|6005,6015|false|false|false|C0016410|folic acid|Folic Acid
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6005,6015|false|false|false|C0523631|Folic acid measurement|Folic Acid
Event|Event|SIMPLE_SEGMENT|6011,6015|false|false|false|||Acid
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6021,6027|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6028,6031|false|false|false|||Sig
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6041,6047|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6041,6047|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|6072,6085|false|false|false|C0002600|amitriptyline|Amitriptyline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6072,6085|false|false|false|C0002600|amitriptyline|Amitriptyline
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6092,6098|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6092,6098|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6112,6118|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6112,6118|false|false|false|||Tablet
Event|Event|SIMPLE_SEGMENT|6130,6137|false|false|false|||bedtime
Drug|Organic Chemical|SIMPLE_SEGMENT|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Vitamin|SIMPLE_SEGMENT|6145,6157|false|false|false|C0301532|Multivitamin preparation|Multivitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6145,6168|false|false|false|C0978787|Multivitamin tablet|Multivitamin     Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6162,6168|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6162,6168|false|false|false|||Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6182,6188|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6182,6188|false|false|false|||Tablet
Drug|Organic Chemical|SIMPLE_SEGMENT|6213,6222|true|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6213,6222|true|false|false|C0022957|lactulose|Lactulose
Event|Event|SIMPLE_SEGMENT|6213,6222|false|false|false|||Lactulose
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6237,6242|true|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|Syrup
Drug|Food|SIMPLE_SEGMENT|6237,6242|true|false|false|C0458173;C0991550|Syrup (dietary);Syrup Drug Form|Syrup
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6243,6246|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|SIMPLE_SEGMENT|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|SIMPLE_SEGMENT|6243,6246|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Organic Chemical|SIMPLE_SEGMENT|6287,6296|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6287,6296|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|SIMPLE_SEGMENT|6287,6296|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6287,6296|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6302,6308|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6322,6328|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|SIMPLE_SEGMENT|6358,6364|false|false|false|||needed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6369,6373|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6369,6373|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6369,6373|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6369,6373|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6380,6389|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6380,6389|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6380,6389|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6380,6401|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6380,6401|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6390,6401|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|6390,6401|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6390,6401|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|SIMPLE_SEGMENT|6403,6407|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|6403,6407|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6403,6407|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6403,6407|false|false|false|C1553498|home health encounter|Home
Event|Event|SIMPLE_SEGMENT|6410,6419|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6410,6419|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6410,6419|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6410,6429|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6420,6429|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|6420,6429|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6420,6429|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6420,6429|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6420,6429|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6440,6447|false|false|false|C0003962|Ascites|Ascites
Event|Event|SIMPLE_SEGMENT|6440,6447|false|false|false|||Ascites
Finding|Pathologic Function|SIMPLE_SEGMENT|6440,6447|false|false|false|C5441966|Peritoneal Effusion|Ascites
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6448,6454|false|false|false|C0205054|Hepatic|Portal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6448,6467|false|false|false|C0020541|Portal Hypertension|Portal hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6455,6467|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|6455,6467|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6468,6487|false|false|false|C0019187|Hepatitis, Alcoholic|Alcoholic hepatitis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6478,6487|false|false|false|C0019158;C0019159|Hepatitis;Hepatitis A|hepatitis
Event|Event|SIMPLE_SEGMENT|6478,6487|false|false|false|||hepatitis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6490,6499|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|6490,6499|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|6490,6499|false|false|false|C1522484|metastatic qualifier|Secondary
Event|Event|SIMPLE_SEGMENT|6501,6508|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|6501,6508|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|6501,6508|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Finding|Sign or Symptom|SIMPLE_SEGMENT|6501,6518|false|true|false|C0740418|Chronic back pain|Chronic back pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6509,6518|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6514,6518|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6514,6518|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6514,6518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6514,6518|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6522,6531|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6522,6531|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6522,6531|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6522,6531|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6522,6531|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6532,6541|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6532,6541|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|6532,6541|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|6532,6541|false|false|false|C1705253|Logical Condition|Condition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6543,6548|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|6543,6548|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6543,6548|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|6543,6548|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|6543,6548|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|6553,6561|false|false|false|||Oriented
Finding|Finding|SIMPLE_SEGMENT|6553,6561|false|false|false|C1961028|Oriented to place|Oriented
Event|Event|SIMPLE_SEGMENT|6564,6574|false|false|false|||Ambulating
Finding|Intellectual Product|SIMPLE_SEGMENT|6575,6587|false|false|false|C3827452|Without Help|without help
Event|Event|SIMPLE_SEGMENT|6583,6587|false|false|false|||help
Finding|Intellectual Product|SIMPLE_SEGMENT|6583,6587|true|false|false|C1552861|Help document|help
Event|Event|SIMPLE_SEGMENT|6607,6613|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6607,6613|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|6615,6623|false|false|false|||afebrile
Finding|Finding|SIMPLE_SEGMENT|6615,6623|false|false|false|C0277797|Apyrexial|afebrile
Event|Event|SIMPLE_SEGMENT|6625,6636|false|false|false|||tachycardic
Event|Event|SIMPLE_SEGMENT|6643,6652|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|6643,6652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6643,6652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6643,6652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6643,6652|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6643,6665|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6643,6665|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|6643,6665|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6653,6665|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|6653,6665|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|6653,6665|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Event|Event|SIMPLE_SEGMENT|6676,6680|false|false|false|||seen
Event|Event|SIMPLE_SEGMENT|6709,6719|false|false|false|||complaints
Finding|Finding|SIMPLE_SEGMENT|6709,6719|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Functional Concept|SIMPLE_SEGMENT|6723,6733|false|false|false|C0442808|Increasing (qualifier value)|increasing
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6734,6743|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|SIMPLE_SEGMENT|6734,6754|false|false|false|C0000731|Abdomen distended|abdominal distention
Finding|Finding|SIMPLE_SEGMENT|6734,6763|false|false|false|C2749840|Abdominal distention and pain|abdominal distention and pain
Event|Event|SIMPLE_SEGMENT|6744,6754|false|false|false|||distention
Finding|Finding|SIMPLE_SEGMENT|6744,6754|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Finding|Pathologic Function|SIMPLE_SEGMENT|6744,6754|false|false|false|C0012359;C3714614|Distention;Pathological Dilatation|distention
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6759,6763|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6759,6763|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6759,6763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6759,6763|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|SIMPLE_SEGMENT|6796,6800|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Finding|SIMPLE_SEGMENT|6796,6806|false|false|false|C0239574|Low grade fever|mild fever
Event|Event|SIMPLE_SEGMENT|6801,6806|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|6801,6806|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|6801,6806|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Finding|SIMPLE_SEGMENT|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Gene or Genome|SIMPLE_SEGMENT|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Molecular Function|SIMPLE_SEGMENT|6808,6812|false|false|false|C0015663;C1366532;C1705510;C2266413;C3889229|FASTK Gene;FASTK wt Allele;FOXD3-AS1 gene;Fas-activated serine/threonine kinase activity;Fasting|fast
Finding|Finding|SIMPLE_SEGMENT|6808,6823|false|false|false|C0039231|Tachycardia|fast heart rate
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6813,6818|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|6813,6818|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|6813,6818|false|false|false|C0795691|HEART PROBLEM|heart
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6813,6823|false|false|false|C0018810;C0488794|heart rate|heart rate
Finding|Finding|SIMPLE_SEGMENT|6813,6823|false|false|false|C2041121||heart rate
Procedure|Health Care Activity|SIMPLE_SEGMENT|6813,6823|false|false|false|C2197023|examination of heart rate|heart rate
Event|Activity|SIMPLE_SEGMENT|6819,6823|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|6819,6823|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|6819,6823|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|6830,6839|false|false|false|||increased
Finding|Finding|SIMPLE_SEGMENT|6840,6857|false|false|false|C1821144|White blood count|white blood count
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6846,6851|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6846,6851|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6846,6851|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6846,6857|false|false|false|C0005771|Blood Cell Count|blood count
Event|Event|SIMPLE_SEGMENT|6852,6857|false|false|false|||count
Event|Event|SIMPLE_SEGMENT|6869,6873|false|false|false|||sent
Event|Event|SIMPLE_SEGMENT|6881,6890|false|false|false|||emergency
Finding|Finding|SIMPLE_SEGMENT|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|SIMPLE_SEGMENT|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|SIMPLE_SEGMENT|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|SIMPLE_SEGMENT|6881,6890|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|6881,6890|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|SIMPLE_SEGMENT|6881,6890|false|false|false|C1553500|emergency encounter|emergency
Event|Event|SIMPLE_SEGMENT|6892,6902|false|false|false|||department
Finding|Idea or Concept|SIMPLE_SEGMENT|6892,6902|false|false|false|C1547537;C1548283;C1549615|Department - Charge type;Department - No suggested values defined;Organization Unit Type - Department|department
Event|Event|SIMPLE_SEGMENT|6907,6915|false|false|false|||admitted
Finding|Idea or Concept|SIMPLE_SEGMENT|6923,6931|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|6944,6950|false|false|false|||workup
Event|Event|SIMPLE_SEGMENT|6965,6980|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|6965,6980|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Body Substance|SIMPLE_SEGMENT|6986,6999|false|false|false|C5441965|Ascitic Fluid|ascitic fluid
Drug|Substance|SIMPLE_SEGMENT|6994,6999|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|6994,6999|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|6994,6999|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7004,7010|false|false|false|||tapped
Event|Event|SIMPLE_SEGMENT|7016,7024|false|false|false|||analyzed
Event|Event|SIMPLE_SEGMENT|7031,7037|false|false|false|||result
Finding|Finding|SIMPLE_SEGMENT|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|7031,7037|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Event|Event|SIMPLE_SEGMENT|7038,7044|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|7062,7066|false|false|false|||have
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7070,7079|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|7070,7079|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|7070,7079|true|false|false|C3714514|Infection|infection
Finding|Body Substance|SIMPLE_SEGMENT|7088,7101|false|false|false|C5441965|Ascitic Fluid|ascitic fluid
Drug|Substance|SIMPLE_SEGMENT|7096,7101|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7096,7101|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7096,7101|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Substance|SIMPLE_SEGMENT|7118,7123|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|SIMPLE_SEGMENT|7118,7123|false|false|false|||fluid
Finding|Intellectual Product|SIMPLE_SEGMENT|7118,7123|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|SIMPLE_SEGMENT|7128,7135|false|false|false|||removed
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7147,7154|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7147,7154|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Event|Event|SIMPLE_SEGMENT|7147,7154|false|false|false|||abdomen
Finding|Finding|SIMPLE_SEGMENT|7147,7154|false|false|false|C0941288|Abdomen problem|abdomen
Event|Event|SIMPLE_SEGMENT|7159,7171|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7159,7171|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|SIMPLE_SEGMENT|7181,7188|false|false|false|||started
Event|Event|SIMPLE_SEGMENT|7197,7202|false|false|false|||urine
Finding|Body Substance|SIMPLE_SEGMENT|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|SIMPLE_SEGMENT|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|SIMPLE_SEGMENT|7197,7202|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Event|Event|SIMPLE_SEGMENT|7204,7214|false|false|false|||collection
Finding|Conceptual Entity|SIMPLE_SEGMENT|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|SIMPLE_SEGMENT|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|SIMPLE_SEGMENT|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|SIMPLE_SEGMENT|7204,7214|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7219,7225|false|false|false|C0009968|copper|copper
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|7219,7225|false|false|false|C0009968|copper|copper
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7219,7225|false|false|false|C0009968|copper|copper
Event|Event|SIMPLE_SEGMENT|7219,7225|false|false|false|||copper
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7219,7225|false|false|false|C0373587|Copper measurement|copper
Event|Event|SIMPLE_SEGMENT|7229,7233|false|false|false|||work
Event|Event|SIMPLE_SEGMENT|7257,7263|false|false|false|||causes
Finding|Functional Concept|SIMPLE_SEGMENT|7257,7263|false|false|false|C0015127;C1314792|Etiology;Etiology aspects|causes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|7273,7278|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|7273,7278|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|7273,7278|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|7273,7278|false|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7273,7286|false|false|false|C0023895;C0267792|Hepatobiliary Disorder;Liver diseases|liver disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7279,7286|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|7279,7286|false|false|false|||disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|7293,7298|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|7293,7298|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|7293,7298|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|7293,7298|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|7311,7317|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|7345,7352|false|false|false|||results
Event|Event|SIMPLE_SEGMENT|7362,7367|false|false|false|||tests
Finding|Intellectual Product|SIMPLE_SEGMENT|7362,7367|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7362,7367|false|false|false|C0022885|Laboratory Procedures|tests
Finding|Sign or Symptom|SIMPLE_SEGMENT|7378,7387|false|false|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7383,7387|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7383,7387|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7383,7387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7383,7387|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7388,7397|false|false|false|||persisted
Event|Event|SIMPLE_SEGMENT|7410,7425|false|false|false|||hospitalization
Procedure|Health Care Activity|SIMPLE_SEGMENT|7410,7425|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7443,7449|false|false|false|C0885876|X-rays, Homeopathic Preparations|x-rays
Event|Event|SIMPLE_SEGMENT|7443,7449|false|false|false|||x-rays
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7443,7449|false|false|false|C0043309|Roentgen Rays|x-rays
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7443,7449|false|false|false|C0043299;C1306645|Diagnostic radiologic examination;Plain x-ray|x-rays
Event|Event|SIMPLE_SEGMENT|7456,7462|false|false|false|||showed
Event|Event|SIMPLE_SEGMENT|7466,7474|false|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|7466,7474|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|7466,7477|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|7478,7486|true|false|false|C0016658|Fracture|fracture
Event|Event|SIMPLE_SEGMENT|7478,7486|false|false|false|||fracture
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7490,7494|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|SIMPLE_SEGMENT|7490,7494|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|SIMPLE_SEGMENT|7490,7494|true|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7496,7505|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|SIMPLE_SEGMENT|7496,7505|false|false|false|||infection
Finding|Pathologic Function|SIMPLE_SEGMENT|7496,7505|false|false|false|C3714514|Infection|infection
Event|Event|SIMPLE_SEGMENT|7515,7523|false|false|false|||continue
Finding|Idea or Concept|SIMPLE_SEGMENT|7529,7533|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7529,7533|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7529,7533|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7534,7538|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7534,7538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7534,7538|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7539,7546|false|false|false|||regimen
Finding|Intellectual Product|SIMPLE_SEGMENT|7539,7546|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7539,7546|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|SIMPLE_SEGMENT|7551,7560|false|false|false|||readdress
Finding|Intellectual Product|SIMPLE_SEGMENT|7572,7584|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|7572,7584|false|false|false|C0033137|Primary Health Care|primary care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7572,7593|false|false|false|C2735025||primary care provider
Finding|Idea or Concept|SIMPLE_SEGMENT|7572,7593|false|false|false|C1547431|Primary Care Provider - Provider role|primary care provider
Event|Activity|SIMPLE_SEGMENT|7580,7584|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|7580,7584|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|7580,7584|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7580,7584|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Functional Concept|SIMPLE_SEGMENT|7585,7593|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Finding|Intellectual Product|SIMPLE_SEGMENT|7585,7593|false|false|false|C1138603;C1555587|Provider;Transaction counts and value totals - provider|provider
Event|Event|SIMPLE_SEGMENT|7600,7607|false|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|7600,7607|false|false|false|C0392747|Changing|changes
Event|Event|SIMPLE_SEGMENT|7613,7617|false|false|false|||made
Finding|Idea or Concept|SIMPLE_SEGMENT|7626,7630|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|7626,7630|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|7626,7630|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7631,7642|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7631,7642|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7631,7642|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7631,7642|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7657,7665|false|false|false|||continue
Event|Event|SIMPLE_SEGMENT|7669,7672|false|false|false|||use
Drug|Organic Chemical|SIMPLE_SEGMENT|7673,7682|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7673,7682|false|false|false|C0022957|lactulose|lactulose
Event|Event|SIMPLE_SEGMENT|7673,7682|false|false|false|||lactulose
Event|Event|SIMPLE_SEGMENT|7687,7699|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|7687,7699|false|false|false|C0009806|Constipation|constipation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7712,7716|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7712,7716|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7712,7716|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7712,7716|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7718,7729|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7718,7729|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7718,7729|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7718,7729|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7742,7746|false|false|false|||stop
Finding|Intellectual Product|SIMPLE_SEGMENT|7757,7763|false|false|false|C0376667|Herbals (publications)|herbal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7767,7772|false|false|false|C3543842|TONICS|tonic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7773,7781|false|false|false|C0920324|Homeopathic Remedies|remedies
Event|Event|SIMPLE_SEGMENT|7773,7781|false|false|false|||remedies
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|SIMPLE_SEGMENT|7793,7798|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|SIMPLE_SEGMENT|7793,7798|false|false|false|||liver
Finding|Finding|SIMPLE_SEGMENT|7793,7798|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|SIMPLE_SEGMENT|7793,7798|false|false|false|C0872387|Procedures on liver|liver
Event|Event|SIMPLE_SEGMENT|7800,7808|false|false|false|||function
Finding|Finding|SIMPLE_SEGMENT|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|SIMPLE_SEGMENT|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|SIMPLE_SEGMENT|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|SIMPLE_SEGMENT|7800,7808|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Event|Event|SIMPLE_SEGMENT|7813,7822|false|false|false|||recovered
Event|Event|SIMPLE_SEGMENT|7838,7847|false|false|false|||therapies
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7838,7847|false|false|false|C0087111|Therapeutic procedure|therapies
Event|Event|SIMPLE_SEGMENT|7852,7860|false|false|false|||interact
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7872,7879|false|false|false|C1705970|Electrical Current|current
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7880,7891|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7880,7891|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|7880,7891|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|7880,7891|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|7895,7899|false|false|false|||make
Event|Event|SIMPLE_SEGMENT|7903,7912|false|false|false|||difficult
Finding|Finding|SIMPLE_SEGMENT|7903,7912|false|false|false|C0332218|Difficult (qualifier value)|difficult
Event|Event|SIMPLE_SEGMENT|7916,7925|false|false|false|||interpret
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7932,7942|false|false|false|C2598148||laboratory
Finding|Functional Concept|SIMPLE_SEGMENT|7932,7942|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Finding|Intellectual Product|SIMPLE_SEGMENT|7932,7942|false|false|false|C1548427;C1571737;C3244292|Diagnostic Service Section ID - Laboratory;Laboratory domain;Referral type - Laboratory|laboratory
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7932,7942|false|false|false|C4283904|Laboratory observation|laboratory
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|7932,7950|false|false|false|C1254595|Laboratory Results|laboratory results
Event|Event|SIMPLE_SEGMENT|7943,7950|false|false|false|||results
Procedure|Health Care Activity|SIMPLE_SEGMENT|7954,7962|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7963,7975|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|7963,7975|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7963,7975|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

