CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Orthopedics|Title|false|false||ORTHOPAEDICSnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Structure of left knee region|Anatomy|false|false|C1549543;C0030193;C0409959;C1552822;C0029408;C0562271|left knee
null|Structure of left knee|Anatomy|false|false|C1549543;C0030193;C0409959;C1552822;C0029408;C0562271|left kneenull|Table Cell Horizontal Align - left|Finding|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Osteoarthritis, Knee|Disorder|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|knee osteoarthritisnull|Examination of knee joint|Procedure|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C0409959;C0029408;C1552822;C0562271;C1549543;C0030193|knee
null|Knee|Anatomy|false|false|C0409959;C0029408;C1552822;C0562271;C1549543;C0030193|knee
null|Lower extremity>Knee|Anatomy|false|false|C0409959;C0029408;C1552822;C0562271;C1549543;C0030193|knee
null|Knee joint|Anatomy|false|false|C0409959;C0029408;C1552822;C0562271;C1549543;C0030193|kneenull|Degenerative polyarthritis|Disorder|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|osteoarthritisnull|Administration Method - Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|pain
null|Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|painnull|null|Attribute|false|false||painnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Arthroplasty, knee, condyle and plateau; medial AND lateral compartments with or without patella resurfacing (total knee arthroplasty)|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|total knee arthroplasty
null|Knee Replacement Arthroplasty|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|total knee arthroplastynull|Total|Modifier|false|false||totalnull|Knee Replacement Arthroplasty|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|knee arthroplastynull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C0086511;C0371178;C5887062;C0003893;C0700235;C0562271;C0086511|knee
null|Knee|Anatomy|false|false|C0086511;C0371178;C5887062;C0003893;C0700235;C0562271;C0086511|knee
null|Lower extremity>Knee|Anatomy|false|false|C0086511;C0371178;C5887062;C0003893;C0700235;C0562271;C0086511|knee
null|Knee joint|Anatomy|false|false|C0086511;C0371178;C5887062;C0003893;C0700235;C0562271;C0086511|kneenull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|arthroplasty
null|Arthroplasty|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|arthroplasty
null|Reconstruction of joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|arthroplastynull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Old|Time|false|false||oldnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|Structure of left knee region|Anatomy|false|false|C1549543;C0030193;C0562271;C0409959;C0029408|left knee
null|Structure of left knee|Anatomy|false|false|C1549543;C0030193;C0562271;C0409959;C0029408|left kneenull|Table Cell Horizontal Align - left|Finding|false|false|C1963703;C0022742;C4299094;C0022745|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Osteoarthritis, Knee|Disorder|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|knee osteoarthritisnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|kneenull|Knee region structure|Anatomy|false|false|C1552822;C0562271;C1549543;C0030193;C0409959;C0029408|knee
null|Knee|Anatomy|false|false|C1552822;C0562271;C1549543;C0030193;C0409959;C0029408|knee
null|Lower extremity>Knee|Anatomy|false|false|C1552822;C0562271;C1549543;C0030193;C0409959;C0029408|knee
null|Knee joint|Anatomy|false|false|C1552822;C0562271;C1549543;C0030193;C0409959;C0029408|kneenull|Degenerative polyarthritis|Disorder|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|osteoarthritisnull|Administration Method - Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|pain
null|Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|painnull|null|Attribute|false|false||painnull|Measures (attribute)|Finding|false|false||measuresnull|Measures|LabModifier|false|false||measuresnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Total|Modifier|false|false||totalnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C0562271|knee
null|Knee|Anatomy|false|false|C0562271|knee
null|Lower extremity>Knee|Anatomy|false|false|C0562271|knee
null|Knee joint|Anatomy|false|false|C0562271|kneenull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false||arthroplasty
null|Arthroplasty|Procedure|false|false||arthroplasty
null|Reconstruction of joint|Procedure|false|false||arthroplastynull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false|C0042449|varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false|C0042449|veinsnull|Veins|Anatomy|false|false|C0042345;C0398102|veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEs
null|PES1 gene|Finding|false|false|C1690938;C3853547;C0687080;C0016504|PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false|C4551530;C1418467;C0687136|PEs
null|Hindfoot of quadruped|Anatomy|false|false|C4551530;C1418467;C0687136|PEs
null|Paw|Anatomy|false|false|C4551530;C1418467;C0687136|PEs
null|Foot|Anatomy|false|false|C4551530;C1418467;C0687136|PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false|C1167408;C3665580|antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false|C1167408;C3665580|antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false|C1167408;C3665580|antiphospholipid antibodynull|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Immunoglobulins|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibody
null|Antibodies|Drug|false|false|C1167408;C3665580|antibodynull|Antibody (immunoassay)|Procedure|false|false|C1167408;C3665580;C1690938;C3853547;C0687080;C0016504|antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false|C4551530;C0162595;C4019436;C0003241;C0021027;C0085278;C0039082|antibody
null|immunoglobulin complex location|Anatomy|false|false|C4551530;C0162595;C4019436;C0003241;C0021027;C0085278;C0039082|antibodynull|Syndrome|Disorder|false|false|C1167408;C3665580|syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false|C0228174;C0006104|A1Cnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false|C0474680|cerebral
null|Brain|Anatomy|false|false|C0474680|cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|true|false|C0009368;C4071907|colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|true|false|C0009368;C4071907|colon
null|Colonic Diseases|Disorder|true|false|C0009368;C4071907|colon
null|Carcinoma in situ of colon|Disorder|true|false|C0009368;C4071907|colonnull|COLON PROBLEM|Finding|true|false|C0009368;C4071907|colonnull|Colon structure (body structure)|Anatomy|false|false|C0009376;C0032584;C0009373;C0154061;C0496907;C0750873|colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false|C0009376;C0032584;C0009373;C0154061;C0496907;C0750873|colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|true|false||colonnull|Colon <Coloninae>|Entity|true|false||colonnull|polyps|Disorder|false|false|C0009368;C4071907|polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false|C3890599|CMC
null|Capillary malformation (disorder)|Disorder|false|false|C3890599|CMCnull|MCC protocol|Procedure|false|false|C3890599|CMCnull|Circulating Melanoma Cell|Anatomy|false|false|C0065772;C0006845;C0340803|CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false|C0392905;C1269611;C0022417|joint arthroplastynull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417|jointnull|null|Anatomy|false|false|C5887062;C0003893;C0700235;C0575044;C0003893|joint
null|Joints|Anatomy|false|false|C5887062;C0003893;C0700235;C0575044;C0003893|joint
null|Articular system|Anatomy|false|false|C5887062;C0003893;C0700235;C0575044;C0003893|jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false|C0392905;C1269611;C0022417|arthroplasty
null|Arthroplasty|Procedure|false|false|C0392905;C1269611;C0022417|arthroplasty
null|Reconstruction of joint|Procedure|false|false|C0392905;C1269611;C0022417|arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false|C0085515;C1550244|rotator cuff repairnull|Rotator Cuff|Anatomy|false|false|C0186666;C0374711;C1705181;C3668885;C0015252;C0728940;C0043240;C4319951|rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false|C1550244;C0085515|cuffnull|Cuff - body part|Anatomy|false|false|C3668885;C0186666|cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false|C0085515|repair
null|Wound Healing|Finding|false|false|C0085515|repairnull|Repair - Remedial Action|Procedure|false|false|C0085515|repair
null|Surgical repair|Procedure|false|false|C0085515|repairnull|Excision|Procedure|false|false|C0085515|excision
null|removal technique|Procedure|false|false|C0085515|excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false|C0582802|digitnull|Digit structure|Anatomy|false|false|C4283905;C1546709;C2700045;C0577573;C0577559;C1414542;C4761764|digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false|C0582802|mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false|C0582802|mass
null|null|Finding|false|false|C0582802|mass
null|FBN1 wt Allele|Finding|false|false|C0582802|mass
null|FBN1 gene|Finding|false|false|C0582802|mass
null|Mass of body region|Finding|false|false|C0582802|massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false|C4482304;C0030288;C0030274;C0687028;C1550227|pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic duct
null|Pancreatic duct|Anatomy|false|false|C0153461;C1280903|pancreatic ductnull|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreatic
null|Pancreatic Hormones|Drug|false|false|C0030274|pancreaticnull|Pancreas|Anatomy|false|false|C0153461;C0030292|pancreaticnull|Duct (organ) structure|Anatomy|false|false|C0153461|duct
null|canal [body parts]|Anatomy|false|false|C0153461|ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false|C4482304;C0030288|explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Entity Name Part Type - family|Finding|false|false|C5239664|family
null|Last Name|Finding|false|false|C5239664|family
null|Living Arrangement - Family|Finding|false|false|C5239664|family
null|Family (taxonomic)|Finding|false|false|C5239664|family
null|Family Collection|Finding|false|false|C5239664|familynull|Family|Subject|false|false||familynull|Deep thrombophlebitis|Disorder|true|false|C5239664|DVT
null|Deep Vein Thrombosis|Disorder|true|false|C5239664|DVTnull|area DVT|Anatomy|false|false|C0149871;C0151950;C2700055;C1546847;C1704727;C1301584;C1563343;C2926618|DVTnull|null|Attribute|true|false|C5239664|DVTnull|Sister|Subject|false|false||sistersnull|Atrial Fibrillation|Disorder|false|false|C0018792|atrial fibrillationnull|null|Attribute|false|false|C0018792|atrial fibrillationnull|Atrial Fibrillation by ECG Finding|Lab|false|false|C0018792|atrial fibrillationnull|Heart Atrium|Anatomy|false|false|C0344434;C0004238;C0232197;C2926591|atrialnull|Fibrillation|Disorder|false|false|C0018792|fibrillationnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Apyrexial|Finding|false|false||Afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Respiratory attachment|Finding|false|false||Respiratory
null|respiratory|Finding|false|false||Respiratory
null|null|Finding|false|false||Respiratory
null|Respiratory specimen|Finding|false|false||Respiratorynull|Respiratory rate|Attribute|false|false||Respiratorynull|cetrimonium bromide|Drug|false|false||CTABnull|Cardiovascular system|Anatomy|false|false||Cardiovascular
null|Cardiovascular|Anatomy|false|false||Cardiovascularnull|Gastrointestinal attachment|Finding|false|false||Gastrointestinalnull|gastrointestinal|Modifier|false|false||Gastrointestinalnull|Genitourinary Route of Administration|Finding|false|false|C3887515;C0042066|Genitourinarynull|Genitourinary system|Anatomy|false|false|C2709258|Genitourinary
null|Genitourinary|Anatomy|false|false|C2709258|Genitourinarynull|Urination|Finding|false|false||Voiding
null|Voids|Finding|false|false||Voidingnull|Neurologic (qualifier value)|Modifier|false|false||Neurologicnull|Gender Status - Intact|Finding|false|false||Intactnull|Intact|Modifier|false|false||Intactnull|Focal|Modifier|false|false||focalnull|Deficit|Modifier|false|false||deficitsnull|Referral type - Psychiatric|Finding|false|false||Psychiatric
null|Psychiatric|Finding|false|false||Psychiatricnull|Psychiatric service|Procedure|false|false||Psychiatricnull|Psychiatry Specialty|Title|false|false||Psychiatricnull|Pleasant|Finding|false|false||Pleasantnull|Musculoskeletal|Finding|false|false|C1548802;C0023216|Musculoskeletalnull|null|Attribute|false|false|C0023216|Musculoskeletalnull|Lower Extremity|Anatomy|false|false|C0497254;C2707260|Lower Extremitynull|Body Site Modifier - Lower|Anatomy|false|false|C0497254;C2003888|Lowernull|Lower (action)|Event|false|false|C1548802|Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Limb structure|Anatomy|false|false||Extremitynull|DRESSING,AQUACEL|Device|false|false||Aquacel dressingnull|Aquacel|Drug|false|false||Aquacelnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Scant|Finding|false|false||scantnull|Smallest|LabModifier|false|false||scantnull|Serosanguineous|Modifier|false|false||serosanguinousnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Full|Modifier|false|false||fullnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|CALF TENDERNESS|Finding|true|false|C0230445;C1305418|calf tendernessnull|Structure of calf of leg|Anatomy|false|false|C0684239;C0234233;C0238883|calf
null|null|Anatomy|false|false|C0684239;C0234233;C0238883|calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Emotional tenderness|Finding|true|false|C0230445;C1305418|tenderness
null|Sore to touch|Finding|true|false|C0230445;C1305418|tendernessnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Lower extremity>Toes|Anatomy|false|false|C0687712;C0582051|Toes
null|Toes|Anatomy|false|false|C0687712;C0582051|Toesnull|Feels warm|Finding|false|false|C0040357;C4299090|warmnull|warming process|Phenomenon|false|false|C0040357;C4299090|warmnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Mandibular right first molar abutment mesial hemisection|Device|false|false||30AMnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Orthopedic Surgical Procedures|Procedure|false|false||Orthopaedic surgerynull|Orthopedics|Title|false|false||Orthopaedicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Operating Room|Device|false|false||operating roomnull|Operating Room|Entity|false|false||operating roomnull|Patient location type - Operating Room|Modifier|false|false||operating roomnull|Operating|Finding|false|false||operatingnull|Room - Patient location type|Modifier|false|false||room
null|Room|Modifier|false|false||roomnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Operative report|Finding|false|false||operative reportnull|Operative|Time|false|false||operativenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Details|Modifier|false|false||detailsnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Uncomplicated|Modifier|false|false||uncomplicatednull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|perioperative|Time|false|false||perioperativenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Postoperative Period|Time|false|false||Postoperativenull|Course|Time|false|false||coursenull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Bolus of ingested food|Finding|false|false||bolus
null|Response Modality - Bolus|Finding|false|false||bolusnull|bolus infusion|Procedure|false|false||bolusnull|Bolus Dosing Unit|LabModifier|false|false||bolusnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Hypotension|Finding|false|false||hypotensionnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|aspects of adverse effects|Finding|false|false||adverse effects
null|Adverse effects|Finding|false|false||adverse effectsnull|Effect|Modifier|false|false||effectsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Lovenox|Drug|false|false||lovenox
null|Lovenox|Drug|false|false||lovenoxnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Daily|Time|false|false||dailynull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Check|Finding|false|false||checknull|null|Event|false|false||checknull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Direct - PostalAddressUse|Finding|false|false||direct
null|direct address|Finding|false|false||directnull|Direct type of relationship|Modifier|false|false||direct
null|Direct (qualifier)|Modifier|false|false||directnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|combination - answer to question|Finding|false|false|C0226896|combinationnull|combination of objects|Entity|false|false||combinationnull|Combined|Modifier|false|false||combinationnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C3811910;C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Daily|Time|false|false||dailynull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Levels (qualifier value)|Modifier|false|false||levelsnull|SURGICAL DRESSINGS|Device|false|false||surgical dressingnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Surgical procedure finding|Finding|false|false||surgery
null|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Daily|Time|false|false||dailynull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Laboratory test finding|Lab|false|false||Labsnull|Hospital course|Finding|false|false||hospital coursenull|null|Attribute|false|false||hospital coursenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Course|Time|false|false||coursenull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Hematocrit level|Finding|false|false||hematocritnull|Hematocrit Measurement|Procedure|false|false||hematocritnull|hematocrit attribute|Attribute|false|false||hematocritnull|Acceptable (foundation metadata concept)|Modifier|false|false||acceptable
null|Acceptable|Modifier|false|false||acceptablenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Operative|Time|false|false||operativenull|Limb structure|Anatomy|false|false||extremitynull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Weight-Bearing state|Subject|false|false||weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||weight
null|Weight symptom (finding)|Finding|false|false||weightnull|Weighing patient|Procedure|false|false||weightnull|null|Attribute|false|false||weightnull|Body Weight|Subject|false|false||weightnull|Importance Weight|Modifier|false|false||weightnull|Weight|LabModifier|false|false||weightnull|Bearing Device|Device|false|false||bearingnull|Operative|Time|false|false||operativenull|Limb structure|Anatomy|false|false||extremitynull|instruction in use of walker|Procedure|false|false||use walkernull|Walkers|Device|false|false||walkernull|Crutches|Device|false|false||crutchesnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Rehabilitation therapy|Procedure|false|false||rehabnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Rehab facility|Device|false|false||rehab facilitynull|Rehab facility|Entity|false|false||rehab facilitynull|Rehabilitation therapy|Procedure|false|false||rehabnull|ADMIN.FACILITY|Finding|false|false||facilitynull|Facility (object)|Device|false|false||facilitynull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|30 days|Time|false|false||30 daysnull|day|Time|false|false||daysnull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Wheezing|Finding|false|false||wheezingnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|econazole|Drug|false|false||econazole
null|econazole|Drug|false|false||econazolenull|Topical Dosage Form|Drug|false|false||topicalnull|Topical Route of Administration|Finding|false|false||topicalnull|Topical surface|Modifier|false|false||topicalnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|enoxaparin sodium|Drug|false|false||Enoxaparin Sodium
null|enoxaparin sodium|Drug|false|false||Enoxaparin Sodiumnull|enoxaparin|Drug|false|false||Enoxaparin
null|enoxaparin|Drug|false|false||Enoxaparinnull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Every twelve hours|Time|false|false||Q12Hnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|next - HtmlLinkType|Finding|false|false||Nextnull|Following|Time|false|false||Next
null|Then|Time|false|false||Nextnull|Adjacent|Modifier|false|false||Nextnull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Administration (procedure)|Procedure|false|false||Administrationnull|Administration occupational activities|Event|false|false||Administrationnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||Time
null|Time (foundation metadata concept)|Finding|false|false||Time
null|Value type - Time|Finding|false|false||Time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||Time
null|Data types - Time|Finding|false|false||Time
null|null|Finding|false|false||Timenull|Time|Time|false|false||Timenull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|leg swellingnull|Leg|Anatomy|false|false|C0581394|leg
null|Lower Extremity|Anatomy|false|false|C0581394|legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|metformin|Drug|false|false||MetFORMIN
null|metformin|Drug|false|false||MetFORMINnull|Glucophage|Drug|false|false||Glucophage
null|Glucophage|Drug|false|false||Glucophagenull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonide
null|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonidenull|triamcinolone|Drug|false|false||Triamcinolone
null|triamcinolone|Drug|false|false||Triamcinolonenull|Ointments|Drug|false|false||Ointmentnull|APPL1 gene|Finding|false|false||Applnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Pruritus|Finding|false|false||itchingnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|hydromorphone|Drug|false|false||HYDROmorphone
null|hydromorphone|Drug|false|false||HYDROmorphonenull|Dilaudid|Drug|false|false||Dilaudid
null|Dilaudid|Drug|false|false||Dilaudidnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Multiple Epiphyseal Dysplasia|Disorder|false|false||mednull|Master of Education|Finding|false|false||med
null|COMP wt Allele|Finding|false|false||med
null|COL9A3 gene|Finding|false|false||med
null|SCN8A wt Allele|Finding|false|false||med
null|COL9A2 gene|Finding|false|false||med
null|COMP gene|Finding|false|false||med
null|SCN8A gene|Finding|false|false||mednull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Daily|Time|false|false||DAILYnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Daily|Time|false|false||DAILYnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|objective (goal)|Finding|false|false||GOAL
null|Act Mood - Goal|Finding|false|false||GOALnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Inhaler (unit of presentation)|Finding|false|false||Inhalernull|Inhaler|Device|false|false||Inhalernull|Inhaler Dosing Unit|LabModifier|false|false||Inhalernull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Dyspnea|Finding|false|false||shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false||breathnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|econazole|Drug|false|false||econazole
null|econazole|Drug|false|false||econazolenull|Topical Dosage Form|Drug|false|false||topicalnull|Topical Route of Administration|Finding|false|false||topicalnull|Topical surface|Modifier|false|false||topicalnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false|C1140621;C0023216|leg swellingnull|Leg|Anatomy|false|false|C0581394|leg
null|Lower Extremity|Anatomy|false|false|C0581394|legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|metformin|Drug|false|false||MetFORMIN
null|metformin|Drug|false|false||MetFORMINnull|Glucophage XR|Drug|false|false||Glucophage XR
null|Glucophage XR|Drug|false|false||Glucophage XRnull|Glucophage|Drug|false|false||Glucophage
null|Glucophage|Drug|false|false||Glucophagenull|Daily|Time|false|false||DAILYnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonide
null|triamcinolone acetonide|Drug|false|false||Triamcinolone Acetonidenull|triamcinolone|Drug|false|false||Triamcinolone
null|triamcinolone|Drug|false|false||Triamcinolonenull|Ointments|Drug|false|false||Ointmentnull|APPL1 gene|Finding|false|false||Applnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Eruption of skin (disorder)|Disorder|false|false||rashnull|Skin rash|Finding|false|false||rash
null|Eruptions|Finding|false|false||rash
null|Exanthema|Finding|false|false||rashnull|Pruritus|Finding|false|false||itchingnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|long-term care|Procedure|false|false||Extended Carenull|Extended (finding)|Finding|false|false||Extended
null|Extension|Finding|false|false||Extendednull|Extended|Modifier|false|false||Extended
null|Extent|Modifier|false|false||Extendednull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Structure of left knee region|Anatomy|false|false|C1552822;C0409959;C0562271;C0029408;C1549543;C0030193|left knee
null|Structure of left knee|Anatomy|false|false|C1552822;C0409959;C0562271;C0029408;C1549543;C0030193|left kneenull|Table Cell Horizontal Align - left|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Osteoarthritis, Knee|Disorder|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|knee osteoarthritisnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|kneenull|Knee region structure|Anatomy|false|false|C0562271;C0029408;C1552822;C1549543;C0030193;C0409959|knee
null|Knee|Anatomy|false|false|C0562271;C0029408;C1552822;C1549543;C0030193;C0409959|knee
null|Lower extremity>Knee|Anatomy|false|false|C0562271;C0029408;C1552822;C1549543;C0030193;C0409959|knee
null|Knee joint|Anatomy|false|false|C0562271;C0029408;C1552822;C1549543;C0030193;C0409959|kneenull|Degenerative polyarthritis|Disorder|false|false|C1963703;C0022742;C4299094;C0022745;C0230432;C4281599|osteoarthritisnull|Administration Method - Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|pain
null|Pain|Finding|false|false|C0230432;C4281599;C1963703;C0022742;C4299094;C0022745|painnull|null|Attribute|false|false||painnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Accident and Emergency department|Device|false|false||emergency departmentnull|interventional services emergency department|Entity|false|false||emergency department
null|Accident and Emergency department|Entity|false|false||emergency departmentnull|Consent Non-Disclosure Reason - Emergency|Finding|false|false||emergency
null|Admission Type - Emergency|Finding|false|false||emergency
null|Referral category - Emergency|Finding|false|false||emergency
null|Emergencies [Disease/Finding]|Finding|false|false||emergency
null|Consent Bypass Reason - Emergency|Finding|false|false||emergency
null|Level of Care - Emergency|Finding|false|false||emergency
null|Certification patient type - Emergency|Finding|false|false||emergency
null|Encounter Admission Source - emergency|Finding|false|false||emergency
null|Patient Class - Emergency|Finding|false|false||emergency
null|Visit Priority Code - Emergency|Finding|false|false||emergencynull|emergency encounter|Procedure|false|false||emergencynull|Specialty Type - Emergency|Title|false|false||emergencynull|Emergency Situation|Phenomenon|false|false||emergencynull|Bale out|Time|false|false||emergencynull|Department - No suggested values defined|Finding|false|false||department
null|Organization Unit Type - Department|Finding|false|false||department
null|Department - Charge type|Finding|false|false||departmentnull|Department|Entity|false|false||departmentnull|Patient location type - Department|Modifier|false|false||department
null|Department - Person location type|Modifier|false|false||departmentnull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Following|Time|false|false||following
null|Status post|Time|false|false||followingnull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Difficult (qualifier value)|Finding|false|false||difficulty withnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Movement|Finding|false|false||movementnull|Fever|Finding|false|false||feversnull|Greater Than|LabModifier|false|false||greater thannull|Greater|LabModifier|false|false||greaternull|Chills|Finding|false|false||chillsnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0741025;C0225386;C1546778;C0013404;C0008031;C1549543;C0030193|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Chest Pain|Finding|false|false|C1527391;C0817096;C1515974|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1515974;C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false|C1515974|pain
null|Pain|Finding|false|false|C1515974|painnull|null|Attribute|false|false||painnull|Dyspnea|Finding|false|false|C1515974|shortness of breathnull|null|Attribute|false|false||shortness of breathnull|Breath|Finding|false|false|C1515974|breathnull|Primary physician|Subject|false|false||primary physiciannull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|New medications|Drug|false|false||new medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|refill|Finding|false|false||refillsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|heavy machinery|Device|false|false||heavy machinerynull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Contact with machinery|Disorder|false|false||machinerynull|Industrial machine|Device|false|false||machinerynull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Tablet Dosage Form|Drug|false|false||tabletsnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Dosage|LabModifier|false|false||dosesnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Constipation|Finding|false|false||constipationnull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false||waternull|Daily|Time|false|false||dailynull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||Colace
null|Colace|Drug|false|false||Colacenull|PREVENT (product)|Drug|false|false||preventnull|Adverse effects|Finding|false|false||side effectnull|Side|Modifier|false|false||sidenull|Effect, Appearance|Modifier|false|false||effect
null|Effect|Modifier|false|false||effectnull|Surgeon|Subject|false|false||surgeonsnull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Diagnostic Service Section ID - Pharmacy|Finding|false|false||pharmacy
null|Pharmacy domain|Finding|false|false||pharmacynull|Pharmaceutical Services|Procedure|false|false||pharmacynull|Pharmacy facility|Device|false|false||pharmacynull|Pharmacy (field)|Title|false|false||pharmacynull|Pharmacy facility|Entity|false|false||pharmacynull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|2 Days|Time|false|false||2 daysnull|day|Time|false|false||daysnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Coxsackievirus and Adenovirus Receptor, human|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Chimeric antigen receptor|Drug|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Drug|false|false|C1166663|carnull|Carney Complex|Disorder|false|false|C1166663|carnull|Car - Mode of Arrival Code|Finding|false|false|C1166663|car
null|Chimeric antigen receptor|Finding|false|false|C1166663|car
null|CASR wt Allele|Finding|false|false|C1166663|car
null|Extracellular Calcium-Sensing Receptor, Human|Finding|false|false|C1166663|car
null|CXADR wt Allele|Finding|false|false|C1166663|car
null|CXADR gene|Finding|false|false|C1166663|car
null|PRKAR1A wt Allele|Finding|false|false|C1166663|car
null|CXADRP1 gene|Finding|false|false|C1166663|car
null|NR1I3 gene|Finding|false|false|C1166663|car
null|SPG7 gene|Finding|false|false|C1166663|car
null|TRIM13 wt Allele|Finding|false|false|C1166663|car
null|Caronte Gene|Finding|false|false|C1166663|car
null|SPG7 wt Allele|Finding|false|false|C1166663|car
null|NR1I3 wt Allele|Finding|false|false|C1166663|carnull|actomyosin contractile ring|Anatomy|false|false|C3540475;C1547285;C3273602;C4039583;C1413828;C3811749;C2239319;C1858724;C1417827;C5890847;C1420354;C5960871;C1706434;C5890846;C0406810;C3539542;C4039583;C5890846|carnull|Automobiles|Device|false|false||carnull|Car <Caridae>|Entity|false|false||car
null|Carib language|Entity|false|false||carnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Address type - Office|Finding|false|false||officenull|Office|Device|false|false||officenull|Organization unit type - Office|Entity|false|false||officenull|Appointments|Event|false|false||appointmentnull|Swelling|Finding|false|false||SWELLING
null|Edema|Finding|false|false||SWELLINGnull|Operative|Time|false|false||operativenull|Joint problem|Finding|false|false|C0392905;C1269611;C0022417|jointnull|null|Anatomy|false|false|C0575044;C5575590;C2024467;C1548318;C1547403;C3541383;C5400024|joint
null|Joints|Anatomy|false|false|C0575044;C5575590;C2024467;C1548318;C1547403;C3541383;C5400024|joint
null|Articular system|Anatomy|false|false|C0575044;C5575590;C2024467;C1548318;C1547403;C3541383;C5400024|jointnull|Joint Device|Device|false|false||jointnull|20 minutes|Time|false|false||20 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|Instructions for Use of the CPT Codebook - Time|Finding|false|false|C0392905;C1269611;C0022417|time
null|Time (foundation metadata concept)|Finding|false|false|C0392905;C1269611;C0022417|time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false|C0392905;C1269611;C0022417|time
null|Value type - Time|Finding|false|false|C0392905;C1269611;C0022417|time
null|Data types - Time|Finding|false|false|C0392905;C1269611;C0022417|time
null|null|Finding|false|false|C0392905;C1269611;C0022417|timenull|Time|Time|false|false||timenull|Physical activity|Finding|false|false||activity
null|Activity (animal life circumstance)|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Ice Pharmaceutical|Drug|false|false|C3496566;C0228434|ice
null|Ice Pharmaceutical|Drug|false|false|C3496566;C0228434|ice
null|Ice|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|methamphetamine|Drug|false|false|C3496566;C0228434|ice
null|Caspase-1, human|Drug|false|false|C3496566;C0228434|ice
null|Caspase-1, human|Drug|false|false|C3496566;C0228434|icenull|caspase-1 activity|Finding|false|false|C3496566;C0228434|ice
null|CASP1 wt Allele|Finding|false|false|C3496566;C0228434|ice
null|CES2 gene|Finding|false|false|C3496566;C0228434|ice
null|CES2 wt Allele|Finding|false|false|C3496566;C0228434|ice
null|CASP1 gene|Finding|false|false|C3496566;C0228434|icenull|cryotherapy using ice|Procedure|false|false|C3496566;C0228434|ice
null|cytarabine/etoposide/idarubicin|Procedure|false|false|C3496566;C0228434|ice
null|AIE Regimen|Procedure|false|false|C3496566;C0228434|ice
null|carboplatin/etoposide/ifosfamide|Procedure|false|false|C3496566;C0228434|icenull|Structure of inferior central nucleus of pons|Anatomy|false|false|C0249492;C1879508;C0280697;C0556917;C0020746;C1873773;C4721557;C0025611;C1705786;C3889432;C1366479;C1150137;C1413348|ice
null|intracentral fissure|Anatomy|false|false|C0249492;C1879508;C0280697;C0556917;C0020746;C1873773;C4721557;C0025611;C1705786;C3889432;C1366479;C1150137;C1413348|icenull|Direct (qualifier)|Modifier|false|false||directlynull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|skinnull|Examination of knee joint|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|kneenull|Knee region structure|Anatomy|false|false|C0050385;C0279078;C0108844;C1879921;C0562271|knee
null|Knee|Anatomy|false|false|C0050385;C0279078;C0108844;C1879921;C0562271|knee
null|Lower extremity>Knee|Anatomy|false|false|C0050385;C0279078;C0108844;C1879921;C0562271|knee
null|Knee joint|Anatomy|false|false|C0050385;C0279078;C0108844;C1879921;C0562271|kneenull|Ace Bandages|Device|false|false||ace bandagenull|ACE protein, human|Drug|false|false||ace
null|ACE protein, human|Drug|false|false||acenull|ACE gene|Finding|false|false||ace
null|Adverse Childhood Experience questionnaire|Finding|false|false||acenull|cisplatin, cytarabine, and etoposide chemotherapy protocol|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|ace
null|cyclophosphamide/doxorubicin protocol|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|ace
null|CDE protocol|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|ace
null|CDE Regimen|Procedure|false|false|C1963703;C0022742;C4299094;C0022745|acenull|Achinese language|Entity|false|false||acenull|Bandage Dosage Form|Drug|false|false||bandagenull|Bandage|Device|false|false||bandagenull|Additional|Finding|false|false||addednull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Anti-Inflammatory Agents|Drug|false|false||anti-inflammatorynull|Anti-inflammatory effect|Modifier|false|false||anti-inflammatorynull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Analgesics and non-steroidal anti-inflammatory drugs|Drug|false|false||NSAIDs
null|Anti-Inflammatory Agents, Non-Steroidal|Drug|false|false||NSAIDsnull|Celebrex|Drug|false|false||Celebrex
null|Celebrex|Drug|false|false||Celebrexnull|ibuprofen|Drug|false|false||ibuprofen
null|ibuprofen|Drug|false|false||ibuprofennull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|Aleve|Drug|false|false||Aleve
null|Aleve|Drug|false|false||Alevenull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|naproxen|Drug|false|false||naproxen
null|naproxen|Drug|false|false||naproxennull|Etc.|Finding|false|false||etcnull|null|Attribute|false|false||physiciannull|Physicians|Subject|false|false||physiciannull|ANTICOAGULATION (finding)|Finding|false|false||ANTICOAGULATION
null|Anticoagulation function|Finding|false|false||ANTICOAGULATION
null|Decreased Coagulation Activity [PE]|Finding|false|false||ANTICOAGULATIONnull|Anticoagulation Therapy|Procedure|false|false||ANTICOAGULATIONnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Coagulation tissue factor induced.INR goal|Attribute|false|false||INR goalnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Daily|Time|false|false||dailynull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Direct - PostalAddressUse|Finding|false|false||direct
null|direct address|Finding|false|false||directnull|Direct type of relationship|Modifier|false|false||direct
null|Direct (qualifier)|Modifier|false|false||directnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||dailynull|Wound care management|Procedure|false|false||WOUND CARE
null|wound care|Procedure|false|false||WOUND CAREnull|Wound Care kit|Device|false|false||WOUND CAREnull|Traumatic Wound|Disorder|false|false||WOUND
null|Wounds and Injuries|Disorder|false|false||WOUND
null|Traumatic injury|Disorder|false|false||WOUNDnull|Route of Administration - Wound|Finding|false|false||WOUND
null|null|Finding|false|false||WOUND
null|Specimen Type - Wound|Finding|false|false||WOUNDnull|In care (finding)|Finding|false|false||CARE
null|Continuity Assessment Record and Evaluation|Finding|false|false||CAREnull|care activity|Event|false|false||CAREnull|DRESSING,AQUACEL|Device|false|false||Aquacel dressingnull|Aquacel|Drug|false|false||Aquacelnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|5 Days|Time|false|false||5 daysnull|day|Time|false|false||daysnull|TUB gene|Finding|false|false||tubnull|Tub - container|Device|false|false||tubnull|Tub Dosing Unit|LabModifier|false|false||tubnull|Bathing|Procedure|false|false||bathsnull|Baths (medical device)|Device|false|false||bathsnull|swimming (history)|Finding|false|false||swimming
null|Swimming|Finding|false|false||swimmingnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0184898;C0332803|incisionnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|checkup examination|Procedure|false|false||checkupnull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Daily|Time|false|false||each daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Open|Modifier|false|false||opennull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Thick|Modifier|false|false||thicknull|Yellow color|Modifier|false|false||yellownull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic Wound|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Activity (animal life circumstance)|Finding|false|false||ACTIVITY
null|Physical activity|Finding|false|false||ACTIVITYnull|Activities|Event|false|false||ACTIVITYnull|null|Modifier|false|false||ACTIVITYnull|Weight-Bearing state|Subject|false|false||Weight bearingnull|infant weight for previous delivery (history)|Finding|false|false||Weight
null|Weight symptom (finding)|Finding|false|false||Weightnull|Weighing patient|Procedure|false|false||Weightnull|null|Attribute|false|false||Weightnull|Body Weight|Subject|false|false||Weightnull|Importance Weight|Modifier|false|false||Weightnull|Weight|LabModifier|false|false||Weightnull|Bearing Device|Device|false|false||bearingnull|Operative|Time|false|false||operativenull|Limb structure|Anatomy|false|false||extremitynull|Crutches|Device|false|false||crutchesnull|Walkers|Device|false|false||walkernull|Self-Help Devices|Device|false|false||assistive devicenull|Participation Type - device|Finding|false|false||devicenull|Medical Devices|Device|false|false||device
null|Devices|Device|false|false||devicenull|Kind of quantity - Device|LabModifier|false|false||devicenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Does mobilize|Finding|false|false||Mobilizenull|Mobilization (procedure)|Procedure|false|false||Mobilizenull|Rupture of Membranes|Finding|false|false||ROM
null|ROM1 gene|Finding|false|false||ROMnull|Range of motion technique (procedure)|Procedure|false|false||ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Strenuous Exercise|Finding|true|false||strenuous exercisenull|Strenuous|Modifier|false|false||strenuousnull|Exercise|Finding|true|false||exercisenull|Exercise Pain Management|Procedure|true|false||exercisenull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|false|false||liftingnull|Follow-up status|Finding|false|false||follow upnull|follow-up|Procedure|false|false||follow upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||Physical Therapynull|Physical therapy|Procedure|false|false||Physical Therapynull|Physical therapy (field)|Title|false|false||Physical Therapynull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Therapy Object (animal model)|Finding|false|false||Therapy
null|therapeutic aspects|Finding|false|false||Therapynull|Therapeutic procedure|Procedure|false|false||Therapynull|Range of motion restrictions|Finding|true|false||range of motion restrictionsnull|Range of motion exercise|Procedure|true|false||range of motionnull|Range of Motion, Articular|Attribute|true|false||range of motionnull|Concept model range (foundation metadata concept)|Finding|true|false||rangenull|Sample Range|LabModifier|false|false||range
null|Range|LabModifier|false|false||rangenull|Motion|Phenomenon|false|false||motionnull|Self-Help Devices|Device|false|false||assistive devicesnull|Medical Devices|Device|false|false||devices
null|device aspects|Device|false|false||devices
null|Devices|Device|false|false||devicesnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Does mobilize|Finding|false|false||Mobilizenull|Mobilization (procedure)|Procedure|false|false||Mobilizenull|Frequently|Time|false|false||frequentlynull|Therapeutic procedure|Procedure|false|false||Treatmentsnull|Frequency|Finding|false|false||Frequency
null|How Often|Finding|false|false||Frequencynull|With frequency|Time|false|false||Frequency
null|Frequencies (time pattern)|Time|false|false||Frequencynull|Kind of quantity - Frequency|LabModifier|false|false||Frequency
null|Statistical Frequency|LabModifier|false|false||Frequency
null|Spatial Frequency|LabModifier|false|false||Frequencynull|Aquacel|Drug|false|false||aquacelnull|post operative (finding)|Finding|false|false||after surgerynull|Postoperative Period|Time|false|false||after surgerynull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Sterility, Reproductive|Finding|false|false||sterile
null|Infertility|Finding|false|false||sterilenull|Sterile (qualifier value)|Modifier|false|false||sterilenull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Daily|Time|false|false||dailynull|Aquacel|Drug|false|false||aquacelnull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Daily|Time|false|false||dailynull|Aquacel|Drug|false|false||aquacelnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions