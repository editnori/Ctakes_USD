 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|155,163|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|178,185|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|Allergies|178,185|false|false|false|C0009214|codeine|Codeine
Drug|Antibiotic|Allergies|188,197|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|188,197|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|Allergies|200,207|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|Allergies|200,207|false|false|false|C0723778|Topamax|Topamax
Finding|Functional Concept|Allergies|210,219|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|Chief Complaint|249,253|false|false|false|C2598155||pain
Finding|Functional Concept|Chief Complaint|249,253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Chief Complaint|249,253|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Chief Complaint|258,266|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Chief Complaint|258,266|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Classification|Chief Complaint|269,274|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|287,305|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|296,305|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|296,305|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|296,305|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|296,305|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|307,317|false|false|false|C0220934|Ultrasonic|Ultrasound
Phenomenon|Natural Phenomenon or Process|Chief Complaint|307,317|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|Ultrasound
Procedure|Diagnostic Procedure|Chief Complaint|307,317|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|Ultrasound
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|307,342|false|false|false|C4305575|Ultrasonography guided steroid injection|Ultrasound guided steroid injection
Drug|Organic Chemical|Chief Complaint|325,332|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Chief Complaint|325,332|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|325,342|false|false|false|C1261311|Injection of steroid|steroid injection
Drug|Biomedical or Dental Material|Chief Complaint|333,342|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|Chief Complaint|333,342|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|333,342|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Functional Concept|Chief Complaint|350,355|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|370,375|false|false|false|C0006441|Synovial bursa|bursa
Finding|Functional Concept|Chief Complaint|377,382|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Chief Complaint|377,386|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|383,386|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Chief Complaint|383,386|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Chief Complaint|383,386|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Chief Complaint|383,386|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Chief Complaint|383,386|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|383,386|false|false|false|C1292890|Procedure on hip|hip
Finding|Conceptual Entity|History of Present Illness|446,453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|446,453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|446,453|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|446,456|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|457,463|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|457,463|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|457,463|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|457,463|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|History of Present Illness|457,470|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|History of Present Illness|464,470|false|false|false|C0006826|Malignant Neoplasms|cancer
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|476,481|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|History of Present Illness|476,481|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Finding|Gene or Genome|History of Present Illness|476,481|false|false|false|C0376571|BRCA1 gene|BRCA1
Finding|Gene or Genome|History of Present Illness|476,486|false|false|false|C0376571|BRCA1 gene|BRCA1 gene
Procedure|Laboratory Procedure|History of Present Illness|476,486|false|false|false|C2010863|BRCA1 gene (lab test)|BRCA1 gene
Disorder|Cell or Molecular Dysfunction|History of Present Illness|476,495|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 gene mutation
Finding|Finding|History of Present Illness|482,486|false|false|false|C0017337;C5849123|Genes;Gross Extranodal Extension|gene
Finding|Gene or Genome|History of Present Illness|482,486|false|false|false|C0017337;C5849123|Genes;Gross Extranodal Extension|gene
Finding|Gene or Genome|History of Present Illness|482,495|false|false|false|C0596611;C0678941|Gene Mutant;Gene Mutation|gene mutation
Finding|Genetic Function|History of Present Illness|482,495|false|false|false|C0596611;C0678941|Gene Mutant;Gene Mutation|gene mutation
Disorder|Cell or Molecular Dysfunction|History of Present Illness|487,495|false|false|false|C1705285|Mutation Abnormality|mutation
Finding|Genetic Function|History of Present Illness|487,495|false|false|false|C0026882|Mutation|mutation
Disorder|Disease or Syndrome|History of Present Illness|497,501|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|497,501|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|History of Present Illness|497,501|false|false|false|C1412502|ARCN1 gene|COPD
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|503,511|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|History of Present Illness|503,520|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Finding|Pathologic Function|History of Present Illness|512,520|false|false|false|C0002940|Aneurysm|aneurysm
Drug|Organic Chemical|History of Present Illness|522,527|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|History of Present Illness|522,527|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|History of Present Illness|522,527|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|History of Present Illness|522,533|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Finding|Sign or Symptom|History of Present Illness|528,533|false|false|false|C0003578|Apnea|apnea
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|535,545|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Finding|Functional Concept|History of Present Illness|535,545|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|History of Present Illness|535,545|false|false|false|C0460137;C1579931|Depression - motion|depression
Disorder|Disease or Syndrome|History of Present Illness|547,561|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|History of Present Illness|547,561|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Disorder|Disease or Syndrome|History of Present Illness|563,588|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid syndrome
Disorder|Disease or Syndrome|History of Present Illness|580,588|false|false|false|C0039082|Syndrome|syndrome
Anatomy|Body Location or Region|History of Present Illness|597,600|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|597,600|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|597,600|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Gene or Genome|History of Present Illness|608,611|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|612,623|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|History of Present Illness|615,623|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|History of Present Illness|615,623|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|History of Present Illness|615,623|false|false|false|C0043031|warfarin|warfarin
Finding|Idea or Concept|History of Present Illness|641,651|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|641,651|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|History of Present Illness|655,661|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|655,661|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|History of Present Illness|662,667|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|662,683|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|668,673|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|668,673|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|668,683|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Sign or Symptom|History of Present Illness|668,688|false|false|false|C0239376|Pain of lower extremities|lower extremity pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|674,683|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|History of Present Illness|674,688|false|false|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Finding|Sign or Symptom|History of Present Illness|674,688|false|false|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Attribute|Clinical Attribute|History of Present Illness|684,688|false|true|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|684,688|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|684,688|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|720,728|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|733,743|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Disorder|Neoplastic Process|History of Present Illness|758,774|false|false|false|C1176475;C1527349|Ductal Breast Carcinoma;Ductal Carcinoma|ductal carcinoma
Disorder|Neoplastic Process|History of Present Illness|765,774|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Functional Concept|History of Present Illness|778,782|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|778,789|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|783,789|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|783,789|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|783,789|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|783,789|false|false|false|C0191838|Procedures on breast|breast
Drug|Hazardous or Poisonous Substance|History of Present Illness|795,803|false|false|false|C0950580|sentinel|sentinel
Drug|Organic Chemical|History of Present Illness|795,803|false|false|false|C0950580|sentinel|sentinel
Finding|Body Substance|History of Present Illness|805,810|false|false|false|C0024202|Lymph|lymph
Finding|Finding|History of Present Illness|816,822|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|History of Present Illness|816,822|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|History of Present Illness|816,822|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|History of Present Illness|816,822|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Finding|Pathologic Function|History of Present Illness|846,854|false|false|false|C0018944|Hematoma|hematoma
Attribute|Clinical Attribute|History of Present Illness|855,861|false|false|false|C5889824||status
Finding|Idea or Concept|History of Present Illness|855,861|false|false|false|C1546481|What subject filter - Status|status
Finding|Gene or Genome|History of Present Illness|862,866|false|false|false|C3469826;C3470073|DESI1 gene;SLC35G1 gene|post
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|867,877|false|false|false|C1282573|Evacuation procedure|evacuation
Finding|Functional Concept|History of Present Illness|901,911|false|false|false|C0025664;C2700391|Methods aspects;Procedure (set of actions)|procedures
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|901,911|false|false|false|C0184661|Interventional procedure|procedures
Finding|Finding|History of Present Illness|922,928|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|922,928|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|History of Present Illness|929,934|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|929,950|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|935,940|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|935,940|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|935,950|false|false|false|C0023216|Lower Extremity|lower extremity
Finding|Sign or Symptom|History of Present Illness|935,955|false|false|false|C0239376|Pain of lower extremities|lower extremity pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|941,950|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|History of Present Illness|941,955|false|true|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Finding|Sign or Symptom|History of Present Illness|941,955|false|true|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Attribute|Clinical Attribute|History of Present Illness|951,955|false|true|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|951,955|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|951,955|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|History of Present Illness|989,992|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|989,992|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|989,992|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Functional Concept|History of Present Illness|993,1003|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|993,1003|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|993,1003|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Classification|History of Present Illness|1021,1029|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1021,1029|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1021,1029|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|History of Present Illness|1035,1050|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|History of Present Illness|1035,1050|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1035,1050|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Idea or Concept|History of Present Illness|1067,1075|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Pathologic Function|History of Present Illness|1087,1095|false|false|false|C0018944|Hematoma|hematoma
Anatomy|Body Location or Region|History of Present Illness|1109,1112|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|1109,1112|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|1109,1112|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1113,1124|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Pathologic Function|History of Present Illness|1155,1177|false|false|false|C0338380|Postoperative hematoma|postoperative hematoma
Finding|Pathologic Function|History of Present Illness|1169,1177|false|true|false|C0018944|Hematoma|hematoma
Finding|Finding|History of Present Illness|1182,1197|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|History of Present Illness|1182,1197|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1182,1197|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1225,1234|false|false|false|C0015385|Limb structure|extremity
Finding|Intellectual Product|History of Present Illness|1225,1239|false|true|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Finding|Sign or Symptom|History of Present Illness|1225,1239|false|true|false|C0030196;C4050173|Extremity Pain question;Pain in limb|extremity pain
Attribute|Clinical Attribute|History of Present Illness|1235,1239|false|true|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1235,1239|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1235,1239|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|1251,1255|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1251,1255|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1251,1255|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1263,1271|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|History of Present Illness|1297,1301|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1297,1301|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1297,1301|false|false|false|C1553498|home health encounter|home
Finding|Finding|History of Present Illness|1317,1323|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|History of Present Illness|1317,1323|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|History of Present Illness|1317,1328|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|History of Present Illness|1324,1328|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1324,1328|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1324,1328|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1353,1359|false|false|false|C0026821|Muscle Cramp|cramps
Anatomy|Body Location or Region|History of Present Illness|1371,1375|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1371,1375|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Functional Concept|History of Present Illness|1383,1388|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Attribute|Clinical Attribute|History of Present Illness|1403,1407|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1403,1407|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1403,1407|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|History of Present Illness|1442,1447|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1442,1453|false|false|false|C0230425|Structure of right thigh|right thigh
Anatomy|Body Location or Region|History of Present Illness|1448,1453|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Finding|Sign or Symptom|History of Present Illness|1477,1483|false|false|false|C0037763|Spasm|spasms
Finding|Finding|History of Present Illness|1501,1509|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1501,1509|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|History of Present Illness|1511,1519|false|false|false|C0030554|Paresthesia|tingling
Finding|Sign or Symptom|History of Present Illness|1511,1519|false|false|false|C2242996|Has tingling sensation|tingling
Finding|Sign or Symptom|History of Present Illness|1524,1532|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|History of Present Illness|1555,1576|false|false|false|C0559998|Seen in breast clinic|seen in breast clinic
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1563,1569|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|History of Present Illness|1563,1569|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|History of Present Illness|1563,1569|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1563,1569|false|false|false|C0191838|Procedures on breast|breast
Attribute|Clinical Attribute|History of Present Illness|1612,1616|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1612,1616|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1612,1616|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|1657,1667|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|History of Present Illness|1657,1667|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|History of Present Illness|1698,1707|false|false|false|C0277899|Absent pulse|pulseless
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1708,1717|false|false|false|C0015385|Limb structure|extremity
Drug|Food|History of Present Illness|1741,1747|false|false|false|C5890763||pulses
Finding|Physiologic Function|History of Present Illness|1741,1747|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|History of Present Illness|1741,1747|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|History of Present Illness|1755,1760|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1755,1765|false|false|false|C0230460|Structure of right foot|right foot
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1761,1765|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|History of Present Illness|1761,1765|false|false|false|C0555980|Foot problem|foot
Drug|Organic Chemical|History of Present Illness|1787,1794|false|false|false|C0699142|Tylenol|Tylenol
Drug|Pharmacologic Substance|History of Present Illness|1787,1794|false|false|false|C0699142|Tylenol|Tylenol
Finding|Finding|History of Present Illness|1798,1802|false|false|false|C5575035|Well (answer to question)|well
Drug|Organic Chemical|History of Present Illness|1806,1814|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|History of Present Illness|1806,1814|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|History of Present Illness|1806,1814|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Attribute|Clinical Attribute|History of Present Illness|1828,1832|false|true|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1828,1832|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1828,1832|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|History of Present Illness|1833,1839|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|1833,1839|false|false|false|C0723011|Relief brand of phenylephrine|relief
Finding|Finding|History of Present Illness|1833,1839|false|false|false|C0564405|Feeling relief|relief
Drug|Hazardous or Poisonous Substance|History of Present Illness|1868,1876|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|History of Present Illness|1868,1876|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|History of Present Illness|1868,1876|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|History of Present Illness|1889,1899|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|History of Present Illness|1889,1899|false|false|false|C0206460|enoxaparin|enoxaparin
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1900,1906|true|false|false|C0399080|Fixation of dental bridge|bridge
Finding|Functional Concept|History of Present Illness|1943,1954|false|false|false|C0332459;C4551657|Compressed structure|compression
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1943,1954|false|false|false|C0728907|Compression|compression
Procedure|Machine Activity|History of Present Illness|1943,1954|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1943,1954|false|false|false|C0565514;C1257972|Compression Therapy;Data Compression|compression
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1983,1986|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Event|Event|History of Present Illness|1993,2000|false|false|false|C1516084|Attempt|attempt
Attribute|Clinical Attribute|History of Present Illness|2016,2020|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|2016,2020|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2016,2020|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Idea or Concept|History of Present Illness|2035,2042|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2090,2093|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|History of Present Illness|2090,2093|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|History of Present Illness|2090,2093|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|History of Present Illness|2090,2093|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Functional Concept|History of Present Illness|2105,2109|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|2105,2109|false|false|false|C0582103|Medical Examination|Exam
Finding|Functional Concept|History of Present Illness|2125,2130|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2125,2146|false|false|false|C0230415|Right lower extremity|Right lower extremity
Anatomy|Body Location or Region|History of Present Illness|2131,2136|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2131,2136|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2131,2146|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2137,2146|false|false|false|C0015385|Limb structure|extremity
Drug|Food|History of Present Illness|2164,2170|false|false|false|C5890763||pulses
Finding|Physiologic Function|History of Present Illness|2164,2170|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|History of Present Illness|2164,2170|false|false|false|C0034107|Pulse taking|pulses
Drug|Food|History of Present Illness|2181,2187|false|false|false|C5890763||pulses
Finding|Physiologic Function|History of Present Illness|2181,2187|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|History of Present Illness|2181,2187|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|History of Present Illness|2196,2200|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2196,2216|false|false|false|C0230416|Left lower extremity|left lower extremity
Anatomy|Body Location or Region|History of Present Illness|2201,2206|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2201,2206|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2201,2216|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2207,2216|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|History of Present Illness|2222,2227|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2222,2243|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|2228,2233|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2228,2233|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2228,2243|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2234,2243|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|History of Present Illness|2247,2251|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2247,2251|false|false|false|C0687712|warming process|warm
Finding|Mental Process|History of Present Illness|2262,2272|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|History of Present Illness|2262,2272|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Procedure|Diagnostic Procedure|History of Present Illness|2276,2285|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|History of Present Illness|2293,2298|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|2293,2303|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|History of Present Illness|2299,2303|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2299,2303|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Mental Process|History of Present Illness|2305,2315|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Finding|Sign or Symptom|History of Present Illness|2305,2315|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|Tenderness
Procedure|Diagnostic Procedure|History of Present Illness|2320,2329|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|History of Present Illness|2337,2342|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2337,2348|false|false|false|C0230425|Structure of right thigh|right thigh
Anatomy|Body Location or Region|History of Present Illness|2343,2348|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Lab|Laboratory or Test Result|History of Present Illness|2353,2357|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Functional Concept|History of Present Illness|2373,2377|false|false|false|C0079107|chemical aspects|Chem
Procedure|Laboratory Procedure|History of Present Illness|2373,2377|false|false|false|C0201682|Chemical procedure|Chem
Finding|Idea or Concept|History of Present Illness|2378,2383|false|false|false|C0441833|Groups|panel
Anatomy|Cell Component|History of Present Illness|2416,2419|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|History of Present Illness|2416,2419|false|false|false|C0009555|Complete Blood Count|CBC
Anatomy|Cell|History of Present Illness|2421,2424|false|false|false|C0023516|Leukocytes|WBC
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2430,2433|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|History of Present Illness|2430,2433|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|History of Present Illness|2430,2433|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|History of Present Illness|2430,2433|false|false|false|C0019029|Hemoglobin concentration|Hgb
Disorder|Virus|History of Present Illness|2444,2447|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|History of Present Illness|2444,2447|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|History of Present Illness|2444,2447|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2444,2447|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Laboratory Procedure|History of Present Illness|2452,2455|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Neoplastic Process|History of Present Illness|2477,2480|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|History of Present Illness|2477,2480|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Attribute|Clinical Attribute|History of Present Illness|2487,2490|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|History of Present Illness|2487,2490|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2487,2490|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|History of Present Illness|2495,2502|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|History of Present Illness|2495,2502|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|History of Present Illness|2495,2502|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|History of Present Illness|2511,2514|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Mod
Finding|Functional Concept|History of Present Illness|2525,2533|false|false|false|C1510439|bacteria aspects|bacteria
Finding|Finding|History of Present Illness|2537,2544|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|2537,2544|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Finding|Functional Concept|History of Present Illness|2565,2575|false|false|false|C0220934|Ultrasonic|Ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2565,2575|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|Ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|2565,2575|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|Ultrasound
Finding|Functional Concept|History of Present Illness|2580,2585|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|History of Present Illness|2580,2590|false|false|false|C0489801|Posterior part of right leg|Right calf
Anatomy|Body Location or Region|History of Present Illness|2586,2590|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2586,2590|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Idea or Concept|History of Present Illness|2627,2635|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|History of Present Illness|2627,2638|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|History of Present Illness|2639,2643|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2644,2650|false|false|false|C0042449|Veins|venous
Finding|Pathologic Function|History of Present Illness|2651,2661|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|History of Present Illness|2669,2674|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2669,2690|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|History of Present Illness|2675,2680|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2675,2680|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2675,2690|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2675,2696|false|false|false|C0226813;C4266545|Lower extremity>Lower extremity veins;Structure of vein of lower extremity|lower extremity veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2681,2690|false|false|false|C0015385|Limb structure|extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2681,2696|false|false|false|C0730267|Venous structure of limb|extremity veins
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2691,2696|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2691,2696|false|true|false|C0398102|Procedure on vein|veins
Attribute|Clinical Attribute|History of Present Illness|2699,2717|false|false|false|C1524365||CT Lower Extremity
Anatomy|Body Location or Region|History of Present Illness|2702,2707|false|false|false|C1548802|Body Site Modifier - Lower|Lower
Event|Activity|History of Present Illness|2702,2707|false|false|false|C2003888|Lower (action)|Lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2702,2717|false|false|false|C0023216|Lower Extremity|Lower Extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2708,2717|false|false|false|C0015385|Limb structure|Extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2708,2723|false|false|false|C0947119|Extremity Right|Extremity Right
Finding|Functional Concept|History of Present Illness|2718,2723|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Drug|Indicator, Reagent, or Diagnostic Aid|History of Present Illness|2741,2749|false|false|false|C0009924|Contrast Media|contrast
Finding|Functional Concept|History of Present Illness|2769,2774|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|History of Present Illness|2769,2779|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|History of Present Illness|2775,2779|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2775,2779|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Location or Region|History of Present Illness|2791,2797|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2791,2797|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2812,2816|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|History of Present Illness|2812,2816|false|false|false|C0555980|Foot problem|foot
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2822,2827|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2822,2827|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|History of Present Illness|2835,2840|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|2835,2840|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2835,2850|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2841,2850|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|History of Present Illness|2920,2926|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Functional Concept|History of Present Illness|2927,2937|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2927,2937|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|2927,2937|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Conceptual Entity|History of Present Illness|2971,2981|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|History of Present Illness|2971,2981|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|History of Present Illness|2971,2981|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|History of Present Illness|2971,2981|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2993,3001|false|false|false|C4083049|Muscle (organ)|muscular
Disorder|Anatomical Abnormality|History of Present Illness|2993,3013|true|false|false|C4021745|Abnormality of the musculature|muscular abnormality
Disorder|Congenital Abnormality|History of Present Illness|3002,3013|true|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|History of Present Illness|3002,3013|true|false|false|C1704258|Abnormality|abnormality
Drug|Organic Chemical|History of Present Illness|3051,3059|false|false|false|C0026549|morphine|Morphine
Drug|Pharmacologic Substance|History of Present Illness|3051,3059|false|false|false|C0026549|morphine|Morphine
Disorder|Disease or Syndrome|History of Present Illness|3067,3071|false|false|false|C1970472|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED|APAP
Drug|Organic Chemical|History of Present Illness|3067,3071|false|false|false|C0000970|acetaminophen|APAP
Drug|Pharmacologic Substance|History of Present Illness|3067,3071|false|false|false|C0000970|acetaminophen|APAP
Drug|Organic Chemical|History of Present Illness|3084,3092|false|false|false|C0728755|Dilaudid|Dilaudid
Drug|Pharmacologic Substance|History of Present Illness|3084,3092|false|false|false|C0728755|Dilaudid|Dilaudid
Drug|Hazardous or Poisonous Substance|History of Present Illness|3114,3122|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|History of Present Illness|3114,3122|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|History of Present Illness|3114,3122|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|History of Present Illness|3129,3141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|History of Present Illness|3129,3141|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|History of Present Illness|3147,3157|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|History of Present Illness|3147,3157|false|false|false|C0028978|omeprazole|Omeprazole
Finding|Finding|History of Present Illness|3164,3171|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|History of Present Illness|3164,3171|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|History of Present Illness|3164,3171|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3164,3171|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3197,3205|false|false|false|C0005847|Blood Vessel|vascular
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3197,3213|false|false|false|C0042381|Vascular Surgical Procedures|vascular surgery
Finding|Finding|History of Present Illness|3206,3213|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|3206,3213|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|3206,3213|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3206,3213|false|false|false|C0543467|Operative Surgical Procedures|surgery
Procedure|Health Care Activity|History of Present Illness|3214,3221|false|false|false|C0009818|Consultation|consult
Finding|Finding|History of Present Illness|3226,3234|false|false|false|C0332149|Possible|possible
Anatomy|Body Location or Region|History of Present Illness|3235,3238|false|false|false|C5239664|area DVT|dvt
Attribute|Clinical Attribute|History of Present Illness|3235,3238|false|true|false|C2926618||dvt
Disorder|Disease or Syndrome|History of Present Illness|3235,3238|false|true|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|dvt
Finding|Conceptual Entity|History of Present Illness|3244,3251|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3244,3251|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|3244,3251|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|3244,3254|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3264,3268|false|false|false|C0042449|Veins|vein
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3264,3278|false|false|false|C0149807|Stripping of vein|vein stripping
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3269,3278|false|false|false|C0185047|Stripping (procedure)|stripping
Finding|Functional Concept|History of Present Illness|3279,3289|false|false|false|C0025664;C2700391|Methods aspects;Procedure (set of actions)|procedures
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3279,3289|false|false|false|C0184661|Interventional procedure|procedures
Disorder|Disease or Syndrome|History of Present Illness|3294,3298|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Procedure|Health Care Activity|History of Present Illness|3315,3324|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Pharmacologic Substance|History of Present Illness|3328,3336|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Attribute|Clinical Attribute|History of Present Illness|3341,3345|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3341,3345|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3341,3345|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|3341,3353|false|false|false|C5548091|Demonstrates adequate pain control|pain control
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3341,3353|false|false|false|C0002766;C1304888|Pain control;Pain management (procedure)|pain control
Drug|Organic Chemical|History of Present Illness|3346,3353|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|History of Present Illness|3346,3353|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|History of Present Illness|3346,3353|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Finding|Conceptual Entity|History of Present Illness|3346,3353|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|History of Present Illness|3346,3353|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|History of Present Illness|3346,3353|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3358,3366|false|false|false|C0005847|Blood Vessel|Vascular
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3358,3374|false|false|false|C0042381|Vascular Surgical Procedures|Vascular surgery
Finding|Finding|History of Present Illness|3367,3374|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|3367,3374|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|3367,3374|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3367,3374|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Idea or Concept|History of Present Illness|3402,3407|true|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3408,3416|false|false|false|C0005847|Blood Vessel|vascular
Finding|Conceptual Entity|History of Present Illness|3417,3425|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Finding|Functional Concept|History of Present Illness|3417,3425|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|etiology
Attribute|Clinical Attribute|History of Present Illness|3434,3438|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3434,3438|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3434,3438|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|History of Present Illness|3459,3467|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|3459,3467|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|3459,3467|false|false|false|C4706767|Transfer (immobility management)|transfer
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|3508,3511|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|History of Present Illness|3508,3511|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|History of Present Illness|3508,3511|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|History of Present Illness|3508,3511|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Event|Activity|History of Present Illness|3527,3534|false|false|false|C1706079||arrival
Finding|Functional Concept|History of Present Illness|3527,3534|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|3542,3547|false|false|false|C3714591|Floor (anatomic)|floor
Finding|Body Substance|History of Present Illness|3553,3560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|3553,3560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|3553,3560|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|History of Present Illness|3573,3577|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3573,3577|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3573,3577|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|3614,3618|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3614,3618|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3614,3618|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|3637,3641|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3637,3641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3637,3641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|History of Present Illness|3666,3670|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Functional Concept|History of Present Illness|3674,3684|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|History of Present Illness|3674,3684|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|History of Present Illness|3674,3684|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Location or Region|History of Present Illness|3695,3698|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|3695,3698|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|3695,3698|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Finding|History of Present Illness|3707,3711|false|false|false|C1299581|Able (qualifier value)|able
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3725,3729|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Attribute|Clinical Attribute|History of Present Illness|3738,3742|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3738,3742|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3738,3742|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3760,3763|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Intellectual Product|History of Present Illness|3788,3792|false|false|false|C1706124|Terminology Kind|kind
Attribute|Clinical Attribute|History of Present Illness|3796,3800|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3796,3800|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3796,3800|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3823,3827|false|false|false|C0042449|Veins|vein
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3823,3837|false|false|false|C0149807|Stripping of vein|vein stripping
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|3828,3837|false|false|false|C0185047|Stripping (procedure)|stripping
Attribute|Clinical Attribute|History of Present Illness|3864,3867|false|false|false|C1114365||age
Drug|Biologically Active Substance|History of Present Illness|3864,3867|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|History of Present Illness|3864,3867|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Location or Region|History of Present Illness|3884,3889|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|3884,3889|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|3884,3894|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|3884,3894|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|3890,3894|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|3890,3894|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|3890,3894|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Body Substance|History of Present Illness|3911,3917|false|false|false|C0225386|Breath|breath
Finding|Daily or Recreational Activity|History of Present Illness|3941,3947|true|false|false|C0040802|travel|travel
Procedure|Health Care Activity|History of Present Illness|3941,3947|true|false|false|C1555670|travel charge|travel
Disorder|Injury or Poisoning|History of Present Illness|3951,3957|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|History of Present Illness|3951,3957|true|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|3965,3968|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|Past Medical History|3996,4008|false|false|false|C0242339|Dyslipidemias|Dyslipidemia
Disorder|Disease or Syndrome|Past Medical History|4011,4025|false|false|false|C0042345|Varicosity|Varicose veins
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4020,4025|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4020,4025|false|false|false|C0398102|Procedure on vein|veins
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4036,4044|false|false|false|C0023690|Ligation|ligation
Disorder|Disease or Syndrome|Past Medical History|4047,4051|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|4047,4051|false|false|false|C1647218|COPD pharmacologic substance|COPD
Finding|Gene or Genome|Past Medical History|4047,4051|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|4054,4057|false|false|false|C0520679|Sleep Apnea, Obstructive|OSA
Drug|Amino Acid, Peptide, or Protein|Past Medical History|4054,4057|false|false|false|C0764906|OSA protein, Drosophila|OSA
Drug|Biologically Active Substance|Past Medical History|4054,4057|false|false|false|C0764906|OSA protein, Drosophila|OSA
Finding|Gene or Genome|Past Medical History|4060,4064|false|false|false|C1424863|CENPJ gene|CPap
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4060,4064|false|false|false|C0199451|Continuous Positive Airway Pressure|CPap
Finding|Finding|Past Medical History|4068,4078|false|false|false|C2169609|recent upper respiratory infection|recent URI
Disorder|Disease or Syndrome|Past Medical History|4075,4078|false|false|false|C0041912|Upper Respiratory Infections|URI
Finding|Gene or Genome|Past Medical History|4075,4078|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|Past Medical History|4075,4078|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Drug|Antibiotic|Past Medical History|4099,4108|false|false|false|C0678143|Zithromax|Zithromax
Drug|Organic Chemical|Past Medical History|4099,4108|false|false|false|C0678143|Zithromax|Zithromax
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4122,4125|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|Past Medical History|4122,4125|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|Past Medical History|4122,4125|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Drug|Amino Acid, Peptide, or Protein|Past Medical History|4134,4159|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Drug|Immunologic Factor|Past Medical History|4134,4159|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Finding|Finding|Past Medical History|4134,4159|false|false|false|C4019436|Antiphospholipid antibody positivity|antiphospholipid antibody
Disorder|Disease or Syndrome|Past Medical History|4134,4168|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid antibody syndrome
Anatomy|Cell Component|Past Medical History|4151,4159|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Past Medical History|4151,4159|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Past Medical History|4151,4159|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Past Medical History|4151,4159|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Past Medical History|4151,4159|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Past Medical History|4160,4168|false|false|false|C0039082|Syndrome|syndrome
Finding|Finding|Past Medical History|4183,4198|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Past Medical History|4183,4198|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4183,4198|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Classification|Past Medical History|4213,4216|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1C
Procedure|Laboratory Procedure|Past Medical History|4213,4216|false|false|false|C0474680|Hemoglobin A1c measurement|A1C
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4230,4238|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|Past Medical History|4230,4247|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Finding|Pathologic Function|Past Medical History|4239,4247|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Finding|Past Medical History|4270,4279|false|false|false|C0442739||unchanged
Disorder|Disease or Syndrome|Past Medical History|4283,4287|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Disorder|Disease or Syndrome|Past Medical History|4290,4304|false|false|false|C1510475|Diverticulosis|diverticulosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4311,4316|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Past Medical History|4311,4316|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Past Medical History|4311,4316|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Past Medical History|4311,4316|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Anatomical Abnormality|Past Medical History|4311,4323|false|false|false|C0009376|Colonic Polyps|colon polyps
Disorder|Anatomical Abnormality|Past Medical History|4317,4323|false|false|false|C0032584|polyps|polyps
Finding|Intellectual Product|Past Medical History|4317,4323|false|false|false|C1546747||polyps
Disorder|Mental or Behavioral Dysfunction|Past Medical History|4326,4336|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Finding|Functional Concept|Past Medical History|4326,4336|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|4326,4336|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Functional Concept|Past Medical History|4343,4348|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Cell|Past Medical History|4349,4352|false|false|false|C3890599|Circulating Melanoma Cell|CMC
Disorder|Congenital Abnormality|Past Medical History|4349,4352|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Disorder|Disease or Syndrome|Past Medical History|4349,4352|false|false|false|C0006845;C0340803|Candidiasis, Chronic Mucocutaneous;Capillary malformation (disorder)|CMC
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4349,4352|false|false|false|C0065772|MCC protocol|CMC
Anatomy|Body Space or Junction|Past Medical History|4353,4358|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Anatomy|Body System|Past Medical History|4353,4358|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|joint
Finding|Finding|Past Medical History|4353,4358|false|false|false|C0575044|Joint problem|joint
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4353,4371|false|false|false|C0003893|Arthroplasty|joint arthroplasty
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4359,4371|false|false|false|C0003893;C0700235;C5887062|Arthroplasty;Reconstruction of joint;Temporomandibular joint arthroplasty by dentist|arthroplasty
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4378,4390|false|false|false|C0085515|Rotator Cuff|rotator cuff
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4378,4397|false|false|false|C0186666|Repair of musculotendinous cuff of shoulder|rotator cuff repair
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4386,4390|false|false|false|C1550244|Cuff - body part|cuff
Finding|Pathologic Function|Past Medical History|4386,4390|false|false|false|C3668885|Cuffing (morphologic abnormality)|cuff
Finding|Functional Concept|Past Medical History|4391,4397|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Past Medical History|4391,4397|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Past Medical History|4391,4397|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4391,4397|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4400,4408|false|false|false|C0015252;C0728940|Excision;removal technique|excision
Finding|Functional Concept|Past Medical History|4409,4414|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4419,4424|false|false|false|C0582802|Digit structure|digit
Finding|Gene or Genome|Past Medical History|4419,4424|false|false|false|C4761764|GSC-DT gene|digit
Finding|Finding|Past Medical History|4425,4429|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Past Medical History|4425,4429|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Past Medical History|4425,4429|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Body Substance|Past Medical History|4438,4443|false|false|false|C0006736|Calculi|stone
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4446,4456|false|false|false|C0030274|Pancreas|pancreatic
Drug|Amino Acid, Peptide, or Protein|Past Medical History|4446,4456|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Hormone|Past Medical History|4446,4456|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Drug|Pharmacologic Substance|Past Medical History|4446,4456|false|false|false|C0030292|Pancreatic Hormones|pancreatic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4446,4461|false|false|false|C0030288;C4482304|Abdomen>Pancreatic duct;Pancreatic duct|pancreatic duct
Disorder|Neoplastic Process|Past Medical History|4446,4461|false|false|false|C0153461|Malignant neoplasm of pancreatic duct|pancreatic duct
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|4457,4461|false|false|false|C0687028;C1550227|Duct (organ) structure;canal [body parts]|duct
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4462,4473|false|false|false|C1280903|Exploration procedure|exploration
Finding|Finding|Past Medical History|4482,4494|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4482,4494|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|4497,4510|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Finding|Idea or Concept|Family Medical History|4551,4557|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4566,4573|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|4566,4580|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|4574,4580|false|false|false|C0006826|Malignant Neoplasms|CANCER
Attribute|Clinical Attribute|Family Medical History|4574,4583|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Family Medical History|4584,4587|false|false|false|C1114365||age
Drug|Biologically Active Substance|Family Medical History|4584,4587|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Family Medical History|4584,4587|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|Family Medical History|4593,4599|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|4593,4599|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4608,4613|false|false|false|C0006104;C4266577|Brain;Head>Brain|BRAIN
Disorder|Disease or Syndrome|Family Medical History|4608,4613|false|false|false|C0006111|Brain Diseases|BRAIN
Disorder|Neoplastic Process|Family Medical History|4608,4620|false|false|false|C0006118;C0153633|Brain Neoplasms;Malignant neoplasm of brain|BRAIN CANCER
Disorder|Neoplastic Process|Family Medical History|4614,4620|false|false|false|C0006826|Malignant Neoplasms|CANCER
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4622,4625|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Drug|Enzyme|Family Medical History|4622,4625|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Drug|Inorganic Chemical|Family Medical History|4622,4625|false|false|false|C0031653;C3815181|PHOSPHOGLUCOMUTASE;Platinum-Group Metal|PGM
Finding|Molecular Function|Family Medical History|4622,4625|false|false|false|C1150365|phosphoglycerate mutase activity|PGM
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4626,4633|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|4626,4640|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|4634,4640|false|false|false|C0006826|Malignant Neoplasms|CANCER
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4647,4654|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Family Medical History|4647,4661|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Family Medical History|4655,4661|false|false|false|C0006826|Malignant Neoplasms|CANCER
Disorder|Neoplastic Process|Family Medical History|4690,4708|false|false|false|C0007103;C0476089|Endometrial Carcinoma;Malignant neoplasm of endometrium|ENDOMETRIAL CANCER
Disorder|Neoplastic Process|Family Medical History|4702,4708|false|false|false|C0006826|Malignant Neoplasms|CANCER
Drug|Amino Acid, Peptide, or Protein|Family Medical History|4710,4713|false|false|false|C1366394;C3712803;C3887684|IGF1 protein, human;Kit Ligand, human;STAT5A protein, human|MGF
Drug|Biologically Active Substance|Family Medical History|4710,4713|false|false|false|C1366394;C3712803;C3887684|IGF1 protein, human;Kit Ligand, human;STAT5A protein, human|MGF
Finding|Gene or Genome|Family Medical History|4710,4713|false|false|false|C1335875;C1366480;C1704887;C1705050|KITLG gene;KITLG wt Allele;STAT5A gene;STAT5A wt Allele|MGF
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4714,4722|false|false|false|C0033572;C4266527|Prostate;Structure of prostate (body structure)|PROSTATE
Disorder|Disease or Syndrome|Family Medical History|4714,4722|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|PROSTATE
Disorder|Neoplastic Process|Family Medical History|4714,4722|false|false|false|C0033575;C0154009;C0154088;C0496923|Benign neoplasm of prostate;Carcinoma in situ of prostate;Neoplasm of uncertain or unknown behavior of prostate;Prostatic Diseases|PROSTATE
Disorder|Neoplastic Process|Family Medical History|4714,4729|false|false|false|C0376358;C0600139|Malignant neoplasm of prostate;Prostate carcinoma|PROSTATE CANCER
Disorder|Neoplastic Process|Family Medical History|4723,4729|false|false|false|C0006826|Malignant Neoplasms|CANCER
Finding|Conceptual Entity|Family Medical History|4731,4738|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|4731,4738|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4747,4753|false|false|false|C0022646;C0227665|Both kidneys;Kidney|KIDNEY
Disorder|Neoplastic Process|Family Medical History|4747,4753|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|KIDNEY
Finding|Sign or Symptom|Family Medical History|4747,4753|false|false|false|C0812426|Kidney problem|KIDNEY
Procedure|Diagnostic Procedure|Family Medical History|4747,4753|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Procedure|Therapeutic or Preventive Procedure|Family Medical History|4747,4753|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|KIDNEY
Disorder|Neoplastic Process|Family Medical History|4747,4760|false|false|false|C0740457;C1378703|Malignant neoplasm of kidney;Renal carcinoma|KIDNEY CANCER
Disorder|Neoplastic Process|Family Medical History|4754,4760|false|false|false|C0006826|Malignant Neoplasms|CANCER
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4763,4768|false|false|false|C0022646|Kidney|RENAL
Disorder|Disease or Syndrome|Family Medical History|4763,4768|false|false|false|C0042075|Urologic Diseases|RENAL
Disorder|Disease or Syndrome|Family Medical History|4763,4776|false|false|false|C0035078|Kidney Failure|RENAL FAILURE
Finding|Functional Concept|Family Medical History|4769,4776|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Family Medical History|4769,4776|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Family Medical History|4769,4776|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|4790,4795|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Family Medical History|4790,4795|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|Family Medical History|4790,4795|false|false|false|C0795691|HEART PROBLEM|HEART
Finding|Functional Concept|Family Medical History|4798,4805|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Family Medical History|4798,4805|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Family Medical History|4798,4805|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Disorder|Disease or Syndrome|Family Medical History|4808,4816|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|DIABETES
Disorder|Disease or Syndrome|Family Medical History|4808,4825|false|false|false|C0011849|Diabetes Mellitus|DIABETES MELLITUS
Drug|Hazardous or Poisonous Substance|Family Medical History|4828,4835|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Immunologic Factor|Family Medical History|4828,4835|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Organic Chemical|Family Medical History|4828,4835|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Drug|Pharmacologic Substance|Family Medical History|4828,4835|false|false|false|C0040329;C2701271|Tobacco;tobacco leaf allergenic extract|TOBACCO
Disorder|Mental or Behavioral Dysfunction|Family Medical History|4828,4841|false|false|false|C0040336|Tobacco Use Disorder|TOBACCO ABUSE
Disorder|Mental or Behavioral Dysfunction|Family Medical History|4836,4841|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Family Medical History|4836,4841|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Family Medical History|4836,4841|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Finding|Conceptual Entity|Substance Abuse Treatment|4859,4865|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|Sister
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|4874,4881|false|false|false|C0205065|Ovarian|OVARIAN
Disorder|Neoplastic Process|Substance Abuse Treatment|4874,4888|false|false|false|C0919267;C1140680|Malignant neoplasm of ovary;ovarian neoplasm|OVARIAN CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|4882,4888|false|false|false|C0006826|Malignant Neoplasms|CANCER
Attribute|Clinical Attribute|Substance Abuse Treatment|4882,4891|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Substance Abuse Treatment|4892,4895|false|false|false|C1114365||age
Drug|Biologically Active Substance|Substance Abuse Treatment|4892,4895|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Substance Abuse Treatment|4892,4895|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|Substance Abuse Treatment|4901,4908|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Substance Abuse Treatment|4901,4908|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Anatomy|Body Location or Region|Substance Abuse Treatment|4913,4919|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|THROAT
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|4913,4919|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|THROAT
Drug|Pharmacologic Substance|Substance Abuse Treatment|4913,4919|false|false|false|C1950455|Throat Homeopathic Medication|THROAT
Finding|Body Substance|Substance Abuse Treatment|4913,4919|false|false|false|C1547926;C1550663|Specimen Type - Throat|THROAT
Finding|Intellectual Product|Substance Abuse Treatment|4913,4919|false|false|false|C1547926;C1550663|Specimen Type - Throat|THROAT
Disorder|Neoplastic Process|Substance Abuse Treatment|4913,4926|false|false|false|C0740339|Throat cancer|THROAT CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|4920,4926|false|false|false|C0006826|Malignant Neoplasms|CANCER
Attribute|Clinical Attribute|Substance Abuse Treatment|4920,4929|false|false|false|C3533909||CANCER dx
Attribute|Clinical Attribute|Substance Abuse Treatment|4930,4933|false|false|false|C1114365||age
Drug|Biologically Active Substance|Substance Abuse Treatment|4930,4933|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Substance Abuse Treatment|4930,4933|false|false|false|C0162574|Glycation End Products, Advanced|age
Finding|Conceptual Entity|Substance Abuse Treatment|4954,4960|false|false|false|C1546515;C1704647|Relationship - Sister;Sister - courtesy title|Sister
Drug|Amino Acid, Peptide, or Protein|Substance Abuse Treatment|4961,4966|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|Substance Abuse Treatment|4961,4966|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Finding|Gene or Genome|Substance Abuse Treatment|4961,4966|false|false|false|C0376571|BRCA1 gene|BRCA1
Disorder|Cell or Molecular Dysfunction|Substance Abuse Treatment|4961,4975|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 MUTATION
Disorder|Cell or Molecular Dysfunction|Substance Abuse Treatment|4967,4975|false|false|false|C1705285|Mutation Abnormality|MUTATION
Finding|Genetic Function|Substance Abuse Treatment|4967,4975|false|false|false|C0026882|Mutation|MUTATION
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|4977,4983|false|false|false|C0006141|Breast|BREAST
Disorder|Neoplastic Process|Substance Abuse Treatment|4977,4983|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|BREAST
Finding|Finding|Substance Abuse Treatment|4977,4983|false|false|false|C0567499|Breast problem|BREAST
Procedure|Therapeutic or Preventive Procedure|Substance Abuse Treatment|4977,4983|false|false|false|C0191838|Procedures on breast|BREAST
Disorder|Neoplastic Process|Substance Abuse Treatment|4977,4990|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|BREAST CANCER
Disorder|Neoplastic Process|Substance Abuse Treatment|4984,4990|false|false|false|C0006826|Malignant Neoplasms|CANCER
Finding|Finding|Substance Abuse Treatment|5012,5020|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Idea or Concept|Substance Abuse Treatment|5012,5020|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|ABNORMAL
Finding|Finding|Substance Abuse Treatment|5012,5030|false|false|false|C0476427|Abnormal cervical smear|ABNORMAL PAP SMEAR
Anatomy|Body Part, Organ, or Organ Component|Substance Abuse Treatment|5021,5024|false|false|false|C3496568|pars anterior of the paramedian lobule|PAP
Drug|Amino Acid, Peptide, or Protein|Substance Abuse Treatment|5021,5024|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Drug|Enzyme|Substance Abuse Treatment|5021,5024|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Drug|Immunologic Factor|Substance Abuse Treatment|5021,5024|false|false|false|C0760170;C1740167|ACPP protein, human;alpha 2-plasmin inhibitor-plasmin complex|PAP
Finding|Finding|Substance Abuse Treatment|5021,5024|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Finding|Gene or Genome|Substance Abuse Treatment|5021,5024|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Finding|Molecular Function|Substance Abuse Treatment|5021,5024|false|false|false|C0428642;C1367456;C1413944;C1413945;C1418410;C1422804;C1423108;C1424700;C1538823;C1705529;C1705530;C1705531;C1863340;C2266415;C3538851;C3889402|ACP3 gene;ACP3 wt Allele;ASAP1 gene;ASAP1 wt Allele;ASAP2 gene;MRPS30 gene;PAPOLA gene;PAPOLA wt Allele;PDAP1 gene;PITUITARY ADENOMA PREDISPOSITION;Pulmonary artery pressure;REG3A gene;REG3A wt Allele;TUSC2 gene;TUSC2 wt Allele|PAP
Procedure|Diagnostic Procedure|Substance Abuse Treatment|5021,5030|false|false|false|C0079104;C3541459|Pap smear;Papanicolaou Test|PAP SMEAR
Procedure|Laboratory Procedure|Substance Abuse Treatment|5021,5030|false|false|false|C0079104;C3541459|Pap smear;Papanicolaou Test|PAP SMEAR
Event|Activity|Substance Abuse Treatment|5025,5030|false|false|false|C1947932|Smear - instruction imperative|SMEAR
Finding|Functional Concept|Substance Abuse Treatment|5025,5030|false|false|false|C3872789|Smearing technique|SMEAR
Procedure|Diagnostic Procedure|Substance Abuse Treatment|5025,5030|false|false|false|C0444186|Smear test|SMEAR
Finding|Gene or Genome|Substance Abuse Treatment|5053,5056|false|false|false|C1420310|SON gene|Son
Attribute|Clinical Attribute|Substance Abuse Treatment|5066,5075|false|false|false|C5889933||SUBSTANCE
Drug|Substance|Substance Abuse Treatment|5066,5075|false|false|false|C0439861|Substance|SUBSTANCE
Finding|Intellectual Product|Substance Abuse Treatment|5066,5075|false|false|false|C5887067|administrative information regarding test substance|SUBSTANCE
Disorder|Mental or Behavioral Dysfunction|Substance Abuse Treatment|5066,5081|false|false|false|C0740858;C5967394|Harmful pattern of substance use;Substance Abuse Problems|SUBSTANCE ABUSE
Disorder|Mental or Behavioral Dysfunction|Substance Abuse Treatment|5076,5081|false|false|false|C0013146|Drug abuse|ABUSE
Event|Event|Substance Abuse Treatment|5076,5081|false|false|false|C1546935|Abuse|ABUSE
Finding|Finding|Substance Abuse Treatment|5076,5081|false|false|false|C0562381|Victim of abuse (finding)|ABUSE
Disorder|Injury or Poisoning|Substance Abuse Treatment|5088,5094|false|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|Substance Abuse Treatment|5088,5094|false|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|Substance Abuse Treatment|5088,5094|false|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|Substance Abuse Treatment|5088,5094|false|false|false|C0011892|heroin|heroin
Disorder|Injury or Poisoning|Substance Abuse Treatment|5088,5103|false|false|false|C0572070|Heroin overdose|heroin overdose
Disorder|Injury or Poisoning|Substance Abuse Treatment|5095,5103|false|false|false|C0029944|Drug Overdose|overdose
Finding|Finding|Substance Abuse Treatment|5095,5103|false|false|false|C1546941;C4018909|Event Qualification - Overdose;Overdose|overdose
Finding|Idea or Concept|Substance Abuse Treatment|5095,5103|false|false|false|C1546941;C4018909|Event Qualification - Overdose;Overdose|overdose
Procedure|Health Care Activity|General Exam|5129,5138|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|General Exam|5139,5143|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5139,5143|false|false|false|C0582103|Medical Examination|EXAM
Drug|Amino Acid, Peptide, or Protein|General Exam|5208,5211|false|false|false|C2744672|SAT1 protein, human|Sat
Drug|Enzyme|General Exam|5208,5211|false|false|false|C2744672|SAT1 protein, human|Sat
Finding|Gene or Genome|General Exam|5208,5211|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Intellectual Product|General Exam|5208,5211|false|false|false|C0871290;C1705827;C1822614|College Entrance Examination Board Scholastic Aptitude Test;SAT1 gene;SAT1 wt Allele|Sat
Finding|Classification|General Exam|5219,5226|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|5219,5226|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|General Exam|5228,5233|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|5228,5233|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|5228,5233|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|5228,5233|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|5228,5233|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|5228,5233|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|5248,5253|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|5254,5262|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|5254,5262|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|5265,5270|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|5272,5275|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|5272,5275|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|5277,5287|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|5288,5293|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|General Exam|5301,5306|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|General Exam|5308,5312|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|5308,5312|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|5308,5312|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|General Exam|5308,5319|false|false|false|C2230237|Supple neck|neck supple
Finding|Functional Concept|General Exam|5313,5319|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|5321,5324|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|General Exam|5338,5343|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|5338,5343|false|false|false|C0741025|Chest problem|Chest
Anatomy|Body Part, Organ, or Organ Component|General Exam|5347,5353|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|5347,5353|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|General Exam|5347,5353|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|5347,5353|false|false|false|C0191838|Procedures on breast|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|5354,5363|false|false|false|C0184898|Surgical incisions|incisions
Finding|Finding|General Exam|5364,5368|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|General Exam|5369,5375|false|false|false|C0205249|Healed|healed
Anatomy|Body Location or Region|General Exam|5383,5389|false|false|false|C0004454|Axilla|axilla
Procedure|Health Care Activity|General Exam|5390,5398|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|General Exam|5390,5398|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Drug|Substance|General Exam|5399,5404|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|5399,5404|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|General Exam|5399,5412|false|false|false|C0411815|Removal of drain|drain removal
Event|Activity|General Exam|5405,5412|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|General Exam|5405,5412|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Activity|General Exam|5426,5430|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|5426,5430|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|5435,5441|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|5435,5441|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|General Exam|5462,5469|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|5470,5475|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|5477,5482|false|false|false|C1550016|Remote control command - Clear|Clear
Procedure|Diagnostic Procedure|General Exam|5486,5498|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|General Exam|5515,5522|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|General Exam|5526,5534|true|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Anatomy|Body Location or Region|General Exam|5535,5542|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|5535,5542|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|5535,5542|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|5544,5548|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|5577,5582|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|5577,5589|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|5583,5589|false|false|false|C0037709||sounds
Finding|Finding|General Exam|5590,5597|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|5590,5597|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Congenital Abnormality|General Exam|5598,5601|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|5598,5601|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|5603,5607|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|5603,5607|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|5609,5613|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|General Exam|5624,5629|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5624,5645|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|General Exam|5630,5635|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5630,5635|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5630,5645|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|5636,5645|false|false|false|C0015385|Limb structure|extremity
Procedure|Diagnostic Procedure|General Exam|5659,5668|false|false|false|C0030247|Palpation|palpation
Finding|Organism Function|General Exam|5673,5681|false|false|false|C0026649|Movement|movement
Attribute|Clinical Attribute|General Exam|5693,5697|false|false|false|C2598155||pain
Finding|Functional Concept|General Exam|5693,5697|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|5693,5697|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|General Exam|5699,5707|false|false|false|C0013604;C0038999|Edema;Swelling|Swelling
Finding|Pathologic Function|General Exam|5699,5707|false|false|false|C0013604;C0038999|Edema;Swelling|Swelling
Drug|Food|General Exam|5738,5744|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|5738,5744|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|5738,5744|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body System|General Exam|5758,5762|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|5758,5762|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|5758,5762|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|5758,5762|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|5758,5762|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Finding|General Exam|5764,5768|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|5764,5768|false|false|false|C0687712|warming process|Warm
Disorder|Disease or Syndrome|General Exam|5775,5789|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|5784,5789|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|5784,5789|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|5799,5804|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5799,5804|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|5799,5816|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|5805,5816|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Finding|General Exam|5835,5841|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Idea or Concept|General Exam|5858,5866|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|General Exam|5871,5880|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|5871,5880|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|5871,5880|false|false|false|C2229507|sensory exam|sensation
Finding|Conceptual Entity|General Exam|5886,5895|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|5886,5895|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Body Substance|General Exam|5909,5918|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5909,5918|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5909,5918|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5909,5918|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|General Exam|5919,5923|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5919,5923|false|false|false|C0582103|Medical Examination|EXAM
Finding|Gene or Genome|General Exam|5950,5954|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|5950,5954|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Finding|Finding|General Exam|6048,6056|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|6048,6056|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|6048,6056|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|6048,6056|false|false|false|C0011209|Obstetric Delivery|delivery
Finding|Classification|General Exam|6066,6073|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|6066,6073|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|General Exam|6075,6080|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|6075,6080|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|6075,6080|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|6075,6080|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|6075,6080|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|6075,6080|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|6095,6100|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|6101,6109|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|6101,6109|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|6112,6117|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|6119,6122|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|6119,6122|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|6124,6134|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|6135,6140|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|General Exam|6148,6153|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|General Exam|6155,6159|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|6155,6159|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|6155,6159|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Finding|General Exam|6155,6166|false|false|false|C2230237|Supple neck|neck supple
Finding|Functional Concept|General Exam|6160,6166|false|false|false|C0332254|Supple|supple
Finding|Finding|General Exam|6168,6171|false|false|false|C0428897|Jugular venous pressure|JVP
Anatomy|Body Location or Region|General Exam|6185,6190|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|General Exam|6185,6190|false|false|false|C0741025|Chest problem|Chest
Anatomy|Body Part, Organ, or Organ Component|General Exam|6194,6200|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|General Exam|6194,6200|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|General Exam|6194,6200|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|6194,6200|false|false|false|C0191838|Procedures on breast|breast
Procedure|Therapeutic or Preventive Procedure|General Exam|6201,6210|false|false|false|C0184898|Surgical incisions|incisions
Finding|Finding|General Exam|6211,6215|false|false|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|General Exam|6216,6222|false|false|false|C0205249|Healed|healed
Anatomy|Body Location or Region|General Exam|6230,6236|false|false|false|C0004454|Axilla|axilla
Procedure|Health Care Activity|General Exam|6237,6245|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Procedure|Therapeutic or Preventive Procedure|General Exam|6237,6245|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|surgical
Drug|Substance|General Exam|6246,6251|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|6246,6251|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|General Exam|6246,6259|false|false|false|C0411815|Removal of drain|drain removal
Event|Activity|General Exam|6252,6259|false|false|false|C1883720|Removing (action)|removal
Procedure|Therapeutic or Preventive Procedure|General Exam|6252,6259|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Finding|Finding|General Exam|6273,6280|true|false|false|C0018808|Heart murmur|murmurs
Anatomy|Body Part, Organ, or Organ Component|General Exam|6281,6286|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|6288,6293|false|false|false|C1550016|Remote control command - Clear|Clear
Anatomy|Body Location or Region|General Exam|6294,6301|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|6294,6301|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|6294,6301|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|6303,6307|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|6336,6341|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|6336,6348|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|6342,6348|false|false|false|C0037709||sounds
Finding|Finding|General Exam|6349,6356|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|6349,6356|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Congenital Abnormality|General Exam|6357,6360|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|6357,6360|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|6362,6366|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|6362,6366|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|6368,6372|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|6397,6405|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|6397,6405|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Procedure|Diagnostic Procedure|General Exam|6427,6436|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|General Exam|6447,6452|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|6453,6471|false|false|false|C0224813|Structure of trochanteric bursa|trochanteric bursa
Anatomy|Body Part, Organ, or Organ Component|General Exam|6466,6471|false|false|false|C0006441|Synovial bursa|bursa
Procedure|Diagnostic Procedure|General Exam|6496,6505|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|General Exam|6516,6521|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|6516,6527|false|false|false|C0817321|Right tibia|right tibia
Anatomy|Body Part, Organ, or Organ Component|General Exam|6522,6527|false|false|false|C0040184|Bone structure of tibia|tibia
Finding|Finding|General Exam|6536,6539|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Finding|Gene or Genome|General Exam|6536,6539|false|false|false|C0948106;C1419600|ROM1 gene;Rupture of Membranes|ROM
Procedure|Laboratory Procedure|General Exam|6536,6539|false|false|false|C1562926|Range of motion technique (procedure)|ROM
Attribute|Clinical Attribute|General Exam|6547,6551|false|true|false|C2598155||pain
Finding|Functional Concept|General Exam|6547,6551|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|6547,6551|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|General Exam|6566,6570|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|6566,6570|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|6566,6570|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|6566,6570|false|false|false|C0562271|Examination of knee joint|knee
Finding|Finding|General Exam|6566,6578|false|false|false|C0240114|Knee flexion|knee flexion
Attribute|Clinical Attribute|General Exam|6571,6578|false|true|false|C1525443|W flexion|flexion
Finding|Organ or Tissue Function|General Exam|6571,6578|false|true|false|C0231452||flexion
Anatomy|Body Part, Organ, or Organ Component|General Exam|6594,6597|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Conceptual Entity|General Exam|6608,6617|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Finding|Functional Concept|General Exam|6608,6617|false|false|false|C0231448;C1880641|Extension;Telephone Extension Number|extension
Drug|Food|General Exam|6635,6641|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|6635,6641|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|6635,6641|false|false|false|C0034107|Pulse taking|pulses
Anatomy|Body System|General Exam|6655,6659|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|6655,6659|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|6655,6659|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|6655,6659|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|6655,6659|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Disorder|Disease or Syndrome|General Exam|6661,6675|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|6670,6675|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|6670,6675|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|6685,6690|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|6685,6690|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|6685,6702|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|6691,6702|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Anatomy|Body Location or Region|General Exam|6712,6717|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|6712,6717|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|6712,6727|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|6718,6727|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|General Exam|6728,6737|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|6728,6737|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|6728,6737|false|false|false|C2229507|sensory exam|sensation
Finding|Intellectual Product|General Exam|6741,6746|false|false|false|C1549782|Relational Operator - Equal|equal
Drug|Amino Acid, Peptide, or Protein|General Exam|6764,6769|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|6764,6769|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|6764,6769|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|6764,6769|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|6764,6769|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|6764,6769|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|6764,6769|false|false|false|C0031765|Phototherapy|light
Finding|Mental Process|General Exam|6770,6775|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|6770,6775|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|6770,6775|false|false|false|C0152054|Therapeutic Touch|touch
Anatomy|Body Location or Region|General Exam|6794,6799|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|6794,6799|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|6794,6809|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|6800,6809|false|false|false|C0015385|Limb structure|extremity
Finding|Idea or Concept|General Exam|6810,6818|false|false|false|C0808080|Strength (attribute)|strength
Finding|Classification|General Exam|6820,6828|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|General Exam|6820,6828|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|General Exam|6820,6828|false|false|false|C5237010|Expression Negative|Negative
Finding|Functional Concept|General Exam|6901,6906|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|6907,6913|false|false|false|C0040184|Bone structure of tibia|tibial
Attribute|Clinical Attribute|General Exam|6914,6918|false|false|false|C2598155||pain
Finding|Functional Concept|General Exam|6914,6918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|6914,6918|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Health Care Activity|General Exam|6940,6949|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|6950,6954|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|6985,6990|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|6985,6990|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|6991,6994|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|6999,7002|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|6999,7002|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|6999,7002|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|7009,7012|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|7009,7012|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|7009,7012|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|7009,7012|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|7019,7022|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|7019,7022|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|7030,7033|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|7030,7033|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|7030,7033|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|7030,7033|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|7037,7040|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|7037,7040|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|7037,7040|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|7037,7040|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|7037,7040|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|7046,7050|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|7077,7080|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|7097,7102|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7097,7102|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|7119,7124|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|7119,7124|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|7119,7124|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|7131,7134|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|7131,7134|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|7234,7239|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7234,7239|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|7244,7247|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|7244,7247|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|7269,7274|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7269,7274|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|7269,7282|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|7269,7282|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|7269,7282|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|7275,7282|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|7275,7282|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|7275,7282|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|7275,7282|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|7275,7282|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|7327,7331|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|7327,7331|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|7327,7331|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|7356,7361|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7356,7361|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|7356,7369|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|7362,7369|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|7362,7369|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|7362,7369|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|7362,7369|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|7362,7369|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|7362,7369|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|7362,7369|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|General Exam|7391,7395|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|7391,7395|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|7391,7395|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|General Exam|7391,7395|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|General Exam|7411,7416|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7411,7416|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|7451,7454|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|7451,7454|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|7451,7454|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|7451,7454|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|7451,7454|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|General Exam|7471,7476|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7471,7476|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|7499,7504|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7499,7504|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|7499,7512|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|7505,7512|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|7505,7512|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|7505,7512|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|General Exam|7518,7527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|7518,7527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|7518,7527|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|7518,7527|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|General Exam|7528,7532|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|7563,7568|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7563,7568|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|7569,7572|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|7577,7580|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7577,7580|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7577,7580|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|7587,7590|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|7587,7590|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|7587,7590|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|7587,7590|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|7597,7600|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|7597,7600|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|7608,7611|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|7608,7611|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|7608,7611|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|7608,7611|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|7615,7618|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|7615,7618|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|7615,7618|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|7615,7618|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|7615,7618|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|7624,7628|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|7655,7658|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|7675,7680|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7675,7680|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|7697,7702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7697,7702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|7697,7710|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|7697,7710|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|7697,7710|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|7703,7710|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|7703,7710|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|7703,7710|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|7703,7710|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|7703,7710|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|7756,7760|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|7756,7760|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|7756,7760|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|7785,7790|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|7785,7790|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|7785,7798|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|7791,7798|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|7791,7798|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|7791,7798|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|7791,7798|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|7791,7798|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|7791,7798|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|7791,7798|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Finding|General Exam|7820,7827|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|7820,7827|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Anatomy|Body Location or Region|General Exam|7856,7861|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7856,7861|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7856,7871|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7856,7876|false|false|false|C0226813;C4266545|Lower extremity>Lower extremity veins;Structure of vein of lower extremity|lower extremity vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|7862,7871|false|false|false|C0015385|Limb structure|extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7862,7876|false|false|false|C0730267|Venous structure of limb|extremity vein
Anatomy|Body Part, Organ, or Organ Component|General Exam|7872,7876|false|false|false|C0042449|Veins|vein
Finding|Functional Concept|General Exam|7884,7889|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Location or Region|General Exam|7884,7894|false|false|false|C0489801|Posterior part of right leg|Right calf
Anatomy|Body Location or Region|General Exam|7890,7894|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|7890,7894|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Idea or Concept|General Exam|7931,7939|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|7931,7942|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|General Exam|7943,7947|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|General Exam|7948,7954|false|false|false|C0042449|Veins|venous
Finding|Finding|General Exam|7948,7965|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|General Exam|7948,7965|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|General Exam|7955,7965|false|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|General Exam|7973,7978|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|7973,7994|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|General Exam|7979,7984|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|7979,7984|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|7979,7994|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7979,8000|false|false|false|C0226813;C4266545|Lower extremity>Lower extremity veins;Structure of vein of lower extremity|lower extremity veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|7985,7994|false|false|false|C0015385|Limb structure|extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|7985,8000|false|false|false|C0730267|Venous structure of limb|extremity veins
Anatomy|Body Part, Organ, or Organ Component|General Exam|7995,8000|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|7995,8000|false|false|false|C0398102|Procedure on vein|veins
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|8027,8035|false|false|false|C0009924|Contrast Media|contrast
Finding|Functional Concept|General Exam|8055,8060|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|8055,8065|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|General Exam|8061,8065|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|8061,8065|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Location or Region|General Exam|8078,8084|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|General Exam|8078,8084|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|General Exam|8099,8103|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|General Exam|8099,8103|false|false|false|C0555980|Foot problem|foot
Anatomy|Body Part, Organ, or Organ Component|General Exam|8110,8115|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|General Exam|8110,8115|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|General Exam|8123,8128|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|8123,8128|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|8123,8138|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|8129,8138|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|General Exam|8210,8216|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Functional Concept|General Exam|8217,8227|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|8217,8227|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|8217,8227|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Conceptual Entity|General Exam|8263,8273|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|8263,8273|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|8263,8273|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|8263,8273|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Part, Organ, or Organ Component|General Exam|8285,8293|false|false|false|C4083049|Muscle (organ)|muscular
Disorder|Anatomical Abnormality|General Exam|8285,8305|true|false|false|C4021745|Abnormality of the musculature|muscular abnormality
Disorder|Congenital Abnormality|General Exam|8294,8305|true|false|false|C0000768|Congenital Abnormality|abnormality
Finding|Finding|General Exam|8294,8305|true|false|false|C1704258|Abnormality|abnormality
Finding|Finding|General Exam|8335,8345|false|false|false|C5453124|Uneventful|Uneventful
Finding|Functional Concept|General Exam|8346,8356|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|General Exam|8346,8356|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|General Exam|8346,8356|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Drug|Biomedical or Dental Material|General Exam|8364,8373|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|General Exam|8364,8373|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|General Exam|8364,8373|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Drug|Pharmacologic Substance|General Exam|8390,8400|false|false|false|C0002932;C5399725|Anesthetic [APC];Anesthetics|anesthetic
Drug|Organic Chemical|General Exam|8405,8412|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|General Exam|8405,8412|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Anatomy|Body Part, Organ, or Organ Component|General Exam|8435,8453|false|false|false|C0224813|Structure of trochanteric bursa|trochanteric bursa
Anatomy|Body Part, Organ, or Organ Component|General Exam|8448,8453|false|false|false|C0006441|Synovial bursa|bursa
Drug|Biomedical or Dental Material|General Exam|8465,8474|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|General Exam|8465,8474|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|General Exam|8465,8474|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Intellectual Product|General Exam|8482,8488|false|false|false|C1561574|Amount class - Amount|amount
Drug|Substance|General Exam|8492,8497|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|8492,8497|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Functional Concept|General Exam|8505,8510|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|General Exam|8533,8538|false|false|false|C0006441|Synovial bursa|bursa
Finding|Functional Concept|General Exam|8543,8553|false|false|false|C0333607|dystrophic|dystrophic
Finding|Finding|General Exam|8543,8567|false|false|false|C0333582|Dystrophic calcification|dystrophic calcification
Finding|Organ or Tissue Function|General Exam|8554,8567|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Finding|Pathologic Function|General Exam|8554,8567|false|false|false|C0006660;C0006663;C1533591|Calcification;Calcinosis;Physiologic calcification|calcification
Phenomenon|Natural Phenomenon or Process|General Exam|8586,8591|false|false|false|C0282173|Space (Astronomy)|space
Finding|Mental Process|Findings|8610,8619|false|false|false|C0242114|Suspicion|suspicion
Finding|Intellectual Product|Findings|8624,8631|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Findings|8624,8631|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Findings|8632,8653|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Findings|8645,8653|false|false|false|C0006444|Bursitis|bursitis
Finding|Intellectual Product|Hospital Course|8680,8687|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Finding|Finding|Hospital Course|8732,8735|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Finding|Idea or Concept|Hospital Course|8736,8747|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Hospital Course|8753,8778|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid syndrome
Disorder|Disease or Syndrome|Hospital Course|8770,8778|false|false|false|C0039082|Syndrome|syndrome
Disorder|Disease or Syndrome|Hospital Course|8784,8788|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8793,8796|false|false|false|C0016504;C0687080;C1690938;C3853547|Foot;Hindfoot of quadruped;Paw;Structure of ankle and/or foot (body structure)|PEs
Finding|Gene or Genome|Hospital Course|8793,8796|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Finding|Intellectual Product|Hospital Course|8793,8796|false|false|false|C0687136;C1418467|PES1 gene;Personal Experience Scales|PEs
Drug|Organic Chemical|Hospital Course|8800,8808|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|8800,8808|false|false|false|C0699129|Coumadin|Coumadin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8826,8832|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|8826,8832|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|8826,8832|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8826,8832|false|false|false|C0191838|Procedures on breast|breast
Disorder|Neoplastic Process|Hospital Course|8826,8839|false|false|false|C0006142;C0678222|Breast Carcinoma;Malignant neoplasm of breast|breast cancer
Disorder|Neoplastic Process|Hospital Course|8833,8839|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8844,8854|false|false|false|C0851238;C1262070|Excision of mass (procedure);Lumpectomy of breast|lumpectomy
Finding|Intellectual Product|Hospital Course|8886,8891|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|8895,8902|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|8895,8902|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|Hospital Course|8903,8908|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8903,8924|false|false|false|C0230415|Right lower extremity|right lower extremity
Anatomy|Body Location or Region|Hospital Course|8909,8914|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|8909,8914|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8909,8924|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8915,8924|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|Hospital Course|8929,8934|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|8929,8938|false|false|false|C0524470|Right hip region structure|right hip
Finding|Sign or Symptom|Hospital Course|8929,8943|false|true|false|C2202100|Pain of right hip joint|right hip pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8935,8938|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8935,8938|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|8935,8938|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|8935,8938|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|8935,8938|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8935,8938|false|false|false|C1292890|Procedure on hip|hip
Attribute|Clinical Attribute|Hospital Course|8935,8943|false|true|false|C1716793||hip pain
Finding|Sign or Symptom|Hospital Course|8935,8943|false|true|false|C0019559;C4551516|Hip joint pain;Hip pain|hip pain
Attribute|Clinical Attribute|Hospital Course|8939,8943|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8939,8943|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8939,8943|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|8956,8965|false|false|false|C0332218|Difficult (qualifier value)|difficult
Finding|Functional Concept|Hospital Course|8979,8984|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8979,9000|false|false|false|C0230415|Right lower extremity|Right lower extremity
Anatomy|Body Location or Region|Hospital Course|8985,8990|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|8985,8990|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8985,9000|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8991,9000|false|false|false|C0015385|Limb structure|extremity
Anatomy|Body Location or Region|Hospital Course|9030,9033|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9030,9033|true|true|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9030,9033|true|true|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Anatomy|Body Location or Region|Hospital Course|9041,9045|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9041,9045|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9046,9051|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9046,9051|false|false|false|C0398102|Procedure on vein|veins
Finding|Finding|Hospital Course|9061,9065|true|true|false|C5575035|Well (answer to question)|well
Finding|Functional Concept|Hospital Course|9117,9122|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|9117,9144|false|false|false|C3862456|right trochanteric bursitis|Right trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|9123,9144|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|9136,9144|false|false|false|C0006444|Bursitis|bursitis
Finding|Functional Concept|Hospital Course|9147,9152|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|9153,9161|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|Hospital Course|9162,9167|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|9162,9167|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9162,9171|false|false|false|C1140621;C4299093|Leg;Lower extremity>Lower leg|lower leg
Finding|Sign or Symptom|Hospital Course|9162,9176|false|true|false|C0023222;C0839480|Pain in limb, lower leg;Pain in lower limb|lower leg pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9168,9171|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|9168,9176|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Hospital Course|9172,9176|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9172,9176|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9172,9176|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|9179,9184|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|9191,9205|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9200,9205|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9200,9205|false|false|false|C0398102|Procedure on vein|veins
Attribute|Clinical Attribute|Hospital Course|9228,9232|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9228,9232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9228,9232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|9260,9265|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Hospital Course|9260,9265|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Hospital Course|9295,9302|false|false|false|C1555582|Initial (abbreviation)|initial
Finding|Functional Concept|Hospital Course|9303,9307|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|9303,9307|false|false|false|C0582103|Medical Examination|exam
Finding|Idea or Concept|Hospital Course|9317,9327|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|9317,9332|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|Hospital Course|9334,9340|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|9334,9340|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|9341,9362|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|9354,9362|false|false|false|C0006444|Bursitis|bursitis
Finding|Functional Concept|Hospital Course|9370,9375|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Attribute|Clinical Attribute|Hospital Course|9402,9406|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9402,9406|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9402,9406|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|9417,9422|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9417,9428|false|false|false|C0817321|Right tibia|right tibia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9423,9428|false|false|false|C0040184|Bone structure of tibia|tibia
Finding|Idea or Concept|Hospital Course|9454,9464|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|9454,9469|false|false|false|C0332290|Consistent with|consistent with
Attribute|Clinical Attribute|Hospital Course|9470,9474|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9470,9474|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9470,9474|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|Hospital Course|9484,9498|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9493,9498|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9493,9498|false|false|false|C0398102|Procedure on vein|veins
Finding|Finding|Hospital Course|9504,9507|false|false|false|C1860232|X-RAY SENSITIVITY|XRs
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9516,9521|false|false|false|C0040184|Bone structure of tibia|tibia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9522,9528|false|false|false|C0016068|Fibula|fibula
Finding|Functional Concept|Hospital Course|9533,9538|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|9533,9542|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9539,9542|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9539,9542|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|9539,9542|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|9539,9542|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|9539,9542|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9539,9542|false|false|false|C1292890|Procedure on hip|hip
Finding|Functional Concept|Hospital Course|9564,9573|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Finding|Pathologic Function|Hospital Course|9564,9573|false|false|false|C0205469;C0677042|Pathological aspects;Pathology processes|pathology
Procedure|Laboratory Procedure|Hospital Course|9564,9573|false|false|false|C0919386|Pathology procedure|pathology
Finding|Sign or Symptom|Hospital Course|9600,9619|true|false|false|C0235031|Neurologic Symptoms|neurologic symptoms
Finding|Functional Concept|Hospital Course|9611,9619|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|9611,9619|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|Hospital Course|9634,9647|false|false|false|C0700594|Radiculopathy|radiculopathy
Finding|Sign or Symptom|Hospital Course|9652,9660|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|Hospital Course|9664,9672|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Hospital Course|9664,9672|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Intellectual Product|Hospital Course|9699,9705|false|false|false|C0542560|Academic degree|degree
Finding|Intellectual Product|Hospital Course|9709,9716|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|9709,9716|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|9709,9725|false|false|false|C0585052|Chronic sciatica|chronic sciatica
Finding|Sign or Symptom|Hospital Course|9717,9725|false|false|false|C0036396|Sciatica|sciatica
Finding|Finding|Hospital Course|9728,9744|false|false|false|C5425896|Mildly decreased|Mildly decreased
Finding|Finding|Hospital Course|9735,9760|false|false|false|C3277184|Decreased patellar reflex|decreased patellar reflex
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9745,9753|false|false|false|C0030647|Patella|patellar
Finding|Finding|Hospital Course|9745,9760|false|false|false|C0234147|Knee reflex|patellar reflex
Finding|Finding|Hospital Course|9754,9760|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Finding|Organ or Tissue Function|Hospital Course|9754,9760|false|false|false|C0034929;C0439840;C0596002|Observation of reflex;Reflex action;Reflex motion descriptor|reflex
Finding|Functional Concept|Hospital Course|9769,9774|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Functional Concept|Hospital Course|9790,9794|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Mental Process|Hospital Course|9816,9823|false|false|false|C0542559|contextual factors|setting
Attribute|Clinical Attribute|Hospital Course|9828,9832|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|9828,9832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|9828,9832|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|9837,9845|false|false|false|C0427198|Protective muscle spasm|guarding
Finding|Idea or Concept|Hospital Course|9847,9855|false|false|false|C0808080|Strength (attribute)|strength
Finding|Finding|Hospital Course|9891,9900|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Hospital Course|9891,9900|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Hospital Course|9891,9900|false|false|false|C2229507|sensory exam|sensation
Drug|Organic Chemical|Hospital Course|9928,9935|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|9928,9935|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9928,9945|false|false|false|C1261311|Injection of steroid|steroid injection
Drug|Biomedical or Dental Material|Hospital Course|9936,9945|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|Hospital Course|9936,9945|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9936,9945|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9967,9972|false|false|false|C0006441|Synovial bursa|bursa
Finding|Idea or Concept|Hospital Course|9976,9987|false|false|false|C0750502|Significant|significant
Finding|Conceptual Entity|Hospital Course|9988,9999|false|false|false|C2986411|Improvement|improvement
Finding|Functional Concept|Hospital Course|10003,10011|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|10003,10011|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Substance|Hospital Course|10045,10050|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|10045,10050|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10060,10065|false|false|false|C0006441|Synovial bursa|bursa
Finding|Functional Concept|Hospital Course|10067,10077|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|10067,10080|false|false|false|C0332299|Suggestive of|suggestive of
Finding|Intellectual Product|Hospital Course|10081,10086|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|10091,10098|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|10091,10098|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|10099,10120|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|10112,10120|false|false|false|C0006444|Bursitis|bursitis
Disorder|Disease or Syndrome|Hospital Course|10126,10134|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|Hospital Course|10135,10139|false|false|false|C0230444|Shin|shin
Finding|Sign or Symptom|Hospital Course|10135,10144|false|false|false|C0241032|shin pain|shin pain
Attribute|Clinical Attribute|Hospital Course|10140,10144|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|10140,10144|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10140,10144|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|10160,10170|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|Hospital Course|10160,10170|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|Hospital Course|10160,10170|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Organic Chemical|Hospital Course|10174,10184|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|10174,10184|false|false|false|C0060926|gabapentin|gabapentin
Drug|Organic Chemical|Hospital Course|10189,10198|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|10189,10198|false|false|false|C0023660|lidocaine|lidocaine
Procedure|Laboratory Procedure|Hospital Course|10189,10198|false|false|false|C0202404|Lidocaine measurement|lidocaine
Drug|Clinical Drug|Hospital Course|10189,10204|false|false|false|C1251704|Lidocaine Patch|lidocaine patch
Drug|Biomedical or Dental Material|Hospital Course|10199,10204|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|Hospital Course|10199,10204|false|false|false|C0332461|Plaque (lesion)|patch
Finding|Functional Concept|Hospital Course|10205,10219|false|false|false|C0332287|In addition to|in addition to
Finding|Functional Concept|Hospital Course|10208,10216|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Finding|Idea or Concept|Hospital Course|10225,10229|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10225,10229|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10225,10229|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10230,10237|false|false|false|C0699142|Tylenol|tylenol
Drug|Pharmacologic Substance|Hospital Course|10230,10237|false|false|false|C0699142|Tylenol|tylenol
Finding|Functional Concept|Hospital Course|10245,10253|false|false|false|C0442805|Increase|increase
Finding|Intellectual Product|Hospital Course|10261,10270|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Finding|Idea or Concept|Hospital Course|10278,10282|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10278,10282|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10278,10282|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10284,10292|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|10284,10292|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|Hospital Course|10284,10292|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Finding|Gene or Genome|Hospital Course|10298,10301|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Gene or Genome|Hospital Course|10309,10312|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Idea or Concept|Hospital Course|10337,10341|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10337,10341|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10337,10341|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10343,10356|false|false|false|C0012306|hydromorphone|hydromorphone
Drug|Pharmacologic Substance|Hospital Course|10343,10356|false|false|false|C0012306|hydromorphone|hydromorphone
Finding|Gene or Genome|Hospital Course|10357,10360|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|10408,10421|false|false|false|C0012306|hydromorphone|hydromorphone
Drug|Pharmacologic Substance|Hospital Course|10408,10421|false|false|false|C0012306|hydromorphone|hydromorphone
Drug|Biomedical or Dental Material|Hospital Course|10436,10445|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|Hospital Course|10436,10445|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10436,10445|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Mental Process|Hospital Course|10453,10460|false|false|false|C0542559|contextual factors|setting
Finding|Intellectual Product|Hospital Course|10467,10472|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|Hospital Course|10474,10478|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|10474,10478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|10474,10478|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|10512,10520|false|false|false|C0040610|tramadol|Tramadol
Drug|Pharmacologic Substance|Hospital Course|10512,10520|false|false|false|C0040610|tramadol|Tramadol
Procedure|Laboratory Procedure|Hospital Course|10512,10520|false|false|false|C1266765|Tramadol measurement (procedure)|Tramadol
Drug|Biomedical or Dental Material|Hospital Course|10530,10537|false|false|false|C0039225|Tablet Dosage Form|tablets
Finding|Pathologic Function|Hospital Course|10545,10566|false|false|false|C0520917|Increased metabolic requirement|increased requirement
Finding|Functional Concept|Hospital Course|10555,10566|false|false|false|C1514873|Requirement|requirement
Finding|Body Substance|Hospital Course|10571,10580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10571,10580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10571,10580|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10571,10580|false|false|false|C0030685|Patient Discharge|discharge
Finding|Finding|Hospital Course|10590,10594|false|false|false|C1299581|Able (qualifier value)|able
Finding|Finding|Hospital Course|10595,10603|false|false|false|C4036205|Ambulate|ambulate
Finding|Intellectual Product|Hospital Course|10618,10622|false|false|false|C4684764|SAFE-Biopharma Standard|safe
Finding|Body Substance|Hospital Course|10627,10636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10627,10636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10627,10636|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10627,10636|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10627,10641|false|false|false|C0184713|Discharge to home|discharge home
Finding|Idea or Concept|Hospital Course|10637,10641|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10637,10641|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10637,10641|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|10663,10673|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|10663,10673|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Mental Process|Hospital Course|10683,10688|false|false|false|C0558083|Enthusiastic|eager
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10725,10733|false|false|false|C0005847|Blood Vessel|vascular
Attribute|Clinical Attribute|Hospital Course|10734,10741|false|false|false|C5444295||surgeon
Event|Activity|Hospital Course|10749,10760|false|false|false|C0003629|Appointments|appointment
Finding|Finding|Hospital Course|10774,10777|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|10774,10777|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|10778,10782|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|10778,10782|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Conceptual Entity|Hospital Course|10788,10797|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|10788,10797|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|10788,10797|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10788,10797|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Sign or Symptom|Hospital Course|10805,10812|false|false|false|C0030193|Pain|painful
Disorder|Disease or Syndrome|Hospital Course|10813,10827|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10822,10827|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10822,10827|false|false|false|C0398102|Procedure on vein|veins
Drug|Biologically Active Substance|Hospital Course|10832,10836|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|10832,10836|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|10832,10836|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|Hospital Course|10832,10836|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|Hospital Course|10832,10847|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|Iron deficiency
Disorder|Disease or Syndrome|Hospital Course|10832,10854|false|false|false|C0162316|Iron deficiency anemia|Iron deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|10837,10847|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|10837,10847|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Hospital Course|10837,10854|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|10848,10854|false|false|false|C0002871|Anemia|anemia
Disorder|Disease or Syndrome|Hospital Course|10856,10862|false|false|false|C0002871|Anemia|Anemia
Finding|Finding|Hospital Course|10866,10869|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|10866,10869|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|10937,10944|true|false|false|C2699424|Concern|concern
Finding|Pathologic Function|Hospital Course|10956,10964|true|false|false|C0019080|Hemorrhage|bleeding
Drug|Biologically Active Substance|Hospital Course|10970,10974|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|10970,10974|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|10970,10974|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|10970,10974|false|false|false|C0337439|Iron measurement|iron
Procedure|Laboratory Procedure|Hospital Course|10970,10982|false|false|false|C2079295|iron studies|iron studies
Procedure|Research Activity|Hospital Course|10975,10982|false|false|false|C0947630|Scientific Study|studies
Drug|Biologically Active Substance|Hospital Course|10992,10996|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|10992,10996|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|10992,10996|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|10992,10996|false|false|false|C0337439|Iron measurement|iron
Finding|Functional Concept|Hospital Course|10997,11006|false|false|false|C0011155|Deficiency|deficient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11014,11022|false|false|false|C0015879|Ferritin|ferritin
Drug|Biologically Active Substance|Hospital Course|11014,11022|false|false|false|C0015879|Ferritin|ferritin
Drug|Pharmacologic Substance|Hospital Course|11014,11022|false|false|false|C0015879|Ferritin|ferritin
Procedure|Laboratory Procedure|Hospital Course|11014,11022|false|false|false|C0373607|Ferritin measurement|ferritin
Finding|Sign or Symptom|Hospital Course|11044,11051|false|false|false|C0015672|Fatigue|fatigue
Finding|Sign or Symptom|Hospital Course|11056,11064|false|false|false|C0085631;C3887611|Agitation;Restlessness|restless
Disorder|Disease or Syndrome|Hospital Course|11056,11068|false|false|false|C0035258|Restless Legs Syndrome|restless leg
Disorder|Disease or Syndrome|Hospital Course|11056,11077|false|false|false|C0035258|Restless Legs Syndrome|restless leg syndrome
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11065,11068|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Disorder|Disease or Syndrome|Hospital Course|11069,11077|false|false|false|C0039082|Syndrome|syndrome
Finding|Conceptual Entity|Hospital Course|11079,11087|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|Hospital Course|11079,11087|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|Hospital Course|11140,11144|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11140,11151|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11145,11151|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|11145,11151|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|11145,11151|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11145,11151|false|false|false|C0191838|Procedures on breast|breast
Finding|Pathologic Function|Hospital Course|11145,11160|false|false|false|C0342095|Breast hematoma|breast hematoma
Finding|Pathologic Function|Hospital Course|11152,11160|false|false|false|C0018944|Hematoma|hematoma
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11169,11175|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|11169,11175|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|11169,11175|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11169,11175|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Hospital Course|11177,11185|false|false|false|C0750558|Unlikely|unlikely
Finding|Intellectual Product|Hospital Course|11197,11203|false|false|false|C1704250|Timing, LOINC Axis 3|timing
Finding|Sign or Symptom|Hospital Course|11204,11208|false|false|false|C0036572|Seizures|fits
Procedure|Diagnostic Procedure|Hospital Course|11217,11220|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Disorder|Disease or Syndrome|Hospital Course|11227,11236|false|false|false|C0017152|Gastritis|gastritis
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11265,11268|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11265,11268|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11265,11268|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11265,11268|false|false|false|C1332410|BID gene|BID
Drug|Pharmacologic Substance|Hospital Course|11269,11272|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|11269,11272|false|false|false|C0871125|Prepulse Inhibition|PPI
Procedure|Diagnostic Procedure|Hospital Course|11281,11292|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|11281,11292|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Attribute|Clinical Attribute|Hospital Course|11302,11310|false|false|false|C2926606||findings
Finding|Functional Concept|Hospital Course|11302,11310|false|false|false|C2607943|findings aspects|findings
Finding|Functional Concept|Hospital Course|11323,11333|false|false|false|C0332299|Suggestive of|suggestive
Finding|Functional Concept|Hospital Course|11323,11336|false|true|false|C0332299|Suggestive of|suggestive of
Disorder|Disease or Syndrome|Hospital Course|11338,11344|false|false|false|C0007570|Celiac Disease|celiac
Disorder|Disease or Syndrome|Hospital Course|11338,11352|false|false|false|C0007570|Celiac Disease|celiac disease
Finding|Gene or Genome|Hospital Course|11338,11352|false|false|false|C1332802|CTLA4 gene|celiac disease
Disorder|Disease or Syndrome|Hospital Course|11345,11352|false|false|false|C0012634|Disease|disease
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11361,11364|false|false|false|C5565118|TGM2 protein, human|ttg
Drug|Enzyme|Hospital Course|11361,11364|false|false|false|C5565118|TGM2 protein, human|ttg
Drug|Pharmacologic Substance|Hospital Course|11361,11364|false|false|false|C5565118|TGM2 protein, human|ttg
Finding|Gene or Genome|Hospital Course|11361,11364|false|false|false|C5575307|TGM2 wt Allele|ttg
Finding|Finding|Hospital Course|11373,11377|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|11373,11377|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|11373,11377|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11404,11407|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Immunologic Factor|Hospital Course|11404,11407|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Drug|Pharmacologic Substance|Hospital Course|11404,11407|false|false|false|C0020835;C2825347|immunoglobulin A;immunoglobulin A, human|IgA
Finding|Gene or Genome|Hospital Course|11404,11407|false|false|false|C1413238;C3273407|CD79A gene;CD79A wt Allele|IgA
Procedure|Laboratory Procedure|Hospital Course|11404,11407|false|false|false|C0202083|Immunoglobulin A measurement|IgA
Disorder|Anatomical Abnormality|Hospital Course|11426,11432|false|false|false|C0032584|polyps|polyps
Finding|Intellectual Product|Hospital Course|11426,11432|false|false|false|C1546747||polyps
Procedure|Health Care Activity|Hospital Course|11468,11477|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Organic Chemical|Hospital Course|11479,11488|false|false|false|C0042839|vitamin A|a vitamin
Drug|Pharmacologic Substance|Hospital Course|11479,11488|false|false|false|C0042839|vitamin A|a vitamin
Drug|Vitamin|Hospital Course|11479,11488|false|false|false|C0042839|vitamin A|a vitamin
Drug|Pharmacologic Substance|Hospital Course|11479,11490|false|false|false|C0310589|Vitamins A and D preparation|a vitamin D
Drug|Organic Chemical|Hospital Course|11481,11488|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|11481,11488|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|11481,11488|false|false|false|C0042890|Vitamins|vitamin
Drug|Hormone|Hospital Course|11481,11490|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Organic Chemical|Hospital Course|11481,11490|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Pharmacologic Substance|Hospital Course|11481,11490|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Vitamin|Hospital Course|11481,11490|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Procedure|Laboratory Procedure|Hospital Course|11481,11490|false|false|false|C0919758|Vitamin D measurement|vitamin D
Finding|Idea or Concept|Hospital Course|11524,11532|false|false|false|C3887511|Evidence|evidence
Disorder|Disease or Syndrome|Hospital Course|11537,11550|false|false|false|C0024523|Malabsorption Syndrome|malabsorption
Finding|Finding|Hospital Course|11537,11550|false|false|false|C3714745|Malabsorption|malabsorption
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11561,11576|false|false|false|C0242297|Dietary Supplementation|supplementation
Drug|Inorganic Chemical|Hospital Course|11607,11613|false|false|false|C3848561|ferric cation|ferric
Drug|Pharmacologic Substance|Hospital Course|11607,11613|false|false|false|C3848561|ferric cation|ferric
Drug|Organic Chemical|Hospital Course|11607,11623|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Pharmacologic Substance|Hospital Course|11607,11623|false|false|false|C0060235|ferric gluconate|ferric gluconate
Drug|Biologically Active Substance|Hospital Course|11614,11623|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Organic Chemical|Hospital Course|11614,11623|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Pharmacologic Substance|Hospital Course|11614,11623|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11638,11641|false|false|false|C5565118|TGM2 protein, human|TTG
Drug|Enzyme|Hospital Course|11638,11641|false|false|false|C5565118|TGM2 protein, human|TTG
Drug|Pharmacologic Substance|Hospital Course|11638,11641|false|false|false|C5565118|TGM2 protein, human|TTG
Finding|Gene or Genome|Hospital Course|11638,11641|false|false|false|C5575307|TGM2 wt Allele|TTG
Finding|Idea or Concept|Hospital Course|11660,11667|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Finding|Body Substance|Hospital Course|11671,11680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11671,11680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11671,11680|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11671,11680|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|Hospital Course|11684,11691|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|11684,11691|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Conceptual Entity|Hospital Course|11722,11729|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|11722,11729|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|11722,11729|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|11722,11732|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|11733,11736|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|11733,11736|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|11733,11736|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11740,11751|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|11743,11751|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|11743,11751|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|11743,11751|false|false|false|C0043031|warfarin|warfarin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11755,11780|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Drug|Immunologic Factor|Hospital Course|11755,11780|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Finding|Finding|Hospital Course|11755,11780|false|false|false|C4019436|Antiphospholipid antibody positivity|Antiphospholipid antibody
Disorder|Disease or Syndrome|Hospital Course|11755,11789|false|false|false|C0085278|Antiphospholipid Syndrome|Antiphospholipid antibody syndrome
Anatomy|Cell Component|Hospital Course|11772,11780|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11772,11780|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Hospital Course|11772,11780|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Hospital Course|11772,11780|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Hospital Course|11772,11780|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Hospital Course|11781,11789|false|false|false|C0039082|Syndrome|syndrome
Finding|Finding|Hospital Course|11793,11811|false|false|false|C1168145|Anticoagulation drug level below therapeutic|Subtherapeutic INR
Attribute|Clinical Attribute|Hospital Course|11808,11811|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|11808,11811|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11808,11811|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Disorder|Disease or Syndrome|Hospital Course|11813,11818|false|false|false|C0024131;C0024138;C0024141;C0409974;C5574816|Chronic discoid lupus erythematosus;Discoid lupus erythematosus;Lupus Erythematosus;Lupus Erythematosus, Systemic;Lupus Vulgaris|Lupus
Disorder|Disease or Syndrome|Hospital Course|11813,11832|false|false|false|C0311370|Lupus anticoagulant disorder|Lupus anticoagulant
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11813,11832|false|false|false|C0085240|Lupus Coagulation Inhibitor|Lupus anticoagulant
Drug|Immunologic Factor|Hospital Course|11813,11832|false|false|false|C0085240|Lupus Coagulation Inhibitor|Lupus anticoagulant
Finding|Finding|Hospital Course|11813,11832|false|false|false|C4321325||Lupus anticoagulant
Procedure|Laboratory Procedure|Hospital Course|11813,11832|false|false|false|C1142517|Lupus anticoagulant assay|Lupus anticoagulant
Lab|Laboratory or Test Result|Hospital Course|11813,11841|false|false|false|C1142516|Lupus anticoagulant positive|Lupus anticoagulant positive
Drug|Pharmacologic Substance|Hospital Course|11819,11832|false|false|false|C0003280;C3536711|Anti-coagulant [EPC];Anticoagulants|anticoagulant
Finding|Idea or Concept|Hospital Course|11875,11879|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11875,11879|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11875,11879|false|false|false|C1553498|home health encounter|home
Drug|Hazardous or Poisonous Substance|Hospital Course|11888,11896|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|11888,11896|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|11888,11896|false|false|false|C0043031|warfarin|warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|11936,11944|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|11936,11944|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|11936,11944|false|false|false|C0043031|warfarin|warfarin
Finding|Pathologic Function|Hospital Course|11967,11975|false|false|false|C0018944|Hematoma|hematoma
Drug|Organic Chemical|Hospital Course|12006,12013|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Hospital Course|12006,12013|false|false|false|C0728963|Lovenox|Lovenox
Attribute|Clinical Attribute|Hospital Course|12033,12036|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|12033,12036|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12033,12036|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Health Care Activity|Hospital Course|12045,12054|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Procedure|Health Care Activity|Hospital Course|12103,12118|false|false|false|C0019993|Hospitalization|hospitalization
Drug|Organic Chemical|Hospital Course|12125,12132|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Hospital Course|12125,12132|false|false|false|C0728963|Lovenox|Lovenox
Finding|Idea or Concept|Hospital Course|12137,12141|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|12137,12141|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Attribute|Clinical Attribute|Hospital Course|12142,12145|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|12142,12145|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12142,12145|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Hazardous or Poisonous Substance|Hospital Course|12187,12195|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|12187,12195|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|12187,12195|false|false|false|C0043031|warfarin|warfarin
Attribute|Clinical Attribute|Hospital Course|12226,12229|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|12226,12229|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12226,12229|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Body Substance|Hospital Course|12233,12242|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|12233,12242|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|12233,12242|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|12233,12242|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|12258,12262|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|Hospital Course|12258,12262|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|12258,12262|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|12258,12262|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Idea or Concept|Hospital Course|12266,12274|false|false|false|C0549178|Continuous|continue
Finding|Idea or Concept|Hospital Course|12275,12279|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|12275,12279|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|12275,12279|false|false|false|C1553498|home health encounter|home
Drug|Hazardous or Poisonous Substance|Hospital Course|12280,12288|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|12280,12288|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|12280,12288|false|false|false|C0043031|warfarin|warfarin
Finding|Intellectual Product|Hospital Course|12289,12296|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12289,12296|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Body Substance|Hospital Course|12298,12305|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|12298,12305|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|12298,12305|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|Hospital Course|12316,12322|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Attribute|Clinical Attribute|Hospital Course|12323,12326|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|12323,12326|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12323,12326|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|Hospital Course|12339,12346|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|12339,12346|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|12339,12346|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|12339,12348|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|12339,12348|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|12339,12348|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|12339,12348|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|12339,12348|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Disorder|Disease or Syndrome|Hospital Course|12339,12359|false|false|false|C0042870|Vitamin D Deficiency|Vitamin D deficiency
Finding|Finding|Hospital Course|12339,12359|false|false|false|C5886864|Decreased circulating vitamin D concentration|Vitamin D deficiency
Disorder|Disease or Syndrome|Hospital Course|12349,12359|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|12349,12359|false|false|false|C0011155|Deficiency|deficiency
Drug|Organic Chemical|Hospital Course|12378,12385|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|12378,12385|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|12378,12385|false|false|false|C0042890|Vitamins|vitamin
Drug|Hormone|Hospital Course|12378,12387|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Organic Chemical|Hospital Course|12378,12387|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Pharmacologic Substance|Hospital Course|12378,12387|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Drug|Vitamin|Hospital Course|12378,12387|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|vitamin D
Procedure|Laboratory Procedure|Hospital Course|12378,12387|false|false|false|C0919758|Vitamin D measurement|vitamin D
Finding|Functional Concept|Hospital Course|12395,12401|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Disorder|Disease or Syndrome|Hospital Course|12438,12451|false|false|false|C0024523|Malabsorption Syndrome|malabsorption
Finding|Finding|Hospital Course|12438,12451|false|false|false|C3714745|Malabsorption|malabsorption
Drug|Biologically Active Substance|Hospital Course|12472,12476|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|12472,12476|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|12472,12476|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|12472,12476|false|false|false|C0337439|Iron measurement|iron
Disorder|Disease or Syndrome|Hospital Course|12472,12487|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|iron deficiency
Disorder|Disease or Syndrome|Hospital Course|12477,12487|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|12477,12487|false|false|false|C0011155|Deficiency|deficiency
Finding|Idea or Concept|Hospital Course|12491,12503|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Occupational Activity|Hospital Course|12533,12537|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|12533,12537|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|Hospital Course|12533,12544|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|Hospital Course|12538,12544|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|12538,12544|false|false|false|C1546481|What subject filter - Status|status
Disorder|Disease or Syndrome|Hospital Course|12561,12564|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Finding|Gene or Genome|Hospital Course|12561,12564|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Functional Concept|Hospital Course|12595,12600|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|12595,12622|false|false|false|C3862456|right trochanteric bursitis|Right trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|12601,12622|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|12614,12622|false|false|false|C0006444|Bursitis|bursitis
Finding|Functional Concept|Hospital Course|12636,12642|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Drug|Biomedical or Dental Material|Hospital Course|12643,12652|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|Hospital Course|12643,12652|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12643,12652|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Finding|Hospital Course|12665,12673|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Hospital Course|12665,12673|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Hospital Course|12665,12673|false|false|false|C0031809|Physical Examination|physical
Finding|Intellectual Product|Hospital Course|12665,12681|false|false|false|C1547999|Diagnostic Service Section ID - Physical Therapy|physical therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12665,12681|false|false|false|C0949766|Physical therapy|physical therapy
Finding|Finding|Hospital Course|12674,12681|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Hospital Course|12674,12681|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12674,12681|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Functional Concept|Hospital Course|12685,12690|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|12691,12699|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12700,12703|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|12700,12708|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Hospital Course|12704,12708|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|12704,12708|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12704,12708|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12726,12736|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|12726,12736|false|false|false|C0060926|gabapentin|gabapentin
Disorder|Disease or Syndrome|Hospital Course|12750,12755|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Drug|Organic Chemical|Hospital Course|12781,12789|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|12781,12789|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|Hospital Course|12781,12789|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Finding|Idea or Concept|Hospital Course|12796,12800|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|12796,12800|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|12796,12800|false|false|false|C1553498|home health encounter|home
Finding|Intellectual Product|Hospital Course|12801,12808|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12801,12808|false|false|false|C0040808|Treatment Protocols|regimen
Procedure|Health Care Activity|Hospital Course|12845,12860|false|false|false|C0019993|Hospitalization|hospitalization
Finding|Idea or Concept|Hospital Course|12876,12879|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|12876,12879|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Activity|Hospital Course|12880,12886|false|false|false|C1999230|Providing (action)|supply
Finding|Functional Concept|Hospital Course|12880,12886|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Finding|Idea or Concept|Hospital Course|12880,12886|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Disorder|Disease or Syndrome|Hospital Course|12907,12911|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|Plan
Finding|Functional Concept|Hospital Course|12907,12911|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Intellectual Product|Hospital Course|12907,12911|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Finding|Mental Process|Hospital Course|12907,12911|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|Plan
Disorder|Disease or Syndrome|Hospital Course|12919,12922|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12919,12922|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|12919,12922|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12919,12922|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|12919,12922|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|12919,12922|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|12919,12922|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|12919,12922|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|12919,12922|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|12919,12922|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Idea or Concept|Hospital Course|12923,12927|false|false|false|C1552851|next - HtmlLinkType|next
Finding|Intellectual Product|Hospital Course|12928,12932|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Classification|Hospital Course|12946,12956|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12946,12956|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Gene or Genome|Hospital Course|12957,12960|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|12957,12960|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|12957,12960|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Location or Region|Hospital Course|12968,12974|false|false|false|C0024090|Lumbar Region|lumbar
Anatomy|Body Location or Region|Hospital Course|12968,12980|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12968,12980|false|false|false|C0024091;C3887615|Bone structure of lumbar vertebra;Lumbar spine structure|lumbar spine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12975,12980|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Hospital Course|12975,12980|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Hospital Course|12975,12980|false|false|false|C0150920|Spine Problem|spine
Finding|Intellectual Product|Hospital Course|12985,12992|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|12985,12992|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|12985,12997|false|false|false|C5700083|chronic pain (diagnosis)|chronic pain
Finding|Sign or Symptom|Hospital Course|12985,12997|false|false|false|C0150055|Chronic pain|chronic pain
Attribute|Clinical Attribute|Hospital Course|12993,12997|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|12993,12997|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12993,12997|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Diagnostic Procedure|Hospital Course|13011,13014|false|false|false|C0013839;C0200204|Electromyogram of eye;Electromyography|EMG
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13018,13026|false|false|false|C0005847|Blood Vessel|Vascular
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13018,13034|false|false|false|C0042381|Vascular Surgical Procedures|Vascular surgery
Finding|Finding|Hospital Course|13027,13034|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Hospital Course|13027,13034|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Hospital Course|13027,13034|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13027,13034|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Conceptual Entity|Hospital Course|13058,13067|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|13058,13067|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|13058,13067|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13058,13067|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Sign or Symptom|Hospital Course|13071,13078|false|false|false|C0030193|Pain|painful
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13080,13085|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13080,13085|false|false|false|C0398102|Procedure on vein|veins
Drug|Biologically Active Substance|Hospital Course|13089,13093|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|13089,13093|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|13089,13093|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|Hospital Course|13089,13093|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|Hospital Course|13089,13104|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|Iron deficiency
Disorder|Disease or Syndrome|Hospital Course|13089,13111|false|false|false|C0162316|Iron deficiency anemia|Iron deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|13094,13104|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|13094,13104|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Hospital Course|13094,13111|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|13105,13111|false|false|false|C0002871|Anemia|anemia
Finding|Functional Concept|Hospital Course|13125,13131|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Drug|Element, Ion, or Isotope|Hospital Course|13132,13139|false|false|false|C0082568|ferryl iron|IV iron
Drug|Biologically Active Substance|Hospital Course|13135,13139|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|13135,13139|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|13135,13139|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|13135,13139|false|false|false|C0337439|Iron measurement|iron
Finding|Functional Concept|Hospital Course|13140,13148|false|false|false|C1827465|Infusion route|infusion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13140,13148|false|false|false|C0574032|Infusion procedures|infusion
Finding|Idea or Concept|Hospital Course|13156,13163|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13164,13167|false|false|false|C5565118|TGM2 protein, human|TTG
Drug|Enzyme|Hospital Course|13164,13167|false|false|false|C5565118|TGM2 protein, human|TTG
Drug|Pharmacologic Substance|Hospital Course|13164,13167|false|false|false|C5565118|TGM2 protein, human|TTG
Finding|Gene or Genome|Hospital Course|13164,13167|false|false|false|C5575307|TGM2 wt Allele|TTG
Drug|Organic Chemical|Hospital Course|13211,13218|false|true|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|13211,13218|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|13211,13218|false|true|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|13222,13226|false|true|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13228,13234|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|13228,13234|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|13228,13234|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13228,13234|false|false|false|C0191838|Procedures on breast|breast
Finding|Pathologic Function|Hospital Course|13228,13243|false|false|false|C0342095|Breast hematoma|breast hematoma
Finding|Pathologic Function|Hospital Course|13235,13243|false|false|false|C0018944|Hematoma|hematoma
Finding|Conceptual Entity|Hospital Course|13248,13255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|13248,13255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|13248,13255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|13248,13258|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|13259,13262|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|13259,13262|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|13259,13262|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13267,13292|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Drug|Immunologic Factor|Hospital Course|13267,13292|false|false|false|C0162595|Antiphospholipid Antibodies|antiphospholipid antibody
Finding|Finding|Hospital Course|13267,13292|false|false|false|C4019436|Antiphospholipid antibody positivity|antiphospholipid antibody
Disorder|Disease or Syndrome|Hospital Course|13267,13301|false|false|false|C0085278|Antiphospholipid Syndrome|antiphospholipid antibody syndrome
Anatomy|Cell Component|Hospital Course|13284,13292|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13284,13292|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Hospital Course|13284,13292|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Hospital Course|13284,13292|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Hospital Course|13284,13292|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Hospital Course|13293,13301|false|false|false|C0039082|Syndrome|syndrome
Finding|Finding|Hospital Course|13304,13322|false|false|false|C1168145|Anticoagulation drug level below therapeutic|subtherapeutic INR
Attribute|Clinical Attribute|Hospital Course|13319,13322|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|13319,13322|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13319,13322|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Body Substance|Hospital Course|13350,13357|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|13350,13357|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|13350,13357|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|13371,13375|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|13371,13375|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|13371,13375|false|false|false|C1553498|home health encounter|home
Drug|Hazardous or Poisonous Substance|Hospital Course|13377,13385|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|13377,13385|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|13377,13385|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|13386,13393|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13386,13393|false|false|false|C0040808|Treatment Protocols|regimen
Attribute|Clinical Attribute|Hospital Course|13396,13407|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|13396,13407|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|13396,13407|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|13396,13420|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|13411,13420|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|13439,13449|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|13439,13449|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|13439,13454|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|13450,13454|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|13471,13479|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|13471,13479|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|13471,13479|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|13471,13479|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|13471,13479|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|13484,13496|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13484,13496|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|13514,13522|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|13514,13522|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|13514,13529|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|13514,13529|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|13523,13529|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13523,13529|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13523,13529|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|13523,13529|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13523,13529|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13540,13543|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13540,13543|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13540,13543|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13540,13543|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13548,13558|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|13548,13558|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13568,13571|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13568,13571|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|13568,13571|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|13568,13571|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|13576,13581|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|13576,13581|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|13599,13609|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|13599,13609|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|13630,13639|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|Hospital Course|13630,13639|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|Hospital Course|13653,13656|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|13657,13662|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|13657,13662|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|Hospital Course|13657,13662|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|13667,13675|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|Hospital Course|13667,13675|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|Hospital Course|13667,13675|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|Hospital Course|13689,13692|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|13693,13697|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|13693,13697|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|13693,13697|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|13700,13708|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|13700,13708|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Idea or Concept|Hospital Course|13712,13718|false|false|false|C0392360|Indication of (contextual qualifier)|Reason
Finding|Idea or Concept|Hospital Course|13712,13722|false|false|false|C0392360|Indication of (contextual qualifier)|Reason for
Finding|Gene or Genome|Hospital Course|13723,13726|false|false|false|C1422467|CIAO3 gene|PRN
Event|Activity|Hospital Course|13727,13736|false|false|false|C1883725|Replicate|duplicate
Finding|Functional Concept|Hospital Course|13727,13736|false|false|false|C0205173;C3539942|Double (qualifier value);Duplicate component (foundation metadata concept)|duplicate
Finding|Intellectual Product|Hospital Course|13727,13736|false|false|false|C0205173;C3539942|Double (qualifier value);Duplicate component (foundation metadata concept)|duplicate
Finding|Functional Concept|Hospital Course|13737,13745|false|false|false|C1547671|Override|override
Drug|Biomedical or Dental Material|Hospital Course|13791,13803|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|13791,13803|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|13791,13810|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|13791,13810|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|13804,13810|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|13804,13810|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Finding|Gene or Genome|Hospital Course|13825,13828|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|13829,13841|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|13851,13855|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|13851,13855|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|13851,13855|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|Hospital Course|13851,13855|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|13860,13866|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|13860,13866|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|13860,13870|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|13860,13870|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|13867,13870|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|13867,13870|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Organic Chemical|Hospital Course|13872,13881|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|13872,13881|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|13872,13889|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|13872,13889|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|13882,13889|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|13882,13889|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|13882,13889|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|Hospital Course|13908,13918|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|13908,13918|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|Hospital Course|13924,13927|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|13933,13946|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|13933,13946|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|13933,13946|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|13962,13965|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|13966,13970|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|13966,13970|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|13966,13970|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|13973,13977|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|13978,13983|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|13978,13983|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|13989,13998|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|13989,13998|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14006,14009|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|14006,14009|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|14006,14009|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|14006,14009|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|14006,14009|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14017,14020|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|14017,14020|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|14017,14020|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|Hospital Course|14017,14020|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|14017,14020|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|14028,14031|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|14032,14037|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|14032,14037|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|14032,14037|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|Hospital Course|14039,14045|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|14051,14058|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|14051,14058|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|14051,14058|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|14051,14060|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|14051,14060|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|14051,14060|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|14051,14060|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|14051,14060|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Antibiotic|Hospital Course|14084,14096|false|false|false|C0014806|erythromycin|Erythromycin
Drug|Organic Chemical|Hospital Course|14084,14096|false|false|false|C0014806|erythromycin|Erythromycin
Finding|Functional Concept|Hospital Course|14102,14107|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|14108,14112|false|false|false|C0028912|Ointments|Oint
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14120,14129|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14125,14129|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|14125,14129|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|14139,14149|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|14139,14149|false|false|false|C0016860|furosemide|Furosemide
Finding|Gene or Genome|Hospital Course|14165,14168|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14169,14172|false|false|false|C0023216;C1140621|Leg;Lower Extremity|Leg
Finding|Pathologic Function|Hospital Course|14169,14181|false|false|false|C0581394|Swelling of lower limb|Leg swelling
Finding|Finding|Hospital Course|14173,14181|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|14173,14181|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Hospital Course|14187,14200|false|false|false|C0012306|hydromorphone|HYDROmorphone
Drug|Pharmacologic Substance|Hospital Course|14187,14200|false|false|false|C0012306|hydromorphone|HYDROmorphone
Drug|Organic Chemical|Hospital Course|14202,14210|false|false|false|C0728755|Dilaudid|Dilaudid
Drug|Pharmacologic Substance|Hospital Course|14202,14210|false|false|false|C0728755|Dilaudid|Dilaudid
Finding|Gene or Genome|Hospital Course|14224,14227|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|14228,14232|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|14228,14232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|14228,14232|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|14235,14241|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|Hospital Course|14235,14241|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Drug|Hazardous or Poisonous Substance|Hospital Course|14247,14255|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|14247,14255|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|14247,14255|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|14269,14273|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Hazardous or Poisonous Substance|Hospital Course|14285,14293|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|14285,14293|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|14285,14293|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|14305,14309|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Finding|Body Substance|Hospital Course|14320,14329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14320,14329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14320,14329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14320,14329|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|14320,14341|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|14330,14341|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|14330,14341|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|14330,14341|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|14347,14357|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|14347,14357|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Organic Chemical|Hospital Course|14377,14387|false|false|false|C0060926|gabapentin|gabapentin
Drug|Pharmacologic Substance|Hospital Course|14377,14387|false|false|false|C0060926|gabapentin|gabapentin
Drug|Biomedical or Dental Material|Hospital Course|14397,14403|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|14407,14415|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|14410,14415|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|14410,14415|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|14422,14427|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Drug|Biomedical or Dental Material|Hospital Course|14445,14451|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|14452,14459|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|14468,14477|false|false|false|C0023660|lidocaine|Lidocaine
Drug|Pharmacologic Substance|Hospital Course|14468,14477|false|false|false|C0023660|lidocaine|Lidocaine
Procedure|Laboratory Procedure|Hospital Course|14468,14477|false|false|false|C0202404|Lidocaine measurement|Lidocaine
Drug|Biomedical or Dental Material|Hospital Course|14481,14486|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|14481,14486|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14489,14493|false|false|false|C4308013|PTCH1 protein, human|PTCH
Finding|Gene or Genome|Hospital Course|14489,14493|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Receptor|Hospital Course|14489,14493|false|false|false|C0694887;C1705339;C1826732;C4308013|PTCH gene;PTCH1 gene;PTCH1 protein, human;PTCH1 wt Allele|PTCH
Finding|Functional Concept|Hospital Course|14501,14506|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Hospital Course|14501,14510|false|false|false|C0524470|Right hip region structure|right hip
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14507,14510|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14507,14510|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Hospital Course|14507,14510|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Hospital Course|14507,14510|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Hospital Course|14507,14510|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Hospital Course|14507,14510|false|false|false|C1292890|Procedure on hip|hip
Drug|Organic Chemical|Hospital Course|14516,14525|false|false|false|C0023660|lidocaine|lidocaine
Drug|Pharmacologic Substance|Hospital Course|14516,14525|false|false|false|C0023660|lidocaine|lidocaine
Procedure|Laboratory Procedure|Hospital Course|14516,14525|false|false|false|C0202404|Lidocaine measurement|lidocaine
Finding|Functional Concept|Hospital Course|14530,14535|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|Apply
Drug|Biomedical or Dental Material|Hospital Course|14564,14569|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|Hospital Course|14564,14569|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Idea or Concept|Hospital Course|14571,14578|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|14587,14595|false|false|false|C0040610|tramadol|TraMADol
Drug|Pharmacologic Substance|Hospital Course|14587,14595|false|false|false|C0040610|tramadol|TraMADol
Procedure|Laboratory Procedure|Hospital Course|14587,14595|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADol
Finding|Gene or Genome|Hospital Course|14609,14612|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|14613,14617|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|14613,14617|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|14613,14617|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|14620,14628|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Finding|Intellectual Product|Hospital Course|14620,14628|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|Moderate
Drug|Organic Chemical|Hospital Course|14634,14642|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|Hospital Course|14634,14642|false|false|false|C0040610|tramadol|tramadol
Procedure|Laboratory Procedure|Hospital Course|14634,14642|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Biomedical or Dental Material|Hospital Course|14651,14657|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|14661,14669|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|14664,14669|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|14664,14669|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Hospital Course|14670,14675|false|false|false|C1720374|Every - dosing instruction fragment|Every
Drug|Biomedical or Dental Material|Hospital Course|14707,14713|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|14714,14721|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|14730,14743|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|14730,14743|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|14730,14743|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|14759,14762|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|14763,14767|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|14763,14767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|14763,14767|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Intellectual Product|Hospital Course|14770,14774|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Finding|Hospital Course|14775,14780|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Hospital Course|14775,14780|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Drug|Organic Chemical|Hospital Course|14787,14796|false|false|false|C0001927|albuterol|Albuterol
Drug|Pharmacologic Substance|Hospital Course|14787,14796|false|false|false|C0001927|albuterol|Albuterol
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14804,14807|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|14804,14807|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|14804,14807|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Finding|Cell Function|Hospital Course|14804,14807|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|14804,14807|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14815,14818|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|14815,14818|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|14815,14818|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Finding|Cell Function|Hospital Course|14815,14818|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|14815,14818|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|14826,14829|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|14830,14835|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|14830,14835|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|14830,14835|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|Hospital Course|14837,14843|false|false|false|C0043144|Wheezing|wheeze
Drug|Organic Chemical|Hospital Course|14850,14862|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|14850,14862|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|14882,14890|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|14882,14890|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|14882,14897|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|14882,14897|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|14891,14897|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|14891,14897|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|14891,14897|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|14891,14897|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|14891,14897|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14908,14911|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14908,14911|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|14908,14911|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|14908,14911|false|false|false|C1332410|BID gene|BID
Drug|Antibiotic|Hospital Course|14918,14930|false|false|false|C0014806|erythromycin|Erythromycin
Drug|Organic Chemical|Hospital Course|14918,14930|false|false|false|C0014806|erythromycin|Erythromycin
Finding|Functional Concept|Hospital Course|14936,14941|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|14942,14946|false|false|false|C0028912|Ointments|Oint
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14954,14963|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14959,14963|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|14959,14963|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|14974,14984|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|14974,14984|false|false|false|C0016860|furosemide|Furosemide
Finding|Gene or Genome|Hospital Course|15000,15003|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|15004,15007|false|false|false|C0023216;C1140621|Leg;Lower Extremity|Leg
Finding|Pathologic Function|Hospital Course|15004,15016|false|false|false|C0581394|Swelling of lower limb|Leg swelling
Finding|Finding|Hospital Course|15008,15016|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|15008,15016|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Drug|Organic Chemical|Hospital Course|15024,15034|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|15024,15034|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|Hospital Course|15044,15047|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|15044,15047|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|15044,15047|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|15044,15047|false|false|false|C1332410|BID gene|BID
Drug|Biomedical or Dental Material|Hospital Course|15055,15067|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|15055,15067|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|15055,15074|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|15055,15074|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|15068,15074|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|15068,15074|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Finding|Gene or Genome|Hospital Course|15089,15092|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|15093,15105|false|false|false|C0009806|Constipation|Constipation
Drug|Biologically Active Substance|Hospital Course|15115,15119|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|15115,15119|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Drug|Substance|Hospital Course|15115,15119|false|false|false|C1517938;C1550648|Line Specimen;Long Interspersed Elements|Line
Finding|Intellectual Product|Hospital Course|15115,15119|false|false|false|C1546701|line source specimen code|Line
Drug|Organic Chemical|Hospital Course|15127,15133|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Pharmacologic Substance|Hospital Course|15127,15133|false|false|false|C0162684;C1739179|Pro-Air Procaterol;ProAir|ProAir
Drug|Organic Chemical|Hospital Course|15127,15137|false|false|false|C1739179|ProAir|ProAir HFA
Drug|Pharmacologic Substance|Hospital Course|15127,15137|false|false|false|C1739179|ProAir|ProAir HFA
Disorder|Disease or Syndrome|Hospital Course|15134,15137|false|false|false|C0015458|Facial Hemiatrophy|HFA
Procedure|Diagnostic Procedure|Hospital Course|15134,15137|false|false|false|C0430649|High frequency audiometry|HFA
Drug|Organic Chemical|Hospital Course|15139,15148|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|15139,15148|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|Hospital Course|15139,15156|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|15139,15156|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|15149,15156|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|15149,15156|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|15149,15156|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|Hospital Course|15175,15185|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|15175,15185|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|Hospital Course|15191,15194|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|15202,15207|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|15202,15207|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|15228,15238|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|Hospital Course|15228,15238|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|Hospital Course|15262,15271|false|false|false|C0040805|trazodone|TraZODone
Drug|Pharmacologic Substance|Hospital Course|15262,15271|false|false|false|C0040805|trazodone|TraZODone
Finding|Gene or Genome|Hospital Course|15285,15288|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|15289,15294|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|15289,15294|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|Hospital Course|15289,15294|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|15302,15309|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|15302,15309|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|15302,15309|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|15302,15311|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|15302,15311|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|15302,15311|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|15302,15311|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|15302,15311|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Hazardous or Poisonous Substance|Hospital Course|15337,15345|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|15337,15345|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|15337,15345|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|15357,15361|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Drug|Hazardous or Poisonous Substance|Hospital Course|15375,15383|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|15375,15383|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|15375,15383|false|false|false|C0043031|warfarin|Warfarin
Finding|Intellectual Product|Hospital Course|15397,15401|false|false|false|C1561540|Transaction counts and value totals - week|WEEK
Finding|Body Substance|Hospital Course|15413,15422|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|15413,15422|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|15413,15422|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|15413,15422|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|15413,15434|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|15413,15434|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|15423,15434|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|15423,15434|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|15436,15440|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|15436,15440|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|15436,15440|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|15446,15453|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|15446,15453|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|Hospital Course|15456,15464|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|15472,15481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|15472,15481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|15472,15481|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|15472,15481|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|15472,15491|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|15482,15491|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|15482,15491|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|15482,15491|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|15482,15491|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Functional Concept|Hospital Course|15520,15525|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|15520,15547|false|false|false|C3862456|right trochanteric bursitis|Right trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|15526,15547|false|false|false|C0151451|Greater trochanteric pain syndrome|trochanteric bursitis
Disorder|Disease or Syndrome|Hospital Course|15539,15547|false|false|false|C0006444|Bursitis|bursitis
Finding|Functional Concept|Hospital Course|15548,15553|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|15554,15562|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|15563,15566|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|15563,15571|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Hospital Course|15567,15571|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|15567,15571|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|15567,15571|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|15572,15577|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Disorder|Disease or Syndrome|Hospital Course|15584,15598|false|false|false|C0042345|Varicosity|varicose veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|15593,15598|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15593,15598|false|false|false|C0398102|Procedure on vein|veins
Disorder|Neoplastic Process|Hospital Course|15601,15610|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Finding|Functional Concept|Hospital Course|15601,15610|false|false|false|C1522484|metastatic qualifier|SECONDARY
Drug|Biologically Active Substance|Hospital Course|15630,15634|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|15630,15634|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|15630,15634|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|Hospital Course|15630,15634|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|Hospital Course|15630,15645|false|false|false|C0162316;C0240066|Iron deficiency;Iron deficiency anemia|Iron deficiency
Disorder|Disease or Syndrome|Hospital Course|15630,15652|false|false|false|C0162316|Iron deficiency anemia|Iron deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|15635,15645|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|15635,15645|false|false|false|C0011155|Deficiency|deficiency
Disorder|Disease or Syndrome|Hospital Course|15635,15652|false|false|false|C0041782|Deficiency anemias|deficiency anemia
Disorder|Disease or Syndrome|Hospital Course|15646,15652|false|false|false|C0002871|Anemia|anemia
Finding|Conceptual Entity|Hospital Course|15653,15660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|15653,15660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|Hospital Course|15653,15660|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|Hospital Course|15653,15663|false|false|false|C0262926|Medical History|History of
Anatomy|Body Location or Region|Hospital Course|15664,15667|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|15664,15667|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|15664,15667|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15671,15682|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|15674,15682|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|15674,15682|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|15674,15682|false|false|false|C0043031|warfarin|warfarin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|15683,15708|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Drug|Immunologic Factor|Hospital Course|15683,15708|false|false|false|C0162595|Antiphospholipid Antibodies|Antiphospholipid antibody
Finding|Finding|Hospital Course|15683,15708|false|false|false|C4019436|Antiphospholipid antibody positivity|Antiphospholipid antibody
Disorder|Disease or Syndrome|Hospital Course|15683,15717|false|false|false|C0085278|Antiphospholipid Syndrome|Antiphospholipid antibody syndrome
Anatomy|Cell Component|Hospital Course|15700,15708|false|false|false|C1167408;C3665580|Immunoglobulin complex location, circulating;immunoglobulin complex location|antibody
Drug|Amino Acid, Peptide, or Protein|Hospital Course|15700,15708|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Immunologic Factor|Hospital Course|15700,15708|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Drug|Pharmacologic Substance|Hospital Course|15700,15708|false|false|false|C0003241;C0021027|Antibodies;Immunoglobulins|antibody
Procedure|Laboratory Procedure|Hospital Course|15700,15708|false|false|false|C4551530|Antibody (immunoassay)|antibody
Disorder|Disease or Syndrome|Hospital Course|15709,15717|false|false|false|C0039082|Syndrome|syndrome
Finding|Finding|Hospital Course|15718,15736|false|false|false|C1168145|Anticoagulation drug level below therapeutic|Subtherapeutic INR
Attribute|Clinical Attribute|Hospital Course|15733,15736|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|15733,15736|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|15733,15736|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|Hospital Course|15737,15744|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|15737,15744|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|15737,15744|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|15737,15746|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|15737,15746|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|15737,15746|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|15737,15746|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|15737,15746|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Disorder|Disease or Syndrome|Hospital Course|15737,15757|false|false|false|C0042870|Vitamin D Deficiency|Vitamin D deficiency
Finding|Finding|Hospital Course|15737,15757|false|false|false|C5886864|Decreased circulating vitamin D concentration|Vitamin D deficiency
Disorder|Disease or Syndrome|Hospital Course|15747,15757|false|false|false|C0162429|Malnutrition|deficiency
Finding|Functional Concept|Hospital Course|15747,15757|false|false|false|C0011155|Deficiency|deficiency
Finding|Mental Process|Discharge Condition|15782,15788|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|15782,15795|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|15782,15795|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|15789,15795|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|15789,15795|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|15797,15802|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|15807,15815|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|15817,15839|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|15817,15839|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|15826,15839|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|15826,15839|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|15841,15846|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|15841,15846|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|15841,15846|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|15841,15846|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|15841,15846|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|15841,15846|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|15851,15862|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|15864,15872|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|15864,15872|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|15864,15872|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|15873,15879|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|15873,15879|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|15881,15891|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|15881,15891|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|15881,15891|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|15881,15891|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Social Behavior|Discharge Condition|15903,15913|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|15917,15920|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|15917,15920|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|Discharge Condition|15917,15920|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|15917,15920|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Gene or Genome|Discharge Instructions|15967,15971|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Finding|Discharge Instructions|16021,16026|false|false|false|C2984081|Very Much|a lot
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16023,16026|false|false|false|C0162435;C0175218|Olfactory tract;nucleus of the lateral olfactory tract|lot
Finding|Idea or Concept|Discharge Instructions|16023,16026|false|false|false|C1710198|Stock (in-store merchandise)|lot
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16030,16033|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Discharge Instructions|16030,16038|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Discharge Instructions|16034,16038|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|16034,16038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|16034,16038|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|16051,16060|false|false|false|C0332218|Difficult (qualifier value)|difficult
Finding|Idea or Concept|Discharge Instructions|16079,16087|false|false|false|C1547192|Organization unit type - Hospital|hospital
Drug|Organic Chemical|Discharge Instructions|16103,16110|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Discharge Instructions|16103,16110|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16103,16120|false|false|false|C1261311|Injection of steroid|steroid injection
Drug|Biomedical or Dental Material|Discharge Instructions|16111,16120|false|false|false|C1272883|Injection|injection
Finding|Functional Concept|Discharge Instructions|16111,16120|false|false|false|C1828121|Injection Route of Administration|injection
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16111,16120|false|false|false|C0021485;C1533685|Injection of therapeutic agent;Injection procedure|injection
Finding|Functional Concept|Discharge Instructions|16131,16136|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|Discharge Instructions|16138,16143|false|false|false|C0039866;C4299091|Lower extremity>Thigh;Thigh structure|thigh
Attribute|Clinical Attribute|Discharge Instructions|16150,16159|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|16150,16159|false|false|false|C0012634|Disease|condition
Finding|Conceptual Entity|Discharge Instructions|16150,16159|false|false|false|C1705253|Logical Condition|condition
Disorder|Disease or Syndrome|Discharge Instructions|16168,16189|false|false|false|C0151451|Greater trochanteric pain syndrome|Trochanteric Bursitis
Disorder|Disease or Syndrome|Discharge Instructions|16181,16189|false|false|false|C0006444|Bursitis|Bursitis
Drug|Pharmacologic Substance|Discharge Instructions|16211,16221|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|16211,16221|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|16229,16239|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Discharge Instructions|16229,16239|false|false|false|C0060926|gabapentin|Gabapentin
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16258,16261|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Attribute|Clinical Attribute|Discharge Instructions|16263,16267|false|true|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|16263,16267|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|16263,16267|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|Discharge Instructions|16268,16273|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Discharge Instructions|16268,16273|false|false|false|C2003888|Lower (action)|lower
Drug|Pharmacologic Substance|Discharge Instructions|16307,16317|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|16307,16317|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|16325,16332|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Discharge Instructions|16325,16332|false|false|false|C0728963|Lovenox|Lovenox
Event|Activity|Discharge Instructions|16336,16341|false|false|false|C1705178|Order (action)|order
Finding|Classification|Discharge Instructions|16336,16341|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Idea or Concept|Discharge Instructions|16336,16341|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Finding|Intellectual Product|Discharge Instructions|16336,16341|false|false|false|C1546465;C1705175;C1705177;C4284072;C5444833|Medical Order;Order (document);Order (record artifact);Order (taxonomic);What subject filter - Order|order
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|16336,16341|false|false|false|C1373200|Order [PK]|order
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16346,16352|false|false|false|C0399080|Fixation of dental bridge|bridge
Drug|Hazardous or Poisonous Substance|Discharge Instructions|16370,16378|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Discharge Instructions|16370,16378|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Discharge Instructions|16370,16378|false|false|false|C0043031|warfarin|warfarin
Drug|Hazardous or Poisonous Substance|Discharge Instructions|16397,16405|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Discharge Instructions|16397,16405|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Discharge Instructions|16397,16405|false|false|false|C0043031|warfarin|warfarin
Attribute|Clinical Attribute|Discharge Instructions|16397,16410|false|false|false|C4082242||warfarin dose
Procedure|Laboratory Procedure|Discharge Instructions|16397,16410|false|false|false|C0366686|warfarin dose|warfarin dose
Attribute|Clinical Attribute|Discharge Instructions|16437,16440|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Discharge Instructions|16437,16440|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|16437,16440|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Body Substance|Discharge Instructions|16452,16461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|16452,16461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|16452,16461|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|16452,16461|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Discharge Instructions|16463,16467|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Discharge Instructions|16463,16467|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Functional Concept|Discharge Instructions|16507,16518|false|false|false|C1522726|Intravenous Route of Administration|intravenous
Drug|Biologically Active Substance|Discharge Instructions|16519,16523|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Discharge Instructions|16519,16523|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Discharge Instructions|16519,16523|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Discharge Instructions|16519,16523|false|false|false|C0337439|Iron measurement|iron
Drug|Biologically Active Substance|Discharge Instructions|16541,16545|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Discharge Instructions|16541,16545|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Discharge Instructions|16541,16545|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Discharge Instructions|16541,16545|false|false|false|C0337439|Iron measurement|iron
Finding|Functional Concept|Discharge Instructions|16546,16555|false|false|false|C0011155|Deficiency|deficient
Finding|Sign or Symptom|Discharge Instructions|16586,16594|false|false|false|C0015672|Fatigue|fatigued
Finding|Idea or Concept|Discharge Instructions|16621,16625|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|16621,16625|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|16621,16625|false|false|false|C1553498|home health encounter|home
Attribute|Clinical Attribute|Discharge Instructions|16644,16655|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|16644,16655|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|16644,16655|false|false|false|C4284232|Medications|medications
Event|Activity|Discharge Instructions|16683,16694|false|false|false|C0003629|Appointments|appointment
Finding|Intellectual Product|Discharge Instructions|16705,16717|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|16705,16717|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Discharge Instructions|16713,16717|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|16713,16717|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|16713,16717|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|16718,16724|false|false|false|C2348314|Doctor - Title|doctor
Anatomy|Body Location or Region|Discharge Instructions|16770,16775|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Discharge Instructions|16770,16775|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16770,16779|false|false|false|C1140621;C4299093|Leg;Lower extremity>Lower leg|lower leg
Finding|Sign or Symptom|Discharge Instructions|16770,16784|false|true|false|C0023222;C0839480|Pain in limb, lower leg;Pain in lower limb|lower leg pain
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16776,16779|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Discharge Instructions|16776,16784|false|true|false|C0023222|Pain in lower limb|leg pain
Attribute|Clinical Attribute|Discharge Instructions|16780,16784|false|true|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|16780,16784|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|16780,16784|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|16806,16810|false|false|true|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Finding|Individual Behavior|Discharge Instructions|16806,16810|false|false|true|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Finding|Organism Function|Discharge Instructions|16806,16810|false|false|true|C0037817;C0234856;C0600118|Does talk;Speaking (function);Speech|talk
Finding|Individual Behavior|Discharge Instructions|16806,16825|false|false|true|C1456713|Talking With Your Doctor|talk to your doctor
Finding|Intellectual Product|Discharge Instructions|16819,16825|false|false|true|C2348314|Doctor - Title|doctor
Finding|Gene or Genome|Discharge Instructions|16842,16845|false|false|true|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Discharge Instructions|16842,16845|false|false|true|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Discharge Instructions|16842,16845|false|false|true|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16854,16859|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|Discharge Instructions|16854,16859|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|Discharge Instructions|16854,16859|false|false|true|C0150920|Spine Problem|spine
Finding|Intellectual Product|Discharge Instructions|16884,16890|false|false|true|C2348314|Doctor - Title|doctor
Drug|Pharmacologic Substance|Discharge Instructions|16911,16921|false|false|true|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|16911,16921|false|false|true|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Drug|Organic Chemical|Discharge Instructions|16930,16940|false|false|false|C0012091|diclofenac|DICLOFENAC
Drug|Pharmacologic Substance|Discharge Instructions|16930,16940|false|false|false|C0012091|diclofenac|DICLOFENAC
Drug|Biomedical or Dental Material|Discharge Instructions|16941,16944|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|GEL
Drug|Indicator, Reagent, or Diagnostic Aid|Discharge Instructions|16941,16944|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|GEL
Drug|Substance|Discharge Instructions|16941,16944|false|false|false|C0017243;C0972569;C1382104;C1551386|Electrophoresis Gel;Gel;Gel - ContainerSeparator;Gel physical state|GEL
Procedure|Laboratory Procedure|Discharge Instructions|16941,16944|false|false|false|C5977403|Blood group antibody screen.GEL|GEL
Drug|Organic Chemical|Discharge Instructions|16958,16966|false|false|false|C0699958|Voltaren|VOLTAREN
Drug|Pharmacologic Substance|Discharge Instructions|16958,16966|false|false|false|C0699958|Voltaren|VOLTAREN
Drug|Organic Chemical|Discharge Instructions|16988,16994|false|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|Discharge Instructions|16988,16994|false|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|Discharge Instructions|16999,17004|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|Discharge Instructions|16999,17004|false|false|false|C0593507|Advil|Advil
Finding|Gene or Genome|Discharge Instructions|16999,17004|false|false|false|C1422473|AVIL gene|Advil
Drug|Biomedical or Dental Material|Discharge Instructions|17010,17017|false|false|false|C1710439|Topical Dosage Form|topical
Finding|Functional Concept|Discharge Instructions|17010,17017|false|false|false|C1522168|Topical Route of Administration|topical
Attribute|Clinical Attribute|Discharge Instructions|17018,17022|false|false|false|C4255237||form
Finding|Functional Concept|Discharge Instructions|17018,17022|false|false|false|C1522492|Formation|form
Attribute|Clinical Attribute|Discharge Instructions|17041,17045|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|17041,17045|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|17041,17045|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|Discharge Instructions|17082,17088|false|false|false|C2348314|Doctor - Title|doctor
Drug|Biologically Active Substance|Discharge Instructions|17111,17115|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Discharge Instructions|17111,17115|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Discharge Instructions|17111,17115|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Discharge Instructions|17111,17115|false|false|false|C0337439|Iron measurement|iron
Finding|Functional Concept|Discharge Instructions|17116,17125|false|false|false|C0011155|Deficiency|deficient
Finding|Intellectual Product|Discharge Instructions|17138,17146|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|17138,17146|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Idea or Concept|Discharge Instructions|17154,17158|false|false|false|C1552020|Role Class - part|part
Event|Activity|Discharge Instructions|17167,17171|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|17167,17171|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|17167,17171|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Disorder|Disease or Syndrome|Discharge Instructions|17194,17198|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Discharge Instructions|17194,17198|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Finding|Idea or Concept|Discharge Instructions|17209,17215|false|false|false|C0018684|Health|health
Procedure|Health Care Activity|Discharge Instructions|17248,17256|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|17257,17269|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|17257,17269|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

