 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
UROLOGY|153,160
<EOL>|160,161
<EOL>|162,163
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
Abdominal|256,265
pain|266,270
,|270,271
distention|272,282
,|282,283
nausea|284,290
<EOL>|290,291
<EOL>|292,293
Major|293,298
Surgical|299,307
or|308,310
Invasive|311,319
Procedure|320,329
:|329,330
<EOL>|330,331
Interventional|331,345
radiology|346,355
placement|356,365
of|366,368
abdominal|369,378
abscess|379,386
drain|387,392
<EOL>|392,393
<EOL>|393,394
<EOL>|395,396
_|424,425
_|425,426
_|426,427
F|428,429
with|430,434
h|435,436
/|436,437
o|437,438
muscle|439,445
invasive|446,454
bladder|455,462
cancer|463,469
,|469,470
returning|471,480
to|481,483
<EOL>|484,485
the|485,488
ED|489,491
POD|492,495
15|496,498
with|499,503
abdominal|504,513
pain|514,518
,|518,519
nausea|520,526
,|526,527
and|528,531
distension|532,542
.|542,543
She|544,547
<EOL>|548,549
has|549,552
been|553,557
obstipated|558,568
for|569,572
nearly|573,579
three|580,585
days|586,590
.|590,591
KUB|592,595
and|596,599
CT|600,602
scan|603,607
<EOL>|608,609
notable|609,616
for|617,620
dilated|621,628
loops|629,634
,|634,635
air|636,639
fluids|640,646
,|646,647
and|648,651
tapering|652,660
small|661,666
bowel|667,672
<EOL>|673,674
without|674,681
an|682,684
obvious|685,692
transition|693,703
point|704,709
.|709,710
Labwork|711,718
notable|719,726
for|727,730
_|731,732
_|732,733
_|733,734
<EOL>|735,736
and|736,739
<EOL>|739,740
leukocytosis|740,752
.|752,753
Concerned|754,763
for|764,767
small|768,773
bowel|774,779
obstruction|780,791
or|792,794
an|795,797
ileus|798,803
<EOL>|804,805
in|805,807
presence|808,816
_|817,818
_|818,819
_|819,820
and|821,824
leukocytosis|825,837
she|838,841
was|842,845
re-admitted|846,857
for|858,861
IVF|862,865
,|865,866
<EOL>|867,868
bowel|868,873
rest|874,878
,|878,879
NGT|880,883
decompression|884,897
.|897,898
<EOL>|899,900
<EOL>|901,902
Hypertension|924,936
,|936,937
laparoscopic|938,950
cholecystectomy|951,966
,|966,967
left|968,972
knee|973,977
<EOL>|978,979
replacement|979,990
six|991,994
to|995,997
_|998,999
_|999,1000
_|1000,1001
years|1002,1007
ago|1008,1011
,|1011,1012
laminectomy|1013,1024
of|1025,1027
L5|1028,1030
-|1030,1031
S1|1031,1033
at|1034,1036
age|1037,1040
<EOL>|1041,1042
_|1042,1043
_|1043,1044
_|1044,1045
,|1045,1046
two|1047,1050
vaginal|1051,1058
deliveries|1059,1069
.|1069,1070
<EOL>|1070,1071
<EOL>|1071,1072
s|1072,1073
/|1073,1074
p|1074,1075
_|1076,1077
_|1077,1078
_|1078,1079
:|1079,1080
<EOL>|1081,1082
1.|1082,1084
Robot|1086,1091
-|1091,1092
assisted|1092,1100
laparoscopic|1101,1113
bilateral|1114,1123
pelvic|1124,1130
lymph|1131,1136
node|1137,1141
<EOL>|1142,1143
dissection|1143,1153
.|1153,1154
<EOL>|1154,1155
2.|1155,1157
Robot|1158,1163
-|1163,1164
assisted|1164,1172
hysterectomy|1173,1185
and|1186,1189
bilateral|1190,1199
oophorectomy|1200,1212
for|1213,1216
<EOL>|1217,1218
large|1218,1223
uterus|1224,1230
,|1230,1231
greater|1232,1239
than|1240,1244
300|1245,1248
grams|1249,1254
,|1254,1255
with|1256,1260
large|1261,1266
fibroid|1267,1274
.|1274,1275
<EOL>|1275,1276
3.|1276,1278
Laparoscopic|1279,1291
radical|1292,1299
cystectomy|1300,1310
and|1311,1314
anterior|1315,1323
vaginectomy|1324,1335
with|1336,1340
<EOL>|1341,1342
vaginal|1342,1349
reconstruction|1350,1364
.|1364,1365
<EOL>|1365,1366
<EOL>|1366,1367
<EOL>|1368,1369
:|1383,1384
<EOL>|1384,1385
_|1385,1386
_|1386,1387
_|1387,1388
<EOL>|1388,1389
:|1403,1404
<EOL>|1404,1405
Negative|1405,1413
for|1414,1417
bladder|1418,1425
CA|1426,1428
.|1428,1429
<EOL>|1429,1430
<EOL>|1430,1431
<EOL>|1432,1433
WdWn|1448,1452
,|1452,1453
NAD|1454,1457
,|1457,1458
AVSS|1459,1463
<EOL>|1463,1464
Abdomen|1464,1471
soft|1472,1476
,|1476,1477
appropriately|1478,1491
tender|1492,1498
along|1499,1504
incision|1505,1513
<EOL>|1513,1514
Incision|1514,1522
is|1523,1525
c|1526,1527
/|1527,1528
d|1528,1529
/|1529,1530
I|1530,1531
<EOL>|1531,1532
Stoma|1532,1537
is|1538,1540
well|1541,1545
perfused|1546,1554
;|1554,1555
Urine|1556,1561
color|1562,1567
is|1568,1570
yellow|1571,1577
<EOL>|1577,1578
Bilateral|1578,1587
lower|1588,1593
extremities|1594,1605
are|1606,1609
warm|1610,1614
,|1614,1615
dry|1616,1619
,|1619,1620
well|1621,1625
perfused|1626,1634
.|1634,1635
There|1637,1642
<EOL>|1643,1644
is|1644,1646
no|1647,1649
reported|1650,1658
calf|1659,1663
pain|1664,1668
to|1669,1671
deep|1672,1676
palpation|1677,1686
.|1686,1687
Bilateral|1688,1697
lower|1698,1703
<EOL>|1704,1705
extremities|1705,1716
have|1717,1721
2|1722,1723
+|1723,1724
pitting|1725,1732
edema|1733,1738
but|1739,1742
no|1743,1745
erythema|1746,1754
,|1754,1755
callor|1756,1762
,|1762,1763
pain|1764,1768
.|1768,1769
<EOL>|1770,1771
<EOL>|1771,1772
Pigtail|1772,1779
drain|1780,1785
has|1786,1789
been|1790,1794
removed|1795,1802
-|1803,1804
dressing|1805,1813
c|1814,1815
/|1815,1816
d|1816,1817
/|1817,1818
i|1818,1819
<EOL>|1819,1820
<EOL>|1821,1822
Pertinent|1822,1831
Results|1832,1839
:|1839,1840
<EOL>|1840,1841
_|1841,1842
_|1842,1843
_|1843,1844
05|1845,1847
:|1847,1848
58AM|1848,1852
BLOOD|1853,1858
WBC|1859,1862
-|1862,1863
9.9|1863,1866
RBC|1867,1870
-|1870,1871
2|1871,1872
.|1872,1873
76|1873,1875
*|1875,1876
Hgb|1877,1880
-|1880,1881
8|1881,1882
.|1882,1883
2|1883,1884
*|1884,1885
Hct|1886,1889
-|1889,1890
26|1890,1892
.|1892,1893
2|1893,1894
*|1894,1895
<EOL>|1896,1897
MCV|1897,1900
-|1900,1901
95|1901,1903
MCH|1904,1907
-|1907,1908
29.7|1908,1912
MCHC|1913,1917
-|1917,1918
31|1918,1920
.|1920,1921
3|1921,1922
*|1922,1923
RDW|1924,1927
-|1927,1928
13.9|1928,1932
RDWSD|1933,1938
-|1938,1939
47|1939,1941
.|1941,1942
3|1942,1943
*|1943,1944
Plt|1945,1948
_|1949,1950
_|1950,1951
_|1951,1952
<EOL>|1952,1953
_|1953,1954
_|1954,1955
_|1955,1956
06|1957,1959
:|1959,1960
45AM|1960,1964
BLOOD|1965,1970
WBC|1971,1974
-|1974,1975
10|1975,1977
.|1977,1978
3|1978,1979
*|1979,1980
RBC|1981,1984
-|1984,1985
2|1985,1986
.|1986,1987
87|1987,1989
*|1989,1990
Hgb|1991,1994
-|1994,1995
8|1995,1996
.|1996,1997
7|1997,1998
*|1998,1999
Hct|2000,2003
-|2003,2004
27|2004,2006
.|2006,2007
7|2007,2008
*|2008,2009
<EOL>|2010,2011
MCV|2011,2014
-|2014,2015
97|2015,2017
MCH|2018,2021
-|2021,2022
30.3|2022,2026
MCHC|2027,2031
-|2031,2032
31|2032,2034
.|2034,2035
4|2035,2036
*|2036,2037
RDW|2038,2041
-|2041,2042
14.0|2042,2046
RDWSD|2047,2052
-|2052,2053
49|2053,2055
.|2055,2056
4|2056,2057
*|2057,2058
Plt|2059,2062
_|2063,2064
_|2064,2065
_|2065,2066
<EOL>|2066,2067
_|2067,2068
_|2068,2069
_|2069,2070
05|2071,2073
:|2073,2074
13AM|2074,2078
BLOOD|2079,2084
WBC|2085,2088
-|2088,2089
11|2089,2091
.|2091,2092
6|2092,2093
*|2093,2094
RBC|2095,2098
-|2098,2099
3|2099,2100
.|2100,2101
27|2101,2103
*|2103,2104
Hgb|2105,2108
-|2108,2109
9|2109,2110
.|2110,2111
8|2111,2112
*|2112,2113
Hct|2114,2117
-|2117,2118
31|2118,2120
.|2120,2121
0|2121,2122
*|2122,2123
<EOL>|2124,2125
MCV|2125,2128
-|2128,2129
95|2129,2131
MCH|2132,2135
-|2135,2136
30.0|2136,2140
MCHC|2141,2145
-|2145,2146
31|2146,2148
.|2148,2149
6|2149,2150
*|2150,2151
RDW|2152,2155
-|2155,2156
13.6|2156,2160
RDWSD|2161,2166
-|2166,2167
47|2167,2169
.|2169,2170
5|2170,2171
*|2171,2172
Plt|2173,2176
_|2177,2178
_|2178,2179
_|2179,2180
<EOL>|2180,2181
_|2181,2182
_|2182,2183
_|2183,2184
07|2185,2187
:|2187,2188
06PM|2188,2192
BLOOD|2193,2198
WBC|2199,2202
-|2202,2203
22|2203,2205
.|2205,2206
5|2206,2207
*|2207,2208
#|2208,2209
RBC|2210,2213
-|2213,2214
3|2214,2215
.|2215,2216
58|2216,2218
*|2218,2219
Hgb|2220,2223
-|2223,2224
10|2224,2226
.|2226,2227
9|2227,2228
*|2228,2229
Hct|2230,2233
-|2233,2234
34.0|2234,2238
<EOL>|2239,2240
MCV|2240,2243
-|2243,2244
95|2244,2246
MCH|2247,2250
-|2250,2251
30.4|2251,2255
MCHC|2256,2260
-|2260,2261
32.1|2261,2265
RDW|2266,2269
-|2269,2270
13.9|2270,2274
RDWSD|2275,2280
-|2280,2281
47|2281,2283
.|2283,2284
9|2284,2285
*|2285,2286
Plt|2287,2290
_|2291,2292
_|2292,2293
_|2293,2294
<EOL>|2294,2295
_|2295,2296
_|2296,2297
_|2297,2298
07|2299,2301
:|2301,2302
06PM|2302,2306
BLOOD|2307,2312
Neuts|2313,2318
-|2318,2319
89|2319,2321
*|2321,2322
Bands|2323,2328
-|2328,2329
1|2329,2330
Lymphs|2331,2337
-|2337,2338
5|2338,2339
*|2339,2340
Monos|2341,2346
-|2346,2347
3|2347,2348
*|2348,2349
<EOL>|2350,2351
Eos|2351,2354
-|2354,2355
0|2355,2356
Baso|2357,2361
-|2361,2362
0|2362,2363
_|2364,2365
_|2365,2366
_|2366,2367
Metas|2368,2373
-|2373,2374
1|2374,2375
*|2375,2376
Myelos|2377,2383
-|2383,2384
0|2384,2385
Hyperse|2386,2393
-|2393,2394
1|2394,2395
*|2395,2396
AbsNeut|2397,2404
-|2404,2405
20|2405,2407
.|2407,2408
48|2408,2410
*|2410,2411
<EOL>|2412,2413
AbsLymp|2413,2420
-|2420,2421
1|2421,2422
.|2422,2423
13|2423,2425
*|2425,2426
AbsMono|2427,2434
-|2434,2435
0|2435,2436
.|2436,2437
68|2437,2439
AbsEos|2440,2446
-|2446,2447
0|2447,2448
.|2448,2449
00|2449,2451
*|2451,2452
AbsBaso|2453,2460
-|2460,2461
0|2461,2462
.|2462,2463
00|2463,2465
*|2465,2466
<EOL>|2466,2467
_|2467,2468
_|2468,2469
_|2469,2470
01|2471,2473
:|2473,2474
04PM|2474,2478
BLOOD|2479,2484
_|2485,2486
_|2486,2487
_|2487,2488
PTT|2489,2492
-|2492,2493
30.9|2493,2497
_|2498,2499
_|2499,2500
_|2500,2501
<EOL>|2501,2502
_|2502,2503
_|2503,2504
_|2504,2505
05|2506,2508
:|2508,2509
58AM|2509,2513
BLOOD|2514,2519
Glucose|2520,2527
-|2527,2528
106|2528,2531
*|2531,2532
UreaN|2533,2538
-|2538,2539
26|2539,2541
*|2541,2542
Creat|2543,2548
-|2548,2549
0.4|2549,2552
Na|2553,2555
-|2555,2556
136|2556,2559
<EOL>|2560,2561
K|2561,2562
-|2562,2563
4.6|2563,2566
Cl|2567,2569
-|2569,2570
107|2570,2573
HCO3|2574,2578
-|2578,2579
26|2579,2581
AnGap|2582,2587
-|2587,2588
8|2588,2589
<EOL>|2589,2590
_|2590,2591
_|2591,2592
_|2592,2593
06|2594,2596
:|2596,2597
45AM|2597,2601
BLOOD|2602,2607
Glucose|2608,2615
-|2615,2616
114|2616,2619
*|2619,2620
UreaN|2621,2626
-|2626,2627
32|2627,2629
*|2629,2630
Creat|2631,2636
-|2636,2637
0.4|2637,2640
Na|2641,2643
-|2643,2644
137|2644,2647
<EOL>|2648,2649
K|2649,2650
-|2650,2651
4.1|2651,2654
Cl|2655,2657
-|2657,2658
106|2658,2661
HCO3|2662,2666
-|2666,2667
25|2667,2669
AnGap|2670,2675
-|2675,2676
10|2676,2678
<EOL>|2678,2679
_|2679,2680
_|2680,2681
_|2681,2682
06|2683,2685
:|2685,2686
00AM|2686,2690
BLOOD|2691,2696
Glucose|2697,2704
-|2704,2705
121|2705,2708
*|2708,2709
UreaN|2710,2715
-|2715,2716
39|2716,2718
*|2718,2719
Creat|2720,2725
-|2725,2726
0.4|2726,2729
Na|2730,2732
-|2732,2733
140|2733,2736
<EOL>|2737,2738
K|2738,2739
-|2739,2740
3.6|2740,2743
Cl|2744,2746
-|2746,2747
107|2747,2750
HCO3|2751,2755
-|2755,2756
26|2756,2758
AnGap|2759,2764
-|2764,2765
11|2765,2767
<EOL>|2767,2768
_|2768,2769
_|2769,2770
_|2770,2771
07|2772,2774
:|2774,2775
06PM|2775,2779
BLOOD|2780,2785
Glucose|2786,2793
-|2793,2794
117|2794,2797
*|2797,2798
UreaN|2799,2804
-|2804,2805
60|2805,2807
*|2807,2808
Creat|2809,2814
-|2814,2815
1|2815,2816
.|2816,2817
7|2817,2818
*|2818,2819
#|2819,2820
Na|2821,2823
-|2823,2824
133|2824,2827
<EOL>|2828,2829
K|2829,2830
-|2830,2831
5.0|2831,2834
Cl|2835,2837
-|2837,2838
96|2838,2840
HCO3|2841,2845
-|2845,2846
21|2846,2848
*|2848,2849
AnGap|2850,2855
-|2855,2856
21|2856,2858
*|2858,2859
<EOL>|2859,2860
_|2860,2861
_|2861,2862
_|2862,2863
08|2864,2866
:|2866,2867
30AM|2867,2871
BLOOD|2872,2877
ALT|2878,2881
-|2881,2882
20|2882,2884
AST|2885,2888
-|2888,2889
19|2889,2891
AlkPhos|2892,2899
-|2899,2900
77|2900,2902
<EOL>|2902,2903
<EOL>|2903,2904
_|2904,2905
_|2905,2906
_|2906,2907
05|2908,2910
:|2910,2911
58AM|2911,2915
BLOOD|2916,2921
Calcium|2922,2929
-|2929,2930
7|2930,2931
.|2931,2932
6|2932,2933
*|2933,2934
Phos|2935,2939
-|2939,2940
2.8|2940,2943
Mg|2944,2946
-|2946,2947
2.2|2947,2950
<EOL>|2950,2951
_|2951,2952
_|2952,2953
_|2953,2954
06|2955,2957
:|2957,2958
45AM|2958,2962
BLOOD|2963,2968
Calcium|2969,2976
-|2976,2977
7|2977,2978
.|2978,2979
7|2979,2980
*|2980,2981
Phos|2982,2986
-|2986,2987
2|2987,2988
.|2988,2989
4|2989,2990
*|2990,2991
Mg|2992,2994
-|2994,2995
2.1|2995,2998
<EOL>|2998,2999
<EOL>|2999,3000
_|3000,3001
_|3001,3002
_|3002,3003
08|3004,3006
:|3006,3007
30AM|3007,3011
BLOOD|3012,3017
Albumin|3018,3025
-|3025,3026
1|3026,3027
.|3027,3028
8|3028,3029
*|3029,3030
Calcium|3031,3038
-|3038,3039
7|3039,3040
.|3040,3041
7|3041,3042
*|3042,3043
Phos|3044,3048
-|3048,3049
3.5|3049,3052
Mg|3053,3055
-|3055,3056
2.1|3056,3059
<EOL>|3060,3061
Iron|3061,3065
-|3065,3066
23|3066,3068
*|3068,3069
<EOL>|3069,3070
_|3070,3071
_|3071,3072
_|3072,3073
07|3074,3076
:|3076,3077
06PM|3077,3081
BLOOD|3082,3087
Calcium|3088,3095
-|3095,3096
8|3096,3097
.|3097,3098
0|3098,3099
*|3099,3100
Phos|3101,3105
-|3105,3106
5|3106,3107
.|3107,3108
5|3108,3109
*|3109,3110
Mg|3111,3113
-|3113,3114
2.2|3114,3117
<EOL>|3117,3118
_|3118,3119
_|3119,3120
_|3120,3121
08|3122,3124
:|3124,3125
30AM|3125,3129
BLOOD|3130,3135
calTIBC|3136,3143
-|3143,3144
116|3144,3147
*|3147,3148
Ferritn|3149,3156
-|3156,3157
789|3157,3160
*|3160,3161
TRF|3162,3165
-|3165,3166
89|3166,3168
*|3168,3169
<EOL>|3169,3170
_|3170,3171
_|3171,3172
_|3172,3173
05|3174,3176
:|3176,3177
09AM|3177,3181
BLOOD|3182,3187
Triglyc|3188,3195
-|3195,3196
106|3196,3199
<EOL>|3199,3200
_|3200,3201
_|3201,3202
_|3202,3203
08|3204,3206
:|3206,3207
30AM|3207,3211
BLOOD|3212,3217
Triglyc|3218,3225
-|3225,3226
89|3226,3228
<EOL>|3228,3229
<EOL>|3229,3230
_|3230,3231
_|3231,3232
_|3232,3233
07|3234,3236
:|3236,3237
06PM|3237,3241
BLOOD|3242,3247
Lactate|3248,3255
-|3255,3256
1.5|3256,3259
<EOL>|3259,3260
<EOL>|3260,3261
_|3261,3262
_|3262,3263
_|3263,3264
03|3265,3267
:|3267,3268
00PM|3268,3272
ASCITES|3273,3280
Creat|3281,3286
-|3286,3287
0.4|3287,3290
Amylase|3291,3298
-|3298,3299
18|3299,3301
Triglyc|3302,3309
-|3309,3310
29|3310,3312
<EOL>|3313,3314
Lipase|3314,3320
-|3320,3321
8|3321,3322
<EOL>|3322,3323
_|3323,3324
_|3324,3325
_|3325,3326
03|3327,3329
:|3329,3330
00PM|3330,3334
OTHER|3335,3340
BODY|3341,3345
FLUID|3346,3351
Creat|3352,3357
-|3357,3358
0.5|3358,3361
<EOL>|3361,3362
<EOL>|3362,3363
_|3363,3364
_|3364,3365
_|3365,3366
7|3367,3368
:|3368,3369
12|3369,3371
pm|3372,3374
BLOOD|3375,3380
CULTURE|3381,3388
<EOL>|3388,3389
<EOL>|3389,3390
*|3418,3419
*|3419,3420
FINAL|3420,3425
REPORT|3426,3432
_|3433,3434
_|3434,3435
_|3435,3436
<EOL>|3436,3437
<EOL>|3437,3438
Blood|3441,3446
Culture|3447,3454
,|3454,3455
Routine|3456,3463
(|3464,3465
Final|3465,3470
_|3471,3472
_|3472,3473
_|3473,3474
:|3474,3475
<EOL>|3476,3477
CITROBACTER|3483,3494
KOSERI|3495,3501
.|3501,3502
FINAL|3506,3511
SENSITIVITIES|3512,3525
.|3525,3526
<EOL>|3527,3528
<EOL>|3528,3529
SENSITIVITIES|3559,3572
:|3572,3573
MIC|3574,3577
expressed|3578,3587
in|3588,3590
<EOL>|3591,3592
MCG|3592,3595
/|3595,3596
ML|3596,3598
<EOL>|3598,3599
<EOL>|3621,3622
_|3622,3623
_|3623,3624
_|3624,3625
_|3625,3626
_|3626,3627
_|3627,3628
_|3628,3629
_|3629,3630
_|3630,3631
_|3631,3632
_|3632,3633
_|3633,3634
_|3634,3635
_|3635,3636
_|3636,3637
_|3637,3638
_|3638,3639
_|3639,3640
_|3640,3641
_|3641,3642
_|3642,3643
_|3643,3644
_|3644,3645
_|3645,3646
_|3646,3647
_|3647,3648
_|3648,3649
_|3649,3650
_|3650,3651
_|3651,3652
_|3652,3653
_|3653,3654
_|3654,3655
_|3655,3656
_|3656,3657
_|3657,3658
_|3658,3659
_|3659,3660
_|3660,3661
_|3661,3662
_|3662,3663
_|3663,3664
_|3664,3665
_|3665,3666
_|3666,3667
_|3667,3668
_|3668,3669
_|3669,3670
_|3670,3671
_|3671,3672
_|3672,3673
_|3673,3674
_|3674,3675
_|3675,3676
_|3676,3677
_|3677,3678
_|3678,3679
<EOL>|3679,3680
CITROBACTER|3709,3720
KOSERI|3721,3727
<EOL>|3727,3728
||3757,3758
<EOL>|3761,3762
CEFEPIME|3762,3770
-|3770,3771
-|3771,3772
-|3772,3773
-|3773,3774
-|3774,3775
-|3775,3776
-|3776,3777
-|3777,3778
-|3778,3779
-|3779,3780
-|3780,3781
-|3781,3782
-|3782,3783
-|3783,3784
<|3787,3788
=|3788,3789
1|3789,3790
S|3791,3792
<EOL>|3792,3793
CEFTAZIDIME|3793,3804
-|3804,3805
-|3805,3806
-|3806,3807
-|3807,3808
-|3808,3809
-|3809,3810
-|3810,3811
-|3811,3812
-|3812,3813
-|3813,3814
-|3814,3815
<|3818,3819
=|3819,3820
1|3820,3821
S|3822,3823
<EOL>|3823,3824
CEFTRIAXONE|3824,3835
-|3835,3836
-|3836,3837
-|3837,3838
-|3838,3839
-|3839,3840
-|3840,3841
-|3841,3842
-|3842,3843
-|3843,3844
-|3844,3845
-|3845,3846
<|3849,3850
=|3850,3851
1|3851,3852
S|3853,3854
<EOL>|3854,3855
CIPROFLOXACIN|3855,3868
-|3868,3869
-|3869,3870
-|3870,3871
-|3871,3872
-|3872,3873
-|3873,3874
-|3874,3875
-|3875,3876
-|3876,3877
<|3877,3878
=|3878,3879
0.25|3879,3883
S|3884,3885
<EOL>|3885,3886
GENTAMICIN|3886,3896
-|3896,3897
-|3897,3898
-|3898,3899
-|3899,3900
-|3900,3901
-|3901,3902
-|3902,3903
-|3903,3904
-|3904,3905
-|3905,3906
-|3906,3907
-|3907,3908
<|3911,3912
=|3912,3913
1|3913,3914
S|3915,3916
<EOL>|3916,3917
MEROPENEM|3917,3926
-|3926,3927
-|3927,3928
-|3928,3929
-|3929,3930
-|3930,3931
-|3931,3932
-|3932,3933
-|3933,3934
-|3934,3935
-|3935,3936
-|3936,3937
-|3937,3938
-|3938,3939
<|3939,3940
=|3940,3941
0.25|3941,3945
S|3946,3947
<EOL>|3947,3948
PIPERACILLIN|3948,3960
/|3960,3961
TAZO|3961,3965
-|3965,3966
-|3966,3967
-|3967,3968
-|3968,3969
-|3969,3970
<|3973,3974
=|3974,3975
4|3975,3976
S|3977,3978
<EOL>|3978,3979
TOBRAMYCIN|3979,3989
-|3989,3990
-|3990,3991
-|3991,3992
-|3992,3993
-|3993,3994
-|3994,3995
-|3995,3996
-|3996,3997
-|3997,3998
-|3998,3999
-|3999,4000
-|4000,4001
<|4004,4005
=|4005,4006
1|4006,4007
S|4008,4009
<EOL>|4009,4010
TRIMETHOPRIM|4010,4022
/|4022,4023
SULFA|4023,4028
-|4028,4029
-|4029,4030
-|4030,4031
-|4031,4032
<|4035,4036
=|4036,4037
1|4037,4038
S|4039,4040
<EOL>|4040,4041
<EOL>|4041,4042
Aerobic|4045,4052
Bottle|4053,4059
Gram|4060,4064
Stain|4065,4070
(|4071,4072
Final|4072,4077
_|4078,4079
_|4079,4080
_|4080,4081
:|4081,4082
<EOL>|4083,4084
GRAM|4090,4094
NEGATIVE|4095,4103
ROD|4104,4107
(|4107,4108
S|4108,4109
)|4109,4110
.|4110,4111
<EOL>|4112,4113
Reported|4119,4127
to|4128,4130
and|4131,4134
read|4135,4139
back|4140,4144
by|4145,4147
_|4148,4149
_|4149,4150
_|4150,4151
_|4152,4153
_|4153,4154
_|4154,4155
,|4155,4156
@|4157,4158
14|4158,4160
:|4160,4161
35|4161,4163
ON|4164,4166
<EOL>|4167,4168
_|4168,4169
_|4169,4170
_|4170,4171
.|4171,4172
<EOL>|4173,4174
<EOL>|4174,4175
_|4175,4176
_|4176,4177
_|4177,4178
3|4179,4180
:|4180,4181
00|4181,4183
pm|4184,4186
ABSCESS|4187,4194
.|4200,4201
PELVIC|4203,4209
ASPIRATION|4210,4220
.|4220,4221
<EOL>|4222,4223
<EOL>|4223,4224
*|4252,4253
*|4253,4254
FINAL|4254,4259
REPORT|4260,4266
_|4267,4268
_|4268,4269
_|4269,4270
<EOL>|4270,4271
<EOL>|4271,4272
GRAM|4275,4279
STAIN|4280,4285
(|4286,4287
Final|4287,4292
_|4293,4294
_|4294,4295
_|4295,4296
:|4296,4297
<EOL>|4298,4299
4|4305,4306
+|4306,4307
(|4310,4311
>|4311,4312
10|4312,4314
per|4315,4318
1000X|4319,4324
FIELD|4325,4330
)|4330,4331
:|4331,4332
POLYMORPHONUCLEAR|4335,4352
<EOL>|4353,4354
LEUKOCYTES|4354,4364
.|4364,4365
<EOL>|4366,4367
1|4373,4374
+|4374,4375
(|4379,4380
<|4380,4381
1|4381,4382
per|4383,4386
1000X|4387,4392
FIELD|4393,4398
)|4398,4399
:|4399,4400
GRAM|4403,4407
NEGATIVE|4408,4416
ROD|4417,4420
(|4420,4421
S|4421,4422
)|4422,4423
.|4423,4424
<EOL>|4425,4426
<EOL>|4426,4427
WOUND|4430,4435
CULTURE|4436,4443
(|4444,4445
Final|4445,4450
_|4451,4452
_|4452,4453
_|4453,4454
:|4454,4455
NO|4459,4461
GROWTH|4462,4468
.|4468,4469
<EOL>|4470,4471
<EOL>|4471,4472
ANAEROBIC|4475,4484
CULTURE|4485,4492
(|4493,4494
Final|4494,4499
_|4500,4501
_|4501,4502
_|4502,4503
:|4503,4504
<EOL>|4505,4506
BACTEROIDES|4512,4523
FRAGILIS|4524,4532
GROUP|4533,4538
.|4538,4539
SPARSE|4543,4549
GROWTH|4550,4556
.|4556,4557
<EOL>|4558,4559
BETA|4568,4572
LACTAMASE|4573,4582
POSITIVE|4583,4591
.|4591,4592
<EOL>|4593,4594
<EOL>|4594,4595
_|4595,4596
_|4596,4597
_|4597,4598
10|4599,4601
:|4601,4602
52|4602,4604
am|4605,4607
STOOL|4608,4613
CONSISTENCY|4618,4629
:|4629,4630
NOT|4631,4634
APPLICABLE|4635,4645
<EOL>|4645,4646
Source|4652,4658
:|4658,4659
Stool|4660,4665
.|4665,4666
<EOL>|4667,4668
<EOL>|4668,4669
*|4697,4698
*|4698,4699
FINAL|4699,4704
REPORT|4705,4711
_|4712,4713
_|4713,4714
_|4714,4715
<EOL>|4715,4716
<EOL>|4716,4717
C.|4720,4722
difficile|4723,4732
DNA|4733,4736
amplification|4737,4750
assay|4751,4756
(|4757,4758
Final|4758,4763
_|4764,4765
_|4765,4766
_|4766,4767
:|4767,4768
<EOL>|4769,4770
Negative|4776,4784
for|4785,4788
toxigenic|4789,4798
C.|4799,4801
difficile|4802,4811
by|4812,4814
the|4815,4818
Illumigene|4819,4829
DNA|4830,4833
<EOL>|4833,4834
amplification|4840,4853
assay|4854,4859
.|4859,4860
<EOL>|4861,4862
(|4873,4874
Reference|4874,4883
Range|4884,4889
-|4889,4890
Negative|4890,4898
)|4898,4899
.|4899,4900
<EOL>|4901,4902
<EOL>|4902,4903
<EOL>|4904,4905
Ms.|4928,4931
_|4932,4933
_|4933,4934
_|4934,4935
was|4936,4939
admitted|4940,4948
to|4949,4951
Dr.|4952,4955
_|4956,4957
_|4957,4958
_|4958,4959
service|4960,4967
for|4968,4971
<EOL>|4972,4973
management|4973,4983
of|4984,4986
ileus|4987,4992
.|4992,4993
Upon|4995,4999
admission|5000,5009
,|5009,5010
a|5011,5012
nasogastric|5013,5024
tube|5025,5029
was|5030,5033
<EOL>|5034,5035
placed|5035,5041
for|5042,5045
decompression|5046,5059
.|5059,5060
On|5062,5064
_|5065,5066
_|5066,5067
_|5067,5068
,|5068,5069
PICC|5070,5074
was|5075,5078
placed|5079,5085
and|5086,5089
TPN|5090,5093
<EOL>|5094,5095
started|5095,5102
.|5102,5103
Blood|5105,5110
cultures|5111,5119
grew|5120,5124
gram|5125,5129
negative|5130,5138
rods|5139,5143
and|5144,5147
ceftriaxone|5148,5159
<EOL>|5160,5161
was|5161,5164
started|5165,5172
.|5172,5173
On|5175,5177
_|5178,5179
_|5179,5180
_|5180,5181
,|5181,5182
pt|5183,5185
started|5186,5193
to|5194,5196
pass|5197,5201
small|5202,5207
amount|5208,5214
of|5215,5217
<EOL>|5218,5219
flatus|5219,5225
.|5225,5226
_|5228,5229
_|5229,5230
_|5230,5231
CT|5232,5234
scan|5235,5239
demonstrated|5240,5252
improving|5253,5262
ileus|5263,5268
,|5268,5269
but|5270,5273
concern|5274,5281
<EOL>|5282,5283
for|5283,5286
possible|5287,5295
urine|5296,5301
leak|5302,5306
and|5307,5310
increased|5311,5320
free|5321,5325
fluid|5326,5331
.|5331,5332
On|5334,5336
_|5337,5338
_|5338,5339
_|5339,5340
,|5340,5341
a|5342,5343
<EOL>|5344,5345
LLQ|5345,5348
drain|5349,5354
was|5355,5358
placed|5359,5365
by|5366,5368
interventional|5369,5383
radiology|5384,5393
.|5393,5394
on|5396,5398
_|5399,5400
_|5400,5401
_|5401,5402
,|5402,5403
pt|5404,5406
<EOL>|5407,5408
passed|5408,5414
clamp|5415,5420
trial|5421,5426
and|5427,5430
NGT|5431,5434
was|5435,5438
removed|5439,5446
.|5446,5447
Pt|5449,5451
continued|5452,5461
to|5462,5464
pass|5465,5469
<EOL>|5470,5471
flatus|5471,5477
and|5478,5481
also|5482,5486
started|5487,5494
to|5495,5497
have|5498,5502
bowel|5503,5508
movements|5509,5518
.|5518,5519
On|5521,5523
_|5524,5525
_|5525,5526
_|5526,5527
,|5527,5528
pt|5529,5531
<EOL>|5532,5533
was|5533,5536
advanced|5537,5545
to|5546,5548
a|5549,5550
clear|5551,5556
liquid|5557,5563
diet|5564,5568
.|5568,5569
Repeat|5571,5577
blood|5578,5583
cultures|5584,5592
were|5593,5597
<EOL>|5598,5599
negative|5599,5607
and|5608,5611
positive|5612,5620
blood|5621,5626
culture|5627,5634
from|5635,5639
admission|5640,5649
grew|5650,5654
<EOL>|5655,5656
citrobacter|5656,5667
.|5667,5668
Diet|5670,5674
was|5675,5678
gradually|5679,5688
advanced|5689,5697
and|5698,5701
ensure|5702,5708
added|5709,5714
.|5714,5715
IV|5716,5718
<EOL>|5719,5720
medications|5720,5731
were|5732,5736
gradually|5737,5746
converted|5747,5756
to|5757,5759
PO|5760,5762
and|5763,5766
she|5767,5770
was|5771,5774
<EOL>|5775,5776
re-evaluated|5776,5788
by|5789,5791
physical|5792,5800
therapy|5801,5808
for|5809,5812
rehabilitative|5813,5827
services|5828,5836
.|5836,5837
<EOL>|5838,5839
She|5839,5842
was|5843,5846
ambulating|5847,5857
with|5858,5862
walker|5863,5869
assistance|5870,5880
and|5881,5884
prepared|5885,5893
for|5894,5897
<EOL>|5898,5899
discharge|5899,5908
to|5909,5911
her|5912,5915
_|5916,5917
_|5917,5918
_|5918,5919
facility|5920,5928
(|5929,5930
_|5930,5931
_|5931,5932
_|5932,5933
)|5933,5934
.|5934,5935
TPN|5936,5939
was|5940,5943
<EOL>|5944,5945
continued|5945,5954
up|5955,5957
until|5958,5963
day|5964,5967
before|5968,5974
discharge|5975,5984
.|5984,5985
At|5986,5988
time|5989,5993
of|5994,5996
discharge|5997,6006
,|6006,6007
<EOL>|6008,6009
she|6009,6012
was|6013,6016
tolerating|6017,6027
regular|6028,6035
diet|6036,6040
,|6040,6041
passing|6042,6049
flatus|6050,6056
regularly|6057,6066
and|6067,6070
<EOL>|6071,6072
having|6072,6078
bowel|6079,6084
movements|6085,6094
.|6094,6095
<EOL>|6096,6097
<EOL>|6098,6099
Medications|6099,6110
on|6111,6113
Admission|6114,6123
:|6123,6124
<EOL>|6124,6125
The|6125,6128
Preadmission|6129,6141
Medication|6142,6152
list|6153,6157
is|6158,6160
accurate|6161,6169
and|6170,6173
complete|6174,6182
.|6182,6183
<EOL>|6183,6184
1.|6184,6186
Atorvastatin|6187,6199
10|6200,6202
mg|6203,6205
PO|6206,6208
QPM|6209,6212
<EOL>|6213,6214
2.|6214,6216
Levothyroxine|6217,6230
Sodium|6231,6237
175|6238,6241
mcg|6242,6245
PO|6246,6248
DAILY|6249,6254
<EOL>|6255,6256
3.|6256,6258
Losartan|6259,6267
Potassium|6268,6277
50|6278,6280
mg|6281,6283
PO|6284,6286
DAILY|6287,6292
<EOL>|6293,6294
4.|6294,6296
Acetaminophen|6297,6310
650|6311,6314
mg|6315,6317
PO|6318,6320
Q6H|6321,6324
<EOL>|6325,6326
5.|6326,6328
Docusate|6329,6337
Sodium|6338,6344
100|6345,6348
mg|6349,6351
PO|6352,6354
BID|6355,6358
<EOL>|6359,6360
6.|6360,6362
Enoxaparin|6363,6373
Sodium|6374,6380
40|6381,6383
mg|6384,6386
SC|6387,6389
DAILY|6390,6395
<EOL>|6396,6397
7.|6397,6399
Nitrofurantoin|6400,6414
Monohyd|6415,6422
(|6423,6424
MacroBID|6424,6432
)|6432,6433
100|6434,6437
mg|6438,6440
PO|6441,6443
DAILY|6444,6449
<EOL>|6450,6451
8.|6451,6453
OxyCODONE|6454,6463
(|6464,6465
Immediate|6465,6474
Release|6475,6482
)|6482,6483
5|6484,6485
mg|6486,6488
PO|6489,6491
Q4H|6492,6495
:|6495,6496
PRN|6496,6499
Pain|6500,6504
-|6505,6506
Moderate|6507,6515
<EOL>|6516,6517
<EOL>|6517,6518
<EOL>|6518,6519
<EOL>|6520,6521
Discharge|6521,6530
Medications|6531,6542
:|6542,6543
<EOL>|6543,6544
1.|6544,6546
Ciprofloxacin|6548,6561
HCl|6562,6565
500|6566,6569
mg|6570,6572
PO|6573,6575
Q12H|6576,6580
Duration|6581,6589
:|6589,6590
7|6591,6592
Days|6593,6597
<EOL>|6598,6599
Last|6599,6603
dose|6604,6608
_|6609,6610
_|6610,6611
_|6611,6612
<EOL>|6614,6615
2.|6615,6617
MetroNIDAZOLE|6619,6632
500|6633,6636
mg|6637,6639
PO|6640,6642
Q6H|6643,6646
Duration|6647,6655
:|6655,6656
7|6657,6658
Days|6659,6663
<EOL>|6664,6665
Last|6665,6669
dose|6670,6674
_|6675,6676
_|6676,6677
_|6677,6678
<EOL>|6680,6681
3.|6681,6683
Senna|6685,6690
8.6|6691,6694
mg|6695,6697
PO|6698,6700
BID|6701,6704
<EOL>|6706,6707
4.|6707,6709
Acetaminophen|6711,6724
650|6725,6728
mg|6729,6731
PO|6732,6734
Q6H|6735,6738
<EOL>|6740,6741
5.|6741,6743
Atorvastatin|6745,6757
10|6758,6760
mg|6761,6763
PO|6764,6766
QPM|6767,6770
<EOL>|6772,6773
6.|6773,6775
Docusate|6777,6785
Sodium|6786,6792
100|6793,6796
mg|6797,6799
PO|6800,6802
BID|6803,6806
<EOL>|6808,6809
7.|6809,6811
Enoxaparin|6813,6823
Sodium|6824,6830
40|6831,6833
mg|6834,6836
SC|6837,6839
DAILY|6840,6845
<EOL>|6846,6847
Start|6847,6852
:|6852,6853
_|6854,6855
_|6855,6856
_|6856,6857
,|6857,6858
First|6859,6864
Dose|6865,6869
:|6869,6870
Next|6871,6875
Routine|6876,6883
Administration|6884,6898
Time|6899,6903
<EOL>|6905,6906
8.|6906,6908
Levothyroxine|6910,6923
Sodium|6924,6930
175|6931,6934
mcg|6935,6938
PO|6939,6941
DAILY|6942,6947
<EOL>|6949,6950
9.|6950,6952
LORazepam|6954,6963
0.25|6964,6968
mg|6969,6971
PO|6972,6974
BID|6975,6978
:|6978,6979
PRN|6979,6982
anxiety|6983,6990
<EOL>|6992,6993
10.|6993,6996
Losartan|6998,7006
Potassium|7007,7016
50|7017,7019
mg|7020,7022
PO|7023,7025
DAILY|7026,7031
<EOL>|7033,7034
11.|7034,7037
Nitrofurantoin|7039,7053
Monohyd|7054,7061
(|7062,7063
MacroBID|7063,7071
)|7071,7072
100|7073,7076
mg|7077,7079
PO|7080,7082
DAILY|7083,7088
<EOL>|7090,7091
12.|7091,7094
OxyCODONE|7096,7105
(|7106,7107
Immediate|7107,7116
Release|7117,7124
)|7124,7125
5|7126,7127
mg|7128,7130
PO|7131,7133
Q4H|7134,7137
:|7137,7138
PRN|7138,7141
Pain|7142,7146
-|7147,7148
<EOL>|7149,7150
Moderate|7150,7158
<EOL>|7160,7161
<EOL>|7161,7162
<EOL>|7163,7164
Discharge|7164,7173
Disposition|7174,7185
:|7185,7186
<EOL>|7186,7187
Extended|7187,7195
Care|7196,7200
<EOL>|7200,7201
<EOL>|7202,7203
Facility|7203,7211
:|7211,7212
<EOL>|7212,7213
_|7213,7214
_|7214,7215
_|7215,7216
<EOL>|7216,7217
<EOL>|7218,7219
Discharge|7219,7228
Diagnosis|7229,7238
:|7238,7239
<EOL>|7239,7240
bladder|7240,7247
cancer|7248,7254
,|7254,7255
post-operative|7256,7270
ileus|7271,7276
,|7276,7277
bacteremia|7278,7288
(|7289,7290
CITROBACTER|7290,7301
<EOL>|7302,7303
KOSERI|7303,7309
)|7309,7310
and|7311,7314
abdominal|7315,7324
-|7324,7325
pelvic|7325,7331
abscess|7332,7339
(|7340,7341
BACTEROIDES|7341,7352
FRAGILIS|7353,7361
<EOL>|7362,7363
GROUP|7363,7368
)|7368,7369
requiring|7370,7379
_|7380,7381
_|7381,7382
_|7382,7383
drainage|7384,7392
<EOL>|7392,7393
<EOL>|7393,7394
<EOL>|7395,7396
Mental|7417,7423
Status|7424,7430
:|7430,7431
Clear|7432,7437
and|7438,7441
coherent|7442,7450
.|7450,7451
<EOL>|7451,7452
Level|7452,7457
of|7458,7460
Consciousness|7461,7474
:|7474,7475
Alert|7476,7481
and|7482,7485
interactive|7486,7497
.|7497,7498
<EOL>|7498,7499
Activity|7499,7507
Status|7508,7514
:|7514,7515
Ambulatory|7516,7526
-|7527,7528
requires|7529,7537
assistance|7538,7548
or|7549,7551
aid|7552,7555
(|7556,7557
walker|7557,7563
<EOL>|7564,7565
or|7565,7567
cane|7568,7572
)|7572,7573
.|7573,7574
<EOL>|7574,7575
<EOL>|7575,7576
<EOL>|7577,7578
-|7602,7603
Please|7603,7609
also|7610,7614
refer|7615,7620
to|7621,7623
the|7624,7627
instructions|7628,7640
provided|7641,7649
to|7650,7652
you|7653,7656
by|7657,7659
the|7660,7663
<EOL>|7664,7665
Ostomy|7665,7671
nurse|7672,7677
specialist|7678,7688
that|7689,7693
details|7694,7701
the|7702,7705
required|7706,7714
care|7715,7719
and|7720,7723
<EOL>|7724,7725
management|7725,7735
of|7736,7738
your|7739,7743
Urostomy|7744,7752
<EOL>|7752,7753
<EOL>|7753,7754
-|7754,7755
Resume|7755,7761
your|7762,7766
pre-admission|7767,7780
/|7780,7781
home|7781,7785
medications|7786,7797
except|7798,7804
as|7805,7807
noted|7808,7813
.|7813,7814
<EOL>|7815,7816
Always|7816,7822
call|7823,7827
to|7828,7830
inform|7831,7837
,|7837,7838
review|7839,7845
and|7846,7849
discuss|7850,7857
any|7858,7861
medication|7862,7872
changes|7873,7880
<EOL>|7881,7882
and|7882,7885
your|7886,7890
post-operative|7891,7905
course|7906,7912
with|7913,7917
your|7918,7922
primary|7923,7930
care|7931,7935
doctor|7936,7942
<EOL>|7942,7943
<EOL>|7943,7944
-|7944,7945
_|7945,7946
_|7946,7947
_|7947,7948
(|7949,7950
acetaminophen|7950,7963
)|7963,7964
and|7965,7968
Ibuprofen|7969,7978
for|7979,7982
pain|7983,7987
control|7988,7995
.|7995,7996
<EOL>|7996,7997
<EOL>|7997,7998
-|7998,7999
Ciprofloxacin|7999,8012
and|8013,8016
Metronidazole|8017,8030
are|8031,8034
new|8035,8038
ANTIBIOTIC|8039,8049
medications|8050,8061
<EOL>|8062,8063
to|8063,8065
treat|8066,8071
your|8072,8076
infection|8077,8086
.|8086,8087
Continue|8088,8096
for|8097,8100
7|8101,8102
days|8103,8107
through|8108,8115
_|8116,8117
_|8117,8118
_|8118,8119
.|8119,8120
<EOL>|8120,8121
<EOL>|8121,8122
-|8122,8123
The|8123,8126
MAXIMUM|8127,8134
dose|8135,8139
of|8140,8142
Tylenol|8143,8150
(|8151,8152
ACETAMINOPHEN|8152,8165
)|8165,8166
is|8167,8169
3|8170,8171
grams|8172,8177
(|8178,8179
from|8179,8183
<EOL>|8184,8185
ALL|8185,8188
sources|8189,8196
)|8196,8197
PER|8198,8201
DAY|8202,8205
<EOL>|8206,8207
<EOL>|8207,8208
-|8208,8209
If|8209,8211
you|8212,8215
are|8216,8219
taking|8220,8226
Ibuprofen|8227,8236
(|8237,8238
Brand|8238,8243
names|8244,8249
include|8250,8257
_|8258,8259
_|8259,8260
_|8260,8261
<EOL>|8262,8263
this|8263,8267
should|8268,8274
always|8275,8281
be|8282,8284
taken|8285,8290
with|8291,8295
food|8296,8300
.|8300,8301
If|8302,8304
you|8305,8308
develop|8309,8316
stomach|8317,8324
<EOL>|8325,8326
pain|8326,8330
or|8331,8333
note|8334,8338
black|8339,8344
stool|8345,8350
,|8350,8351
stop|8352,8356
the|8357,8360
Ibuprofen|8361,8370
.|8370,8371
<EOL>|8371,8372
<EOL>|8372,8373
-|8373,8374
Please|8374,8380
do|8381,8383
NOT|8384,8387
drive|8388,8393
,|8393,8394
operate|8395,8402
dangerous|8403,8412
machinery|8413,8422
,|8422,8423
or|8424,8426
consume|8427,8434
<EOL>|8435,8436
alcohol|8436,8443
while|8444,8449
taking|8450,8456
narcotic|8457,8465
pain|8466,8470
medications|8471,8482
.|8482,8483
<EOL>|8483,8484
<EOL>|8484,8485
-|8485,8486
Do|8486,8488
NOT|8489,8492
drive|8493,8498
and|8499,8502
until|8503,8508
you|8509,8512
are|8513,8516
cleared|8517,8524
to|8525,8527
resume|8528,8534
such|8535,8539
<EOL>|8540,8541
activities|8541,8551
by|8552,8554
your|8555,8559
PCP|8560,8563
or|8564,8566
urologist|8567,8576
.|8576,8577
You|8578,8581
may|8582,8585
be|8586,8588
a|8589,8590
passenger|8591,8600
<EOL>|8600,8601
<EOL>|8601,8602
-|8602,8603
Colace|8603,8609
may|8610,8613
have|8614,8618
been|8619,8623
prescribed|8624,8634
to|8635,8637
avoid|8638,8643
post|8644,8648
surgical|8649,8657
<EOL>|8658,8659
constipation|8659,8671
and|8672,8675
constipation|8676,8688
related|8689,8696
to|8697,8699
narcotic|8700,8708
pain|8709,8713
<EOL>|8714,8715
medication|8715,8725
.|8725,8726
Discontinue|8727,8738
if|8739,8741
loose|8742,8747
stool|8748,8753
or|8754,8756
diarrhea|8757,8765
develops|8766,8774
.|8774,8775
<EOL>|8776,8777
Colace|8777,8783
is|8784,8786
a|8787,8788
stool|8789,8794
-|8794,8795
softener|8795,8803
,|8803,8804
NOT|8805,8808
a|8809,8810
laxative|8811,8819
.|8819,8820
<EOL>|8820,8821
<EOL>|8821,8822
-|8822,8823
No|8823,8825
heavy|8826,8831
lifting|8832,8839
for|8840,8843
4|8844,8845
weeks|8846,8851
(|8852,8853
no|8853,8855
more|8856,8860
than|8861,8865
10|8866,8868
pounds|8869,8875
)|8875,8876
.|8876,8877
Do|8878,8880
"|8881,8882
not|8882,8885
"|8885,8886
<EOL>|8887,8888
be|8888,8890
sedentary|8891,8900
.|8900,8901
Walk|8902,8906
frequently|8907,8917
.|8917,8918
Light|8919,8924
household|8925,8934
chores|8935,8941
(|8942,8943
cooking|8943,8950
,|8950,8951
<EOL>|8952,8953
folding|8953,8960
laundry|8961,8968
,|8968,8969
washing|8970,8977
dishes|8978,8984
)|8984,8985
are|8986,8989
generally|8990,8999
|9000,9001
ok|9001,9003
|9003,9004
but|9005,9008
AGAIN|9009,9014
,|9014,9015
<EOL>|9016,9017
avoid|9017,9022
straining|9023,9032
,|9032,9033
pulling|9034,9041
,|9041,9042
twisting|9043,9051
(|9052,9053
do|9053,9055
NOT|9056,9059
vacuum|9060,9066
)|9066,9067
.|9067,9068
<EOL>|9068,9069
<EOL>|9069,9070
<EOL>|9071,9072
Followup|9072,9080
Instructions|9081,9093
:|9093,9094
<EOL>|9094,9095
_|9095,9096
_|9096,9097
_|9097,9098
<EOL>|9098,9099

