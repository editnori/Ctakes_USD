 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|44,53|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|44,58|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|78,87|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|78,87|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|78,92|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|110,115|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|134,137|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|134,137|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|145,152|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|145,152|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|154,162|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|186,195|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|186,195|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|198,220|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|206,210|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|206,210|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|206,220|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|223,232|false|false|false|C1999232|Attending (action)|Attending
Finding|Pathologic Function|Chief Complaint|257,266|false|false|false|C0014591|Epistaxis|Epistaxis
Finding|Classification|Chief Complaint|269,274|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|275,283|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|287,305|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|296,305|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|296,305|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|296,305|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|296,305|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|366,373|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|366,376|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|History of Present Illness|377,380|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|History of Present Illness|377,380|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|History of Present Illness|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|History of Present Illness|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|History of Present Illness|377,380|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Finding|Gene or Genome|History of Present Illness|377,380|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Finding|Functional Concept|History of Present Illness|385,391|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|History of Present Illness|385,391|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|History of Present Illness|385,391|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|385,391|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|History of Present Illness|412,424|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|History of Present Illness|430,444|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|History of Present Illness|430,444|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Finding|Functional Concept|History of Present Illness|464,472|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|464,472|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|464,472|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Idea or Concept|History of Present Illness|486,494|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|500,505|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|500,505|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|500,505|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|500,505|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|History of Present Illness|506,515|false|false|false|C0016658|Fracture|fractures
Finding|Finding|History of Present Illness|506,515|false|false|false|C4554413|Fractured|fractures
Finding|Pathologic Function|History of Present Illness|521,530|false|false|false|C0014591|Epistaxis|epistaxis
Disorder|Neoplastic Process|History of Present Illness|531,540|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|History of Present Illness|531,540|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Finding|History of Present Illness|544,548|false|false|false|C0085639|Falls|fall
Finding|Body Substance|History of Present Illness|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|554,561|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|History of Present Illness|653,657|false|false|false|C0263940|Curb|curb
Disorder|Injury or Poisoning|History of Present Illness|671,677|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|History of Present Illness|671,677|false|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Location or Region|History of Present Illness|685,689|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|History of Present Illness|685,689|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|History of Present Illness|685,689|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Finding|Finding|History of Present Illness|701,705|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|History of Present Illness|710,723|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|History of Present Illness|710,723|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Disorder|Injury or Poisoning|History of Present Illness|791,797|false|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|History of Present Illness|791,797|false|false|false|C0548346|Trauma assessment and care|trauma
Anatomy|Body Location or Region|History of Present Illness|805,809|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|History of Present Illness|805,809|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|History of Present Illness|805,809|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Activity|History of Present Illness|852,856|false|false|false|C1947933|care activity|care
Finding|Finding|History of Present Illness|852,856|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|852,856|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Procedure|Diagnostic Procedure|History of Present Illness|867,874|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|History of Present Illness|870,874|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Anatomy|Body Location or Region|History of Present Illness|883,887|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|883,887|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|883,887|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|883,887|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|History of Present Illness|889,893|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|889,893|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|889,893|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Location or Region|History of Present Illness|899,903|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|History of Present Illness|899,903|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Finding|Gene or Genome|History of Present Illness|899,903|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|926,931|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|926,931|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|926,931|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|926,931|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|926,936|false|false|false|C0027422|Nasal bone structure|nasal bone
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|932,936|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|History of Present Illness|932,936|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|History of Present Illness|932,936|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Injury or Poisoning|History of Present Illness|949,957|false|false|false|C0016658|Fracture|fracture
Finding|Pathologic Function|History of Present Illness|976,985|false|false|false|C0014591|Epistaxis|epistaxis
Disorder|Injury or Poisoning|History of Present Illness|1039,1047|false|false|false|C0043242;C0518443;C1302752|Abrasion;Superficial abrasion;skin abrasion|abrasion
Drug|Pharmacologic Substance|History of Present Illness|1039,1047|false|false|false|C1627366|Abrasion Pharmacologic Substance|abrasion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1039,1047|false|false|false|C0580209|Surgical abrasion|abrasion
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1055,1061|false|false|false|C0399080|Fixation of dental bridge|bridge
Finding|Pathologic Function|History of Present Illness|1097,1105|false|false|false|C0019080|Hemorrhage|Bleeding
Finding|Finding|History of Present Illness|1110,1114|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|History of Present Illness|1170,1176|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|1170,1176|false|false|false|C0027497|Nausea|nausea
Disorder|Disease or Syndrome|History of Present Illness|1198,1203|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|History of Present Illness|1198,1203|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|History of Present Illness|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1213,1217|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Sign or Symptom|History of Present Illness|1236,1247|false|false|false|C0220870|Lightheadedness|lightheaded
Finding|Pathologic Function|History of Present Illness|1269,1280|false|false|false|C0857353|Hypotensive|hypotensive
Attribute|Clinical Attribute|History of Present Illness|1302,1308|false|false|false|C4255046||report
Finding|Intellectual Product|History of Present Illness|1302,1308|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|History of Present Illness|1302,1308|false|false|false|C0700287|Reporting|report
Finding|Intellectual Product|History of Present Illness|1320,1325|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1320,1347|false|false|false|C0234431|Brief loss of consciousness|brief loss of consciousness
Finding|Finding|History of Present Illness|1326,1330|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Finding|History of Present Illness|1326,1347|false|false|false|C0041657|Unconscious State|loss of consciousness
Finding|Finding|History of Present Illness|1334,1347|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Finding|Mental Process|History of Present Illness|1334,1347|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|consciousness
Drug|Biomedical or Dental Material|History of Present Illness|1381,1389|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|History of Present Illness|1381,1389|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Classification|History of Present Illness|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|1395,1401|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1417,1421|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|History of Present Illness|1417,1421|false|false|false|C5848506||eyes
Anatomy|Body Location or Region|History of Present Illness|1444,1448|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1444,1448|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1444,1448|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1444,1448|false|false|false|C0876917|Procedure on head|head
Finding|Body Substance|History of Present Illness|1454,1461|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1454,1461|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1454,1461|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1474,1479|false|false|false|C0441471|Event|event
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1503,1512|false|false|false|C0009676|Confusion|confusion
Finding|Finding|History of Present Illness|1503,1512|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Sign or Symptom|History of Present Illness|1544,1551|true|false|false|C0039070|Syncope|syncope
Finding|Organ or Tissue Function|History of Present Illness|1555,1566|false|false|false|C0019010|Hemodynamics|hemodynamic
Procedure|Laboratory Procedure|History of Present Illness|1555,1566|false|false|false|C4281788|hemodynamics (procedure)|hemodynamic
Finding|Functional Concept|History of Present Illness|1568,1575|false|false|false|C0392747|Changing|changes
Event|Event|History of Present Illness|1597,1602|false|false|false|C0441471|Event|event
Finding|Pathologic Function|History of Present Illness|1607,1616|false|false|false|C0014591|Epistaxis|epistaxis
Finding|Body Substance|History of Present Illness|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1622,1629|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Activity|History of Present Illness|1659,1663|false|false|false|C1947933|care activity|care
Finding|Finding|History of Present Illness|1659,1663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|History of Present Illness|1659,1663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|History of Present Illness|1677,1684|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|1685,1690|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|1685,1696|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|1685,1696|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|History of Present Illness|1691,1696|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|1691,1696|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Lab|Laboratory or Test Result|History of Present Illness|1724,1728|false|false|false|C0587081|Laboratory test finding|Labs
Anatomy|Cell|History of Present Illness|1747,1750|false|false|false|C0023516|Leukocytes|WBC
Procedure|Laboratory Procedure|History of Present Illness|1779,1782|false|false|false|C0201617|Primed lymphocyte test|plt
Drug|Biologically Active Substance|History of Present Illness|1788,1791|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|1788,1791|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|History of Present Illness|1788,1791|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Finding|Intellectual Product|History of Present Illness|1834,1840|false|false|false|C1547311|Patient Condition Code - Stable|stable
Procedure|Laboratory Procedure|History of Present Illness|1844,1854|false|false|false|C0042014;C0373521|Urinalysis;Urinalysis; qualitative or semiquantitative, except immunoassays|urinalysis
Finding|Classification|History of Present Illness|1860,1868|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1860,1868|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1860,1868|false|false|false|C5237010|Expression Negative|negative
Procedure|Diagnostic Procedure|History of Present Illness|1872,1875|false|false|false|C0039985|Plain chest X-ray|CXR
Disorder|Disease or Syndrome|History of Present Illness|1897,1910|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|History of Present Illness|1918,1922|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|1924,1928|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1924,1928|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|History of Present Illness|1924,1928|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|History of Present Illness|1924,1928|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1924,1933|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|History of Present Illness|1929,1933|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|History of Present Illness|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|History of Present Illness|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|1929,1933|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|History of Present Illness|1929,1933|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|History of Present Illness|1929,1933|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Finding|History of Present Illness|1935,1943|false|false|false|C0332149|Possible|possibly
Disorder|Injury or Poisoning|History of Present Illness|1957,1967|false|false|false|C1720922|Respiratory Aspiration|aspiration
Finding|Finding|History of Present Illness|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|History of Present Illness|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|History of Present Illness|1957,1967|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1957,1967|false|false|false|C0349707||aspiration
Disorder|Disease or Syndrome|History of Present Illness|1983,1992|false|false|false|C0032285|Pneumonia|pneumonia
Finding|Body Substance|History of Present Illness|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1998,2005|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Immunologic Factor|History of Present Illness|2016,2020|false|false|false|C3526553;C3644171|diphtheria, tetanus toxoids and acellular pertussis vaccine;tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Tdap
Drug|Pharmacologic Substance|History of Present Illness|2016,2020|false|false|false|C3526553;C3644171|diphtheria, tetanus toxoids and acellular pertussis vaccine;tetanus toxoid, reduced diphtheria toxoid, and acellular pertussis vaccine, adsorbed|Tdap
Drug|Antibiotic|History of Present Illness|2022,2033|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Organic Chemical|History of Present Illness|2022,2033|false|false|false|C0002645|amoxicillin|amoxicillin
Drug|Pharmacologic Substance|History of Present Illness|2022,2045|false|false|false|C0054066|amoxicillin / clavulanate|amoxicillin-clavulanate
Drug|Antibiotic|History of Present Illness|2034,2045|false|false|false|C0110038|clavulanate|clavulanate
Drug|Organic Chemical|History of Present Illness|2034,2045|false|false|false|C0110038|clavulanate|clavulanate
Drug|Antibiotic|History of Present Illness|2051,2061|false|false|false|C0003232|Antibiotics|antibiotic
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2051,2073|false|false|false|C0282638|Antibiotic Prophylaxis|antibiotic prophylaxis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|2062,2073|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Drug|Organic Chemical|History of Present Illness|2075,2086|false|false|false|C0061851|ondansetron|ondansetron
Drug|Pharmacologic Substance|History of Present Illness|2075,2086|false|false|false|C0061851|ondansetron|ondansetron
Drug|Organic Chemical|History of Present Illness|2103,2113|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|History of Present Illness|2103,2113|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|History of Present Illness|2103,2122|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|History of Present Illness|2103,2122|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|History of Present Illness|2114,2122|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|History of Present Illness|2114,2122|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Organic Chemical|History of Present Illness|2129,2140|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|History of Present Illness|2129,2140|false|false|false|C0070166|clopidogrel|Clopidogrel
Disorder|Anatomical Abnormality|Past Medical History|2184,2187|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Past Medical History|2184,2187|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Past Medical History|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Past Medical History|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Past Medical History|2184,2187|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Finding|Gene or Genome|Past Medical History|2184,2187|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Finding|Functional Concept|Past Medical History|2188,2194|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Past Medical History|2188,2194|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Past Medical History|2188,2194|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2188,2194|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|Past Medical History|2215,2218|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Past Medical History|2219,2239|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Finding|Finding|Past Medical History|2219,2239|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Finding|Body Substance|Family Medical History|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Family Medical History|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Family Medical History|2278,2285|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Research Activity|Family Medical History|2289,2296|false|false|false|C0150114|unaware|unaware
Finding|Classification|Family Medical History|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2302,2308|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Finding|Family Medical History|2302,2316|false|false|false|C0241889|Family Medical History|family history
Finding|Finding|Family Medical History|2302,2319|false|false|false|C0241889|Family Medical History|family history of
Finding|Conceptual Entity|Family Medical History|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|2309,2316|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|2309,2319|false|false|false|C0262926|Medical History|history of
Finding|Pathologic Function|Family Medical History|2320,2328|false|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|Family Medical History|2320,2338|false|false|false|C0005779|Blood Coagulation Disorders|bleeding diathesis
Finding|Pathologic Function|Family Medical History|2320,2338|false|false|false|C1458140|Bleeding tendency|bleeding diathesis
Attribute|Clinical Attribute|Family Medical History|2329,2338|false|false|false|C0012655|Disease susceptibility|diathesis
Procedure|Health Care Activity|General Exam|2358,2367|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Classification|General Exam|2396,2403|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2396,2403|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|General Exam|2405,2410|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|2405,2410|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|2405,2410|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|2405,2410|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|2405,2410|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2405,2410|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2425,2430|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|2431,2439|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2431,2439|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2442,2447|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2457,2466|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2468,2471|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|2468,2471|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|2473,2483|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|2484,2489|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Injury or Poisoning|General Exam|2491,2499|false|false|false|C0009938|Contusions|bruising
Finding|Finding|General Exam|2491,2499|false|false|false|C2136686|reported bruising (history)|bruising
Anatomy|Body Part, Organ, or Organ Component|General Exam|2507,2516|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|General Exam|2512,2516|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|2512,2516|false|false|false|C5848506||eyes
Finding|Finding|General Exam|2518,2525|false|false|false|C0038999|Swelling|swollen
Finding|Finding|General Exam|2518,2530|false|false|false|C0240577|Swollen nose|swollen nose
Finding|Intellectual Product|General Exam|2536,2540|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Mental Process|General Exam|2541,2551|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|2541,2551|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Activity|General Exam|2570,2575|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|2570,2575|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|2570,2575|false|false|false|C1533810||place
Anatomy|Body Location or Region|General Exam|2578,2582|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|2578,2582|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|2578,2582|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|2584,2590|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|2600,2603|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|2600,2603|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|General Exam|2600,2603|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|General Exam|2606,2610|false|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|General Exam|2606,2610|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Drug|Amino Acid, Peptide, or Protein|General Exam|2622,2625|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|General Exam|2622,2625|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|2622,2625|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|2669,2672|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|2669,2672|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|2674,2678|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Disorder|Congenital Abnormality|General Exam|2720,2723|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Finding|Gene or Genome|General Exam|2720,2723|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Finding|General Exam|2725,2729|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2725,2729|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2731,2735|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|2749,2755|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|2749,2755|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|2749,2755|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|2760,2768|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|General Exam|2770,2778|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|2783,2788|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|2783,2788|false|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|2816,2822|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|General Exam|2824,2829|false|false|false|C1513492|motor movement|motor
Finding|Finding|General Exam|2824,2838|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|General Exam|2824,2838|false|false|false|C0234130|Motor function (observable entity)|motor function
Finding|Finding|General Exam|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|2830,2838|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Anatomy|Body System|General Exam|2854,2858|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|2854,2858|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|2854,2858|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|2854,2858|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|2854,2858|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Injury or Poisoning|General Exam|2863,2875|true|false|false|C0015256|Excoriation|excoriations
Disorder|Disease or Syndrome|General Exam|2879,2883|true|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|General Exam|2879,2883|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|2879,2883|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Body Substance|General Exam|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2886,2895|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2886,2895|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Classification|General Exam|2924,2931|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2924,2931|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|General Exam|2933,2938|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|2933,2938|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|2933,2938|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|2933,2938|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|2933,2938|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2933,2938|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2953,2958|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|2959,2967|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2959,2967|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2970,2975|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2985,2994|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2996,2999|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|2996,2999|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3001,3011|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|3012,3017|false|false|false|C1550016|Remote control command - Clear|clear
Disorder|Injury or Poisoning|General Exam|3019,3027|false|false|false|C0009938|Contusions|bruising
Finding|Finding|General Exam|3019,3027|false|false|false|C2136686|reported bruising (history)|bruising
Anatomy|Body Part, Organ, or Organ Component|General Exam|3035,3044|false|false|false|C0229118|Structure of both eyes|both eyes
Anatomy|Body Part, Organ, or Organ Component|General Exam|3040,3044|false|false|false|C0015392|Eye|eyes
Attribute|Clinical Attribute|General Exam|3040,3044|false|false|false|C5848506||eyes
Finding|Finding|General Exam|3046,3053|false|false|false|C0038999|Swelling|swollen
Finding|Finding|General Exam|3046,3058|false|false|false|C0240577|Swollen nose|swollen nose
Finding|Intellectual Product|General Exam|3064,3068|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Mental Process|General Exam|3069,3079|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3069,3079|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Activity|General Exam|3098,3103|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|3098,3103|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3098,3103|false|false|false|C1533810||place
Anatomy|Body Location or Region|General Exam|3106,3110|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3106,3110|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3106,3110|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|General Exam|3112,3118|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3128,3131|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3128,3131|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|General Exam|3128,3131|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Attribute|Clinical Attribute|General Exam|3134,3138|false|false|false|C0231832|Respiratory rate|RESP
Disorder|Disease or Syndrome|General Exam|3134,3138|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|RESP
Drug|Amino Acid, Peptide, or Protein|General Exam|3150,3153|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|General Exam|3150,3153|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|3150,3153|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|3197,3200|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|3197,3200|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Disorder|Disease or Syndrome|General Exam|3202,3206|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Disorder|Congenital Abnormality|General Exam|3248,3251|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Finding|Gene or Genome|General Exam|3248,3251|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Finding|Finding|General Exam|3253,3257|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3253,3257|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3259,3263|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|3277,3283|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3277,3283|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3277,3283|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|3288,3296|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|General Exam|3298,3306|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|3311,3316|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3311,3316|false|false|false|C0013604|Edema|edema
Finding|Finding|General Exam|3344,3350|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Functional Concept|General Exam|3352,3357|false|false|false|C1513492|motor movement|motor
Finding|Finding|General Exam|3352,3366|false|false|false|C5551447|Motor function (finding)|motor function
Phenomenon|Biologic Function|General Exam|3352,3366|false|false|false|C0234130|Motor function (observable entity)|motor function
Finding|Finding|General Exam|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|General Exam|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|General Exam|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|General Exam|3358,3366|false|false|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Anatomy|Body System|General Exam|3382,3386|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|General Exam|3382,3386|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|General Exam|3382,3386|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|General Exam|3382,3386|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|General Exam|3382,3386|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Disorder|Injury or Poisoning|General Exam|3391,3403|true|false|false|C0015256|Excoriation|excoriations
Disorder|Disease or Syndrome|General Exam|3407,3411|true|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|General Exam|3407,3411|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|General Exam|3407,3411|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Procedure|Health Care Activity|General Exam|3434,3443|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Disorder|Disease or Syndrome|General Exam|3457,3462|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3457,3462|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3463,3466|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3473,3476|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3473,3476|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3473,3476|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3483,3486|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3483,3486|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3483,3486|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3483,3486|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3492,3495|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3492,3495|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3502,3505|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3502,3505|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3502,3505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3502,3505|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3509,3512|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3509,3512|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3509,3512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3509,3512|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3509,3512|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3519,3523|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3539,3542|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3559,3564|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3559,3564|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3577,3583|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3589,3594|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3599,3602|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|3599,3602|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3629,3634|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3629,3634|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3639,3642|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|3639,3642|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3664,3669|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3664,3669|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3664,3677|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3664,3677|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3664,3677|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3670,3677|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3670,3677|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3670,3677|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3670,3677|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3670,3677|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3725,3729|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3725,3729|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3725,3729|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|3755,3760|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3755,3760|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3764,3767|false|false|false|C0010287|Creatine Kinase|CPK
Drug|Enzyme|General Exam|3764,3767|false|false|false|C0010287|Creatine Kinase|CPK
Finding|Gene or Genome|General Exam|3764,3767|false|false|false|C1418571|PIK3C2A gene|CPK
Procedure|Laboratory Procedure|General Exam|3764,3767|false|false|false|C0201973|Creatine kinase measurement|CPK
Anatomy|Body Part, Organ, or Organ Component|General Exam|3775,3782|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3775,3782|false|false|false|C1314974|Cardiac attachment|CARDIAC
Procedure|Laboratory Procedure|General Exam|3775,3789|false|false|false|C1271630|Cardiac markers|CARDIAC MARKER
Attribute|Clinical Attribute|General Exam|3790,3795|false|false|false|C4554533||TREND
Disorder|Disease or Syndrome|General Exam|3809,3814|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3809,3814|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|3841,3846|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3841,3846|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3847,3852|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3847,3852|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3847,3852|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3847,3852|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|3896,3901|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3896,3901|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3902,3907|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3902,3907|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3902,3907|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3902,3907|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|3950,3955|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3950,3955|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3956,3961|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3956,3961|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3956,3961|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3956,3961|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|3990,3995|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3990,3995|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3996,4001|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|3996,4001|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|3996,4001|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|3996,4001|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|General Exam|3999,4003|false|false|false|C0602256|MB 5|MB-5
Disorder|Disease or Syndrome|General Exam|4030,4035|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4030,4035|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4036,4041|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4036,4041|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4036,4041|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4036,4041|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|4070,4075|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4070,4075|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4076,4081|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|4076,4081|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|4076,4081|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|4076,4081|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Drug|Organic Chemical|General Exam|4079,4083|false|false|false|C0602249|MB 2|MB-2
Finding|Body Substance|General Exam|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4099,4108|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4099,4108|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|General Exam|4109,4113|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4127,4132|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4127,4132|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4133,4136|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4141,4144|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4141,4144|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4151,4154|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4151,4154|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4151,4154|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4151,4154|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4161,4164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4161,4164|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4172,4175|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4172,4175|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4172,4175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4172,4175|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4179,4182|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4179,4182|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4179,4182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4179,4182|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4179,4182|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4189,4193|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4208,4211|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4228,4233|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4228,4233|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4228,4241|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4228,4241|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4228,4241|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4234,4241|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4234,4241|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4234,4241|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4234,4241|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4234,4241|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4289,4293|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4289,4293|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4289,4293|false|false|false|C0202059|Bicarbonate measurement|HCO3
Finding|Finding|General Exam|4307,4314|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4307,4314|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Procedure|Diagnostic Procedure|General Exam|4320,4323|false|false|false|C0039985|Plain chest X-ray|CXR
Anatomy|Body Location or Region|General Exam|4352,4357|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|General Exam|4352,4357|false|false|false|C0741025|Chest problem|chest
Anatomy|Body Part, Organ, or Organ Component|General Exam|4372,4377|false|false|false|C0024109|Lung|lungs
Disorder|Disease or Syndrome|General Exam|4421,4434|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|General Exam|4442,4446|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4442,4451|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|General Exam|4442,4456|false|false|false|C0225732|Structure of base of left lung|left lung base
Anatomy|Body Location or Region|General Exam|4447,4451|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|4447,4451|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|4447,4451|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|4447,4451|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|4447,4456|false|false|false|C0225704|Basal segment of lung|lung base
Anatomy|Body Location or Region|General Exam|4452,4456|false|false|false|C2987514|Anatomical base|base
Drug|Biomedical or Dental Material|General Exam|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Chemical Viewed Functionally|General Exam|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4452,4456|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|base
Finding|Gene or Genome|General Exam|4452,4456|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Finding|Idea or Concept|General Exam|4452,4456|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|base
Anatomy|Body Part, Organ, or Organ Component|General Exam|4482,4495|false|false|false|C1269845|Structure of hemidiaphragm|hemidiaphragm
Finding|Intellectual Product|General Exam|4506,4510|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|4511,4519|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|General Exam|4521,4532|false|false|false|C0020452|Hyperemia|engorgement
Finding|Finding|General Exam|4521,4532|false|false|false|C1706102|Tick Engorgement|engorgement
Finding|Finding|General Exam|4553,4578|false|false|false|C5139173|Apical pulmonary opacity|apical pleural thickening
Anatomy|Tissue|General Exam|4560,4567|false|false|false|C0032225|Pleura|pleural
Disorder|Disease or Syndrome|General Exam|4560,4567|false|false|false|C0032226|Pleural Diseases|pleural
Disorder|Disease or Syndrome|General Exam|4560,4578|false|false|false|C0264545|Thickening of pleura|pleural thickening
Finding|Finding|General Exam|4568,4578|false|false|false|C0205400|Thickened|thickening
Anatomy|Body Part, Organ, or Organ Component|General Exam|4632,4638|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4632,4643|false|false|false|C0003489;C4037976|Aortic arch structure;Chest>Aortic arch|aortic arch
Disorder|Anatomical Abnormality|General Exam|4632,4643|false|false|false|C4759703|Aortic arch malformation|aortic arch
Anatomy|Body Location or Region|General Exam|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|4639,4643|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|4639,4643|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|4639,4643|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Finding|General Exam|4645,4659|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Finding|Organ or Tissue Function|General Exam|4645,4659|false|false|false|C0006660;C2242558|Pathologic calcification, calcified structure;Physiologic calcification|calcifications
Anatomy|Body Part, Organ, or Organ Component|General Exam|4665,4670|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|General Exam|4665,4670|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|General Exam|4665,4670|false|false|false|C0795691|HEART PROBLEM|heart
Procedure|Health Care Activity|General Exam|4700,4704|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|General Exam|4700,4704|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Finding|Functional Concept|General Exam|4709,4713|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4709,4720|false|false|false|C0225860|Left atrial structure|left atrium
Anatomy|Body Part, Organ, or Organ Component|General Exam|4714,4720|false|false|false|C0018792|Heart Atrium|atrium
Finding|Functional Concept|General Exam|4740,4744|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4740,4761|false|false|false|C0504053|Wall of left ventricle|Left ventricular wall
Anatomy|Body Part, Organ, or Organ Component|General Exam|4745,4756|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|4745,4761|false|false|false|C0507618|Wall of ventricle|ventricular wall
Anatomy|Body Space or Junction|General Exam|4779,4785|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|4779,4785|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|4779,4785|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Intellectual Product|General Exam|4812,4816|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|General Exam|4827,4831|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Disorder|Disease or Syndrome|General Exam|4827,4864|false|false|false|C1277187|Left ventricular systolic dysfunction|left ventricular systolic dysfunction
Anatomy|Body Part, Organ, or Organ Component|General Exam|4832,4843|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|General Exam|4844,4852|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|4844,4864|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|4853,4864|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|General Exam|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|4853,4864|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Finding|General Exam|4884,4895|false|false|false|C0086439|Hypokinesia|hypokinesis
Attribute|Clinical Attribute|General Exam|4939,4943|false|false|false|C0428772|Left ventricular ejection fraction|LVEF
Procedure|Diagnostic Procedure|General Exam|4939,4943|false|false|false|C3837267|LVEF (procedure)|LVEF
Finding|Pathologic Function|General Exam|4967,4974|true|false|false|C0087086|Thrombus|thrombi
Finding|Functional Concept|General Exam|4991,4995|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4991,5005|false|false|false|C0225897;C4266612|Chest>Heart.ventricle.left;Left ventricular structure|left ventricle
Anatomy|Body Part, Organ, or Organ Component|General Exam|4996,5005|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Anatomy|Body Space or Junction|General Exam|4996,5005|false|false|false|C0007799;C0018827;C2355627|Cerebral Ventricles;Heart Ventricle;Ventricle|ventricle
Finding|Functional Concept|General Exam|5007,5012|false|false|false|C1552823|Table Cell Horizontal Align - right|Right
Anatomy|Body Part, Organ, or Organ Component|General Exam|5014,5025|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Part, Organ, or Organ Component|General Exam|5026,5033|false|false|false|C0935616|chamber [body part]|chamber
Finding|Functional Concept|General Exam|5043,5047|false|false|false|C0332296|Free of (attribute)|free
Attribute|Clinical Attribute|General Exam|5048,5059|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|General Exam|5053,5059|false|false|false|C0026597|Motion|motion
Anatomy|Body Part, Organ, or Organ Component|General Exam|5089,5095|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5089,5101|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5096,5101|false|false|false|C1186983|Anatomical valve|valve
Finding|Intellectual Product|General Exam|5121,5125|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|5126,5132|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5126,5138|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5133,5138|false|false|false|C1186983|Anatomical valve|valve
Finding|Pathologic Function|General Exam|5140,5148|false|false|false|C1261287|Stenosis|stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5150,5155|false|false|false|C1186983|Anatomical valve|valve
Finding|Finding|General Exam|5150,5160|false|false|false|C4687749|Valve Area|valve area
Event|Governmental or Regulatory Activity|General Exam|5156,5160|false|false|false|C1510751|Academic Research Enhancement Awards|area
Disorder|Congenital Abnormality|General Exam|5164,5167|false|false|false|C0555206|Chiari malformation type II|cm2
Finding|Intellectual Product|General Exam|5170,5174|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|5180,5186|false|false|false|C0003483|Aorta|aortic
Disorder|Disease or Syndrome|General Exam|5180,5200|false|false|false|C0003504|Aortic Valve Insufficiency|aortic regurgitation
Finding|Finding|General Exam|5187,5200|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5187,5200|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5187,5200|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5215,5227|false|false|false|C0026264|Mitral Valve|mitral valve
Anatomy|Body Part, Organ, or Organ Component|General Exam|5222,5227|false|false|false|C1186983|Anatomical valve|valve
Disorder|Disease or Syndrome|General Exam|5268,5288|false|false|false|C0026266|Mitral Valve Insufficiency|mitral regurgitation
Finding|Finding|General Exam|5275,5288|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5275,5288|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5275,5288|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|General Exam|5302,5311|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|General Exam|5302,5311|false|false|false|C2707265||pulmonary
Finding|Finding|General Exam|5302,5311|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Anatomy|Body Part, Organ, or Organ Component|General Exam|5302,5318|false|false|false|C0034052|Pulmonary artery structure|pulmonary artery
Anatomy|Body Part, Organ, or Organ Component|General Exam|5312,5318|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|General Exam|5312,5318|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Organ or Tissue Function|General Exam|5319,5327|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|5329,5337|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|General Exam|5329,5337|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|General Exam|5329,5337|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|General Exam|5329,5337|false|false|false|C0033095||pressure
Finding|Functional Concept|General Exam|5382,5393|false|false|false|C0205463|Physiological|physiologic
Anatomy|Body Location or Region|General Exam|5395,5406|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|General Exam|5395,5406|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|General Exam|5395,5415|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|General Exam|5395,5415|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Finding|Body Substance|General Exam|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|General Exam|5407,5415|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|General Exam|5419,5429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|General Exam|5419,5429|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Functional Concept|General Exam|5438,5442|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Space or Junction|General Exam|5438,5461|false|false|false|C0503990|Cavity of left ventricle|left ventricular cavity
Attribute|Clinical Attribute|General Exam|5438,5466|false|false|false|C0455830|Left ventricular cavity size|left ventricular cavity size
Anatomy|Body Part, Organ, or Organ Component|General Exam|5443,5454|false|false|false|C0018827|Heart Ventricle|ventricular
Anatomy|Body Space or Junction|General Exam|5443,5461|false|false|false|C0507083|Cavity of ventricle|ventricular cavity
Anatomy|Body Space or Junction|General Exam|5455,5461|false|false|false|C0333343|Body cavities|cavity
Disorder|Anatomical Abnormality|General Exam|5455,5461|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Disorder|Disease or Syndrome|General Exam|5455,5461|false|false|false|C0011334;C1510420|Cavitation;Dental caries|cavity
Finding|Intellectual Product|General Exam|5472,5476|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Organ or Tissue Function|General Exam|5487,5495|false|false|false|C0039155|Systole|systolic
Finding|Pathologic Function|General Exam|5487,5507|false|false|false|C0749225|Systolic dysfunction|systolic dysfunction
Disorder|Disease or Syndrome|General Exam|5496,5507|false|false|false|C3887505|DYSFUNCTION - SKIN DISORDERS|dysfunction
Finding|Conceptual Entity|General Exam|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Functional Concept|General Exam|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Finding|Pathologic Function|General Exam|5496,5507|false|false|false|C0031847;C0277785;C3887504|Dysfunction;Functional disorder;physiopathological|dysfunction
Disorder|Disease or Syndrome|General Exam|5517,5520|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|General Exam|5517,5520|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|General Exam|5517,5520|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|General Exam|5517,5520|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|General Exam|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|General Exam|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|General Exam|5517,5520|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Attribute|Clinical Attribute|General Exam|5522,5528|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|General Exam|5529,5532|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|5529,5532|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|General Exam|5529,5532|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Cell Function|General Exam|5534,5546|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|General Exam|5534,5546|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Intellectual Product|General Exam|5549,5553|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Disorder|Disease or Syndrome|General Exam|5549,5575|false|false|false|C3276923|Mild aortic valve stenosis|Mild aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5554,5560|false|false|false|C0003483|Aorta|aortic
Anatomy|Body Part, Organ, or Organ Component|General Exam|5554,5566|false|false|false|C0003501;C4533215|Aortic valve structure;Chest>Aortic valve|aortic valve
Disorder|Congenital Abnormality|General Exam|5554,5575|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Disorder|Disease or Syndrome|General Exam|5554,5575|false|false|false|C5193127;C5700069|AORTIC VALVE DISEASE 3;Stenosis of aorta|aortic valve stenosis
Finding|Pathologic Function|General Exam|5554,5575|false|false|false|C0003507|Aortic Valve Stenosis|aortic valve stenosis
Anatomy|Body Part, Organ, or Organ Component|General Exam|5561,5566|false|false|false|C1186983|Anatomical valve|valve
Finding|Pathologic Function|General Exam|5567,5575|false|false|false|C1261287|Stenosis|stenosis
Finding|Intellectual Product|General Exam|5577,5581|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Anatomy|Body Part, Organ, or Organ Component|General Exam|5582,5588|false|false|false|C0003483|Aorta|aortic
Finding|Finding|General Exam|5590,5603|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|General Exam|5590,5603|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|General Exam|5590,5603|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Finding|Conceptual Entity|Hospital Course|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5654,5661|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5654,5664|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|Hospital Course|5665,5668|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Hospital Course|5665,5668|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Hospital Course|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Hospital Course|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Hospital Course|5665,5668|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Finding|Gene or Genome|Hospital Course|5665,5668|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Finding|Functional Concept|Hospital Course|5673,5679|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Hospital Course|5673,5679|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Hospital Course|5673,5679|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5673,5679|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|Hospital Course|5700,5712|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Hospital Course|5718,5732|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Finding|Finding|Hospital Course|5718,5732|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5753,5758|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|5753,5758|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|5753,5758|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|5753,5758|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|Hospital Course|5759,5768|false|false|false|C0016658|Fracture|fractures
Finding|Finding|Hospital Course|5759,5768|false|false|false|C4554413|Fractured|fractures
Finding|Pathologic Function|Hospital Course|5773,5782|false|false|false|C0014591|Epistaxis|epistaxis
Finding|Functional Concept|Hospital Course|5789,5799|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5789,5799|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|Hospital Course|5801,5805|false|false|false|C0085639|Falls|fall
Finding|Idea or Concept|Hospital Course|5811,5819|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|Hospital Course|5811,5826|false|false|false|C0488549||hospital course
Finding|Finding|Hospital Course|5811,5826|false|false|false|C0489547|Hospital course|hospital course
Disorder|Disease or Syndrome|Hospital Course|5842,5848|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|5842,5848|false|false|false|C3537184||NSTEMI
Finding|Pathologic Function|Hospital Course|5852,5861|false|false|false|C0014591|Epistaxis|Epistaxis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5863,5868|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|5863,5868|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|5863,5868|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|5863,5868|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|Hospital Course|5869,5878|false|false|false|C0016658|Fracture|fractures
Finding|Finding|Hospital Course|5869,5878|false|false|false|C4554413|Fractured|fractures
Finding|Body Substance|Hospital Course|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|5879,5886|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|Hospital Course|5904,5914|false|false|false|C0443254|mechanical method|mechanical
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5904,5914|false|false|false|C0699886|Mechanical Treatments|mechanical
Finding|Finding|Hospital Course|5915,5919|false|false|false|C0085639|Falls|fall
Finding|Idea or Concept|Hospital Course|5957,5965|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Hospital Course|5970,5977|false|false|false|C0549178|Continuous|ongoing
Finding|Pathologic Function|Hospital Course|5978,5987|false|false|false|C0014591|Epistaxis|epistaxis
Procedure|Diagnostic Procedure|Hospital Course|5989,5996|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|Hospital Course|5992,5996|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Idea or Concept|Hospital Course|6008,6016|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6030,6035|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|6030,6035|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|6030,6035|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|6030,6035|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6030,6040|false|false|false|C0027422|Nasal bone structure|nasal bone
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6036,6040|false|false|false|C0262950;C1442209|Skeletal bone;XXX bone|bone
Finding|Body Substance|Hospital Course|6036,6040|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Finding|Intellectual Product|Hospital Course|6036,6040|false|false|false|C1546560;C1550616|Specimen Type - Bone|bone
Disorder|Injury or Poisoning|Hospital Course|6052,6061|false|false|false|C0016658|Fracture|fractures
Finding|Finding|Hospital Course|6052,6061|false|false|false|C4554413|Fractured|fractures
Finding|Idea or Concept|Hospital Course|6103,6112|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|6103,6112|false|false|false|C1555324|inpatient encounter|inpatient
Finding|Body Substance|Hospital Course|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6140,6149|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6140,6149|false|false|false|C0030685|Patient Discharge|discharge
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6190,6195|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|6190,6195|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|6190,6195|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|6190,6195|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Biomedical or Dental Material|Hospital Course|6197,6202|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|6197,6202|false|false|false|C2003858|Spray (action)|spray
Finding|Functional Concept|Hospital Course|6197,6202|false|false|false|C4521772|Spray (administration method)|spray
Event|Activity|Hospital Course|6207,6211|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|Hospital Course|6207,6211|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|Hospital Course|6207,6211|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Finding|Hospital Course|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Hospital Course|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Hospital Course|6212,6220|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Hospital Course|6212,6220|false|false|false|C0033095||pressure
Finding|Pathologic Function|Hospital Course|6228,6236|false|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|Hospital Course|6249,6255|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|6249,6255|false|false|false|C3537184||NSTEMI
Finding|Body Substance|Hospital Course|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6256,6263|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6278,6282|false|false|false|C1547225|Mild Severity of Illness Code|mild
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6283,6292|false|false|false|C0439775|Elevation procedure|elevation
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6296,6304|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Hospital Course|6296,6304|false|false|false|C0041199|Troponin|troponin
Procedure|Laboratory Procedure|Hospital Course|6296,6304|false|false|false|C0523952|Troponin measurement|troponin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6372,6381|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|6372,6381|false|false|false|C1179435|Protein Component|component
Finding|Conceptual Entity|Hospital Course|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|6372,6381|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Procedure|Health Care Activity|Hospital Course|6412,6421|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Body Substance|Hospital Course|6427,6434|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6427,6434|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6427,6434|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Body Location or Region|Hospital Course|6448,6453|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|6448,6453|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|6448,6458|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|6448,6458|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|6454,6458|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6454,6458|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6454,6458|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6468,6475|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|6468,6475|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Sign or Symptom|Hospital Course|6468,6484|false|false|false|C0741933|cardiac symptom|cardiac symptoms
Finding|Functional Concept|Hospital Course|6476,6484|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|6476,6484|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body System|Hospital Course|6486,6496|false|false|false|C0007226|Cardiovascular system|Cardiology
Finding|Idea or Concept|Hospital Course|6538,6549|false|false|false|C0750501|most likely|most likely
Finding|Finding|Hospital Course|6543,6549|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6543,6549|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|Hospital Course|6550,6559|false|true|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|6550,6559|false|true|false|C1522484|metastatic qualifier|secondary
Finding|Idea or Concept|Hospital Course|6563,6569|false|false|false|C0699784|Economic demand|demand
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6563,6569|false|false|false|C0441516|Demand (clinical)|demand
Finding|Pathologic Function|Hospital Course|6571,6579|false|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6571,6579|false|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Gene or Genome|Hospital Course|6581,6585|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Hospital Course|6581,6585|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Disorder|Neoplastic Process|Hospital Course|6593,6602|false|false|false|C0027627|Neoplasm Metastasis|secondary
Finding|Functional Concept|Hospital Course|6593,6602|false|false|false|C1522484|metastatic qualifier|secondary
Finding|Finding|Hospital Course|6610,6614|false|false|false|C0085639|Falls|fall
Procedure|Diagnostic Procedure|Hospital Course|6619,6633|false|false|false|C0013516|Echocardiography|echocardiogram
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6648,6654|false|false|false|C0003483|Aorta|aortic
Finding|Pathologic Function|Hospital Course|6648,6663|false|false|false|C0003507|Aortic Valve Stenosis|aortic stenosis
Finding|Pathologic Function|Hospital Course|6655,6663|false|false|false|C1261287|Stenosis|stenosis
Finding|Finding|Hospital Course|6668,6674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6668,6674|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Attribute|Clinical Attribute|Hospital Course|6675,6681|false|true|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6682,6685|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|6682,6685|false|true|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|6682,6685|false|true|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Hospital Course|6686,6693|false|true|false|C0012634|Disease|disease
Attribute|Clinical Attribute|Hospital Course|6704,6715|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|Hospital Course|6709,6715|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|Hospital Course|6716,6729|false|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|Hospital Course|6716,6729|false|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|Hospital Course|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6735,6742|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|6745,6755|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|6745,6755|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|6777,6788|false|false|false|C0085542|pravastatin|pravastatin
Drug|Pharmacologic Substance|Hospital Course|6777,6788|false|false|false|C0085542|pravastatin|pravastatin
Drug|Organic Chemical|Hospital Course|6806,6818|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|6806,6818|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Organic Chemical|Hospital Course|6825,6836|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|6825,6836|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Organic Chemical|Hospital Course|6875,6882|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|6875,6882|false|false|false|C0004057|aspirin|aspirin
Finding|Finding|Hospital Course|6886,6895|false|false|false|C0700292;C5548348|Blood oxygen concentration below reference range (finding);Hypoxemia|Hypoxemia
Disorder|Disease or Syndrome|Hospital Course|6906,6919|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Body Substance|Hospital Course|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6920,6927|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Pathologic Function|Hospital Course|6950,6957|false|false|false|C0242184|Hypoxia|hypoxic
Drug|Biologically Active Substance|Hospital Course|6998,7004|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Hospital Course|6998,7004|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Hospital Course|6998,7004|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6998,7004|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Attribute|Clinical Attribute|Hospital Course|6998,7016|false|false|false|C0483415|Oxygen Saturation|oxygen saturations
Phenomenon|Natural Phenomenon or Process|Hospital Course|7005,7016|false|false|false|C0522534|Saturated|saturations
Finding|Finding|Hospital Course|7017,7028|false|false|false|C2709070|on room air|on room air
Drug|Inorganic Chemical|Hospital Course|7020,7028|false|false|false|C3846005|Room Air|room air
Drug|Inorganic Chemical|Hospital Course|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|7025,7028|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Hospital Course|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|7025,7028|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Attribute|Clinical Attribute|Hospital Course|7041,7060|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|7041,7060|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|7054,7060|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|7064,7069|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|7064,7069|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|Hospital Course|7064,7069|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|Hospital Course|7071,7077|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|Hospital Course|7088,7098|false|false|false|C0009450|Communicable Diseases|infectious
Finding|Functional Concept|Hospital Course|7100,7108|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|7100,7108|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Disorder|Disease or Syndrome|Hospital Course|7120,7132|true|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|7120,7132|true|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Procedure|Diagnostic Procedure|Hospital Course|7136,7139|false|false|false|C0039985|Plain chest X-ray|CXR
Disorder|Disease or Syndrome|Hospital Course|7149,7162|false|false|false|C0521530|Lung consolidation|consolidation
Finding|Functional Concept|Hospital Course|7167,7171|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7167,7176|false|false|false|C0225730|Left lung|left lung
Anatomy|Body Location or Region|Hospital Course|7172,7176|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7172,7176|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|7172,7176|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|7172,7176|false|false|false|C0740941|Lung Problem|lung
Finding|Idea or Concept|Hospital Course|7178,7185|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|Hospital Course|7178,7185|false|false|false|C0039869;C4319827|Thought|thought
Finding|Finding|Hospital Course|7192,7200|false|false|false|C0332149|Possible|possibly
Drug|Organic Chemical|Hospital Course|7201,7208|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|7201,7208|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|7201,7208|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Injury or Poisoning|Hospital Course|7212,7221|false|false|false|C1720922|Respiratory Aspiration|aspirated
Finding|Organ or Tissue Function|Hospital Course|7212,7221|false|false|false|C0700198|Pulmonary aspiration|aspirated
Disorder|Disease or Syndrome|Hospital Course|7222,7227|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|7222,7227|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Hazardous or Poisonous Substance|Hospital Course|7231,7238|false|false|false|C0728873|Monitor brand of insecticide|monitor
Drug|Organic Chemical|Hospital Course|7231,7238|false|false|false|C0728873|Monitor brand of insecticide|monitor
Procedure|Laboratory Procedure|Hospital Course|7239,7252|false|false|false|C0523807|Oxygen saturation measurement|O2 saturation
Phenomenon|Natural Phenomenon or Process|Hospital Course|7242,7252|false|false|false|C0522534|Saturated|saturation
Procedure|Health Care Activity|Hospital Course|7254,7265|false|false|false|C0886414|Body temperature measurement|temperature
Attribute|Clinical Attribute|Hospital Course|7267,7272|false|false|false|C4554533||trend
Anatomy|Cell|Hospital Course|7273,7276|false|false|false|C0023516|Leukocytes|WBC
Drug|Antibiotic|Hospital Course|7300,7311|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Idea or Concept|Hospital Course|7318,7327|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|7318,7327|false|false|false|C1555324|inpatient encounter|inpatient
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7343,7354|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Finding|Body Substance|Hospital Course|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|7409,7418|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|7409,7418|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|Hospital Course|7422,7427|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|7422,7441|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Disorder|Injury or Poisoning|Hospital Course|7422,7441|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute kidney injury
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7428,7434|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|7428,7434|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|7428,7434|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|7428,7434|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7428,7434|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|Hospital Course|7428,7441|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|Hospital Course|7435,7441|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Finding|Body Substance|Hospital Course|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7442,7449|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|Hospital Course|7465,7475|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|7465,7475|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|Hospital Course|7465,7475|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|7465,7475|false|false|false|C0201975|Creatinine measurement|creatinine
Drug|Biologically Active Substance|Hospital Course|7493,7503|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|7493,7503|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|Hospital Course|7493,7503|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|7493,7503|false|false|false|C0201975|Creatinine measurement|creatinine
Disorder|Disease or Syndrome|Hospital Course|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|7508,7511|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|7508,7511|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|7508,7511|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|7508,7511|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|Hospital Course|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7517,7524|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Procedure|Research Activity|Hospital Course|7529,7536|false|false|false|C0150114|unaware|unaware
Finding|Conceptual Entity|Hospital Course|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7542,7549|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7542,7552|false|false|false|C0262926|Medical History|history of
Finding|Finding|Hospital Course|7542,7567|false|false|false|C0455686||history of kidney disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7553,7559|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|7553,7559|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|7553,7559|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|7553,7559|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7553,7559|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|7553,7567|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|7560,7567|false|false|false|C0012634|Disease|disease
Finding|Body Substance|Hospital Course|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7574,7581|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|7604,7610|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Biologically Active Substance|Hospital Course|7611,7621|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|7611,7621|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|Hospital Course|7611,7621|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|7611,7621|false|false|false|C0201975|Creatinine measurement|creatinine
Disorder|Disease or Syndrome|Hospital Course|7625,7652|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7636,7644|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|Hospital Course|7636,7652|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|Hospital Course|7645,7652|false|false|false|C0012634|Disease|disease
Finding|Body Substance|Hospital Course|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7653,7660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Conceptual Entity|Hospital Course|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7667,7674|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7667,7677|false|false|false|C0262926|Medical History|history of
Disorder|Anatomical Abnormality|Hospital Course|7678,7681|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Disorder|Disease or Syndrome|Hospital Course|7678,7681|false|false|false|C0003486;C0162871|Aortic Aneurysm;Aortic Aneurysm, Abdominal|AAA
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7678,7681|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Biologically Active Substance|Hospital Course|7678,7681|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Organic Chemical|Hospital Course|7678,7681|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Drug|Pharmacologic Substance|Hospital Course|7678,7681|false|false|false|C0611285;C0731345|AAA brand of benzocaine-cetalkonium chloride combination;APP protein, human|AAA
Finding|Gene or Genome|Hospital Course|7678,7681|false|false|false|C1364818;C1705543;C5780959|AAAS wt Allele;APP gene;APP wt Allele|AAA
Finding|Functional Concept|Hospital Course|7682,7688|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Hospital Course|7682,7688|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Hospital Course|7682,7688|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7682,7688|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Finding|Conceptual Entity|Hospital Course|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7704,7711|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7704,7714|true|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|7723,7726|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7723,7726|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|7723,7726|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7723,7726|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|7723,7726|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|7723,7726|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|7723,7726|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|7723,7726|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|7723,7726|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|7723,7726|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Body Substance|Hospital Course|7728,7735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7728,7735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7728,7735|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Conceptual Entity|Hospital Course|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7743,7750|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7743,7753|false|false|false|C0262926|Medical History|history of
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7754,7758|true|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7762,7769|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|7762,7769|true|false|false|C1314974|Cardiac attachment|cardiac
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7792,7799|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Hospital Course|7792,7799|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Intellectual Product|Hospital Course|7800,7807|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7800,7807|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Idea or Concept|Hospital Course|7826,7831|false|false|false|C1552828|Table Frame - above|above
Finding|Idea or Concept|Hospital Course|7834,7846|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Classification|Hospital Course|7855,7865|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|7855,7865|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Attribute|Clinical Attribute|Hospital Course|7866,7872|false|false|false|C1718621|W stress|stress
Drug|Organic Chemical|Hospital Course|7866,7872|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Hospital Course|7866,7872|false|false|false|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Hospital Course|7866,7872|false|false|false|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Hospital Course|7866,7877|false|false|false|C0920208|Echocardiography, Stress|stress echo
Procedure|Health Care Activity|Hospital Course|7873,7877|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7873,7877|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Idea or Concept|Hospital Course|7889,7899|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|7889,7899|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Attribute|Clinical Attribute|Hospital Course|7900,7906|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7907,7910|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|Hospital Course|7907,7910|false|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|Hospital Course|7907,7910|false|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Disorder|Disease or Syndrome|Hospital Course|7911,7918|false|false|false|C0012634|Disease|disease
Finding|Finding|Hospital Course|7921,7929|false|false|false|C0332149|Possible|possibly
Finding|Gene or Genome|Hospital Course|7932,7937|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Tissue|Hospital Course|7938,7948|false|false|false|C0027061|Myocardium|myocardial
Finding|Idea or Concept|Hospital Course|7962,7966|false|false|false|C0035647|Risk|risk
Finding|Functional Concept|Hospital Course|7971,7977|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Procedure|Diagnostic Procedure|Hospital Course|7978,7992|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Intellectual Product|Hospital Course|8017,8021|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Pathologic Function|Hospital Course|8033,8042|false|false|false|C0014591|Epistaxis|epistaxis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8074,8079|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8074,8079|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8074,8079|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8074,8079|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Drug|Pharmacologic Substance|Hospital Course|8074,8085|false|false|false|C2608294|Nasal Spray brand of phenylephrine|nasal spray
Drug|Biomedical or Dental Material|Hospital Course|8080,8085|false|false|false|C1154182|Spray Dosage Form|spray
Event|Activity|Hospital Course|8080,8085|false|false|false|C2003858|Spray (action)|spray
Finding|Functional Concept|Hospital Course|8080,8085|false|false|false|C4521772|Spray (administration method)|spray
Finding|Functional Concept|Hospital Course|8088,8094|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Anatomy|Body Location or Region|Hospital Course|8095,8100|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|8095,8100|false|false|false|C0741025|Chest problem|chest
Procedure|Diagnostic Procedure|Hospital Course|8095,8106|false|false|false|C0039985|Plain chest X-ray|chest x-ray
Finding|Functional Concept|Hospital Course|8101,8106|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Finding|Intellectual Product|Hospital Course|8101,8106|false|false|false|C0034571;C3244296|ActClaimAttachmentCategoryCode - x-ray;roentgenographic|x-ray
Phenomenon|Natural Phenomenon or Process|Hospital Course|8101,8106|false|false|false|C0043309|Roentgen Rays|x-ray
Procedure|Diagnostic Procedure|Hospital Course|8101,8106|false|false|false|C0043299;C1306645;C1962945|Diagnostic radiologic examination;Plain x-ray;Radiographic imaging procedure|x-ray
Finding|Conceptual Entity|Hospital Course|8130,8140|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Finding|Pathologic Function|Hospital Course|8130,8140|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|resolution
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8148,8151|false|false|false|C1261077|Structure of left lower lobe of lung|LLL
Finding|Finding|Hospital Course|8153,8165|false|false|false|C4527217|Infiltrative Tumor Margin|infiltrative
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8166,8173|false|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|Hospital Course|8166,8173|false|false|false|C1951340|Process Pharmacologic Substance|process
Finding|Functional Concept|Hospital Course|8166,8173|false|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|Hospital Course|8166,8173|false|false|false|C1522240|Process|process
Finding|Idea or Concept|Hospital Course|8176,8184|false|false|false|C0750591|consider|Consider
Finding|Functional Concept|Hospital Course|8185,8191|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|8185,8191|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|8185,8194|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|8185,8194|false|false|false|C1522577|follow-up|follow-up
Anatomy|Body Location or Region|Hospital Course|8200,8203|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8200,8203|false|false|false|C0150934;C0175196|Ear, nose and throat;Structure of entorhinal cortex|ENT
Finding|Gene or Genome|Hospital Course|8200,8203|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Finding|Sign or Symptom|Hospital Course|8200,8203|false|false|false|C0262471;C1417861;C3889152|ENT problem;NT5E gene;NT5E wt Allele|ENT
Drug|Substance|Hospital Course|8207,8214|false|false|false|C0032167|Plastics|Plastic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8207,8222|false|false|false|C0677616|Plastic Surgical Procedures|Plastic Surgery
Finding|Finding|Hospital Course|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Functional Concept|Hospital Course|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Finding|Idea or Concept|Hospital Course|8215,8222|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|Surgery
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8215,8222|false|false|false|C0543467|Operative Surgical Procedures|Surgery
Finding|Idea or Concept|Hospital Course|8234,8244|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|8234,8244|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8248,8253|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|Hospital Course|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|Hospital Course|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|Hospital Course|8248,8253|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|Hospital Course|8248,8253|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|Hospital Course|8248,8253|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Disorder|Injury or Poisoning|Hospital Course|8254,8263|false|false|false|C0016658|Fracture|fractures
Finding|Finding|Hospital Course|8254,8263|false|false|false|C4554413|Fractured|fractures
Finding|Functional Concept|Hospital Course|8266,8272|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Anatomy|Cell Component|Hospital Course|8273,8276|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|8273,8276|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Intellectual Product|Hospital Course|8284,8288|false|false|false|C1561540|Transaction counts and value totals - week|week
Procedure|Laboratory Procedure|Hospital Course|8312,8315|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8312,8315|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|HCT
Anatomy|Cell|Hospital Course|8321,8330|false|false|false|C0005821|Blood Platelets|platelets
Drug|Pharmacologic Substance|Hospital Course|8321,8330|false|false|false|C0443116|Platelets Product|platelets
Procedure|Laboratory Procedure|Hospital Course|8321,8330|false|false|false|C0032181|Platelet count (procedure)|platelets
Finding|Idea or Concept|Hospital Course|8333,8341|false|false|false|C0750591|consider|Consider
Finding|Functional Concept|Hospital Course|8342,8352|false|false|false|C0439836|Conversions (qualifier value)|conversion
Drug|Organic Chemical|Hospital Course|8356,8366|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8356,8366|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|8356,8375|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|Hospital Course|8356,8375|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|Hospital Course|8367,8375|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|Hospital Course|8367,8375|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Organic Chemical|Hospital Course|8379,8388|false|false|false|C0038617;C0220918|Succinates;succinate|succinate
Finding|Mental Process|Hospital Course|8394,8398|false|false|false|C1331418|Comfort|ease
Event|Occupational Activity|Hospital Course|8402,8416|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8402,8416|false|false|false|C1533734|Administration (procedure)|administration
Attribute|Clinical Attribute|Hospital Course|8420,8431|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8420,8431|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8420,8431|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|8420,8444|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|8435,8444|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|8463,8473|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|8463,8473|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|8463,8478|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|8474,8478|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|8495,8503|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|8495,8503|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8495,8503|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|8508,8519|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|8508,8519|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|8539,8549|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|8539,8558|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|8550,8558|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Organic Chemical|Hospital Course|8576,8587|false|false|false|C0085542|pravastatin|Pravastatin
Drug|Pharmacologic Substance|Hospital Course|8576,8587|false|false|false|C0085542|pravastatin|Pravastatin
Finding|Body Substance|Hospital Course|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|8605,8614|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|8605,8614|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|8605,8626|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|8615,8626|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|8615,8626|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|8615,8626|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|8631,8642|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|8631,8642|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|8662,8675|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8662,8675|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8662,8675|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8690,8693|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8694,8698|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|8694,8698|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|8694,8698|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|8713,8718|false|false|false|C0003211;C3536840|Anti-Inflammatory Agents, Non-Steroidal|NSAID
Attribute|Clinical Attribute|Hospital Course|8719,8730|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|8719,8730|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|8719,8730|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Hospital Course|8736,8745|false|false|false|C0020740|ibuprofen|ibuprofen
Drug|Pharmacologic Substance|Hospital Course|8736,8745|false|false|false|C0020740|ibuprofen|ibuprofen
Finding|Pathologic Function|Hospital Course|8758,8766|false|false|false|C0019080|Hemorrhage|bleeding
Drug|Organic Chemical|Hospital Course|8772,8779|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8772,8779|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8795,8803|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Drug|Organic Chemical|Hospital Course|8817,8827|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Pharmacologic Substance|Hospital Course|8817,8827|false|false|false|C0025859|metoprolol|Metoprolol
Drug|Organic Chemical|Hospital Course|8817,8836|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Pharmacologic Substance|Hospital Course|8817,8836|false|false|false|C0700548|metoprolol tartrate|Metoprolol Tartrate
Drug|Organic Chemical|Hospital Course|8828,8836|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Pharmacologic Substance|Hospital Course|8828,8836|false|false|false|C0039328;C0144544|Tartrates;tartrate|Tartrate
Drug|Organic Chemical|Hospital Course|8855,8865|false|false|false|C0025859|metoprolol|metoprolol
Drug|Pharmacologic Substance|Hospital Course|8855,8865|false|false|false|C0025859|metoprolol|metoprolol
Drug|Organic Chemical|Hospital Course|8855,8874|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Pharmacologic Substance|Hospital Course|8855,8874|false|false|false|C0700548|metoprolol tartrate|metoprolol tartrate
Drug|Organic Chemical|Hospital Course|8866,8874|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Pharmacologic Substance|Hospital Course|8866,8874|false|false|false|C0039328;C0144544|Tartrates;tartrate|tartrate
Drug|Biomedical or Dental Material|Hospital Course|8883,8889|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|8893,8901|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|8896,8901|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|8896,8901|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Disorder|Disease or Syndrome|Hospital Course|8908,8913|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Drug|Biomedical or Dental Material|Hospital Course|8932,8938|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|8939,8946|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|8953,8965|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8953,8965|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|8984,8996|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8984,8996|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Biomedical or Dental Material|Hospital Course|9005,9011|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Hospital Course|9015,9023|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|9018,9023|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|9018,9023|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|9038,9042|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|9038,9042|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|9049,9055|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|9056,9063|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|9070,9083|false|false|false|C0030071|oxymetazoline|Oxymetazoline
Drug|Pharmacologic Substance|Hospital Course|9070,9083|false|false|false|C0030071|oxymetazoline|Oxymetazoline
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9094,9097|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9094,9097|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9094,9097|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9094,9097|false|false|false|C1332410|BID gene|BID
Finding|Gene or Genome|Hospital Course|9098,9101|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Hazardous or Poisonous Substance|Hospital Course|9144,9151|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Hospital Course|9144,9151|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Intellectual Product|Hospital Course|9157,9167|false|false|false|C0592503|Proprietary Name|brand name
Finding|Intellectual Product|Hospital Course|9163,9167|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Finding|Body Substance|Hospital Course|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9181,9190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9181,9190|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|9181,9202|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|9181,9202|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|9191,9202|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|9191,9202|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|Hospital Course|9204,9208|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9204,9208|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9204,9208|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|9214,9221|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|9214,9221|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Finding|Intellectual Product|Hospital Course|9224,9232|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9240,9249|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9240,9249|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9240,9259|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|9250,9259|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|9250,9259|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|9250,9259|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|9250,9259|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9261,9266|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|Hospital Course|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|Hospital Course|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|Hospital Course|9261,9266|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|Hospital Course|9261,9266|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|Hospital Course|9261,9266|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Disorder|Injury or Poisoning|Hospital Course|9261,9275|false|false|false|C0339848|Fractured nasal bones|Nasal fracture
Disorder|Injury or Poisoning|Hospital Course|9267,9275|false|false|false|C0016658|Fracture|fracture
Finding|Pathologic Function|Hospital Course|9276,9285|false|false|false|C0014591|Epistaxis|Epistaxis
Disorder|Disease or Syndrome|Hospital Course|9286,9292|false|false|false|C4255010||NSTEMI
Finding|Finding|Hospital Course|9286,9292|false|false|false|C3537184||NSTEMI
Finding|Mental Process|Discharge Condition|9317,9323|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9317,9330|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9317,9330|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9324,9330|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9324,9330|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|9332,9337|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|9342,9350|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|9352,9374|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9352,9374|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|9361,9374|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9361,9374|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9376,9381|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9376,9381|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9376,9381|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9376,9381|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9386,9397|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9399,9407|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9399,9407|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9399,9407|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9408,9414|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9408,9414|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9416,9426|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9416,9426|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|Discharge Condition|9429,9440|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|9429,9440|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Pathologic Function|Discharge Instructions|9546,9552|false|false|false|C0019080|Hemorrhage|bleeds
Finding|Finding|Discharge Instructions|9563,9572|false|false|false|C0332218|Difficult (qualifier value)|difficult
Finding|Pathologic Function|Discharge Instructions|9634,9642|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Idea or Concept|Discharge Instructions|9656,9664|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|Discharge Instructions|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Discharge Instructions|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Discharge Instructions|9697,9701|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|9702,9711|false|false|false|C0041199|Troponin|troponins
Drug|Biologically Active Substance|Discharge Instructions|9702,9711|false|false|false|C0041199|Troponin|troponins
Disorder|Disease or Syndrome|Discharge Instructions|9715,9720|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|9715,9720|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Laboratory Procedure|Discharge Instructions|9715,9725|false|false|false|C0018941|Hematologic Tests|blood test
Anatomy|Body Location or Region|Discharge Instructions|9721,9725|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Discharge Instructions|9721,9725|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|9721,9725|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|9721,9725|false|false|false|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|9721,9725|false|false|false|C0022885|Laboratory Procedures|test
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9735,9740|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|9735,9740|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|9735,9740|false|false|false|C0795691|HEART PROBLEM|heart
Finding|Functional Concept|Discharge Instructions|9744,9754|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|9744,9754|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Discharge Instructions|9744,9754|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|9763,9768|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|Discharge Instructions|9763,9768|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|Discharge Instructions|9763,9768|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Disease or Syndrome|Discharge Instructions|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Discharge Instructions|9816,9819|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Discharge Instructions|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Discharge Instructions|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Discharge Instructions|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Discharge Instructions|9816,9819|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Discharge Instructions|9816,9819|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Discharge Instructions|9816,9819|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|Discharge Instructions|9831,9837|false|false|true|C1718621|W stress|stress
Drug|Organic Chemical|Discharge Instructions|9831,9837|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Drug|Pharmacologic Substance|Discharge Instructions|9831,9837|false|false|true|C0723460|Stress bismuth subsalicylate|stress
Finding|Finding|Discharge Instructions|9831,9837|false|false|true|C0038435|Stress|stress
Procedure|Diagnostic Procedure|Discharge Instructions|9831,9842|false|false|true|C0015260;C3494508|Exercise stress test;Stress Test|stress test
Anatomy|Body Location or Region|Discharge Instructions|9838,9842|false|false|false|C4318744|Test - temporal region|test
Finding|Functional Concept|Discharge Instructions|9838,9842|false|false|true|C0039593;C0392366|Testing;Tests (qualifier value)|test
Finding|Intellectual Product|Discharge Instructions|9838,9842|false|false|true|C0039593;C0392366|Testing;Tests (qualifier value)|test
Lab|Laboratory or Test Result|Discharge Instructions|9838,9842|false|false|true|C0456984|Test Result|test
Procedure|Laboratory Procedure|Discharge Instructions|9838,9842|false|false|true|C0022885|Laboratory Procedures|test
Finding|Intellectual Product|Discharge Instructions|9854,9862|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|9854,9862|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|9885,9889|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|9885,9889|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|9885,9889|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Activity|Discharge Instructions|9906,9914|false|false|false|C1707391|Choose (action)|choosing
Procedure|Health Care Activity|Discharge Instructions|9922,9930|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|9931,9943|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|9931,9943|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

