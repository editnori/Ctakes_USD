 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|155,163|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|166,175|false|false|false|C1717415||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|166,175|false|false|false|C0020517|Hypersensitivity|Allergies
Drug|Organic Chemical|SIMPLE_SEGMENT|178,185|false|false|false|C0009214|codeine|Codeine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|178,185|false|false|false|C0009214|codeine|Codeine
Drug|Antibiotic|SIMPLE_SEGMENT|188,197|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|SIMPLE_SEGMENT|188,197|false|false|false|C0591132|Augmentin|Augmentin
Drug|Organic Chemical|SIMPLE_SEGMENT|200,207|false|false|false|C0723778|Topamax|Topamax
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|200,207|false|false|false|C0723778|Topamax|Topamax
Finding|Functional Concept|SIMPLE_SEGMENT|210,219|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|228,243|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|234,243|false|false|false|C3864418||Complaint
Finding|Finding|SIMPLE_SEGMENT|234,243|false|false|false|C5441521|Complaint (finding)|Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|245,264|false|false|false|C2707305||Shortness of Breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|245,264|false|false|false|C0013404|Dyspnea|Shortness of Breath
Finding|Body Substance|SIMPLE_SEGMENT|258,264|false|false|false|C0225386|Breath|Breath
Finding|Classification|SIMPLE_SEGMENT|267,272|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|273,281|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|273,281|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|285,303|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|294,303|false|false|false|C0945766||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|294,303|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|294,303|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|294,303|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Conceptual Entity|SIMPLE_SEGMENT|313,320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|313,320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|313,320|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|313,323|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|313,339|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|313,339|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|324,331|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|324,331|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|324,339|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|332,339|false|false|false|C0221423|Illness (finding)|Illness
Finding|Conceptual Entity|SIMPLE_SEGMENT|363,370|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|363,370|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|363,370|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|363,373|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|363,391|false|false|false|C5192533|History of cerebral aneurysm|history of cerebral aneurysm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|374,382|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|374,391|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|383,391|false|false|false|C0002940|Aneurysm|aneurysm
Attribute|Clinical Attribute|SIMPLE_SEGMENT|410,429|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|410,429|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|423,429|false|false|false|C0225386|Breath|breath
Event|Occupational Activity|SIMPLE_SEGMENT|490,500|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|490,500|false|false|false|C0376636|Disease Management|management
Finding|Idea or Concept|SIMPLE_SEGMENT|518,523|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|SIMPLE_SEGMENT|518,523|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Finding|SIMPLE_SEGMENT|538,546|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|538,546|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|SIMPLE_SEGMENT|559,565|false|false|false|C0392197;C0518610|Physiologic warmth;Social warmth|warmth
Finding|Physiologic Function|SIMPLE_SEGMENT|559,565|false|false|false|C0392197;C0518610|Physiologic warmth;Social warmth|warmth
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|570,578|false|false|false|C0041834|Erythema|erythema
Finding|Idea or Concept|SIMPLE_SEGMENT|580,590|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|580,595|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|596,606|false|false|false|C0007642|Cellulitis|cellulitis
Finding|Finding|SIMPLE_SEGMENT|596,606|false|false|false|C2025995|cellulitis on exam (physical finding)|cellulitis
Finding|Finding|SIMPLE_SEGMENT|622,626|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|622,626|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|622,626|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|SIMPLE_SEGMENT|651,654|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|651,654|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|651,654|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Antibiotic|SIMPLE_SEGMENT|689,699|false|false|false|C0007716|cephalexin|cephalexin
Drug|Organic Chemical|SIMPLE_SEGMENT|689,699|false|false|false|C0007716|cephalexin|cephalexin
Finding|Conceptual Entity|SIMPLE_SEGMENT|706,717|false|false|false|C2986411|Improvement|improvement
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|721,729|false|false|false|C0041834|Erythema|erythema
Attribute|Clinical Attribute|SIMPLE_SEGMENT|734,738|false|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|734,738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|734,738|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|753,761|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|753,761|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Gene or Genome|SIMPLE_SEGMENT|804,807|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Finding|Finding|SIMPLE_SEGMENT|840,847|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|840,847|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|SIMPLE_SEGMENT|840,859|false|false|false|C0231807|Dyspnea on exertion|dyspnea on exertion
Finding|Organism Function|SIMPLE_SEGMENT|851,859|false|false|false|C0015264|Exertion|exertion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|870,875|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|870,875|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|894,898|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|894,898|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|894,898|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|913,916|false|false|false|C0041912|Upper Respiratory Infections|URI
Finding|Gene or Genome|SIMPLE_SEGMENT|913,916|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Intellectual Product|SIMPLE_SEGMENT|913,916|false|false|false|C1421895;C1548524;C3272713|URI1 gene;URI1 wt Allele;Uniform Resource Identifier|URI
Finding|Functional Concept|SIMPLE_SEGMENT|917,925|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|SIMPLE_SEGMENT|917,925|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Anatomy|Body Location or Region|SIMPLE_SEGMENT|943,946|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|943,946|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|943,946|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Body Substance|SIMPLE_SEGMENT|951,958|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|951,958|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|951,958|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|SIMPLE_SEGMENT|970,975|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|970,975|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|977,983|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|SIMPLE_SEGMENT|985,994|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|985,999|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|995,999|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|995,999|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|995,999|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1001,1006|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1011,1018|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1011,1018|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1011,1018|false|false|false|C0872388|Procedures on bladder|bladder
Finding|Functional Concept|SIMPLE_SEGMENT|1019,1026|false|false|false|C0392747|Changing|changes
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1046,1049|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1046,1049|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|1046,1049|false|false|false|C0162574|Glycation End Products, Advanced|age
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1062,1068|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Finding|SIMPLE_SEGMENT|1070,1079|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|SIMPLE_SEGMENT|1070,1079|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1070,1079|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|SIMPLE_SEGMENT|1070,1079|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|SIMPLE_SEGMENT|1070,1079|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1091,1097|false|false|false|C0944911||weight
Finding|Finding|SIMPLE_SEGMENT|1091,1097|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|SIMPLE_SEGMENT|1091,1097|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|SIMPLE_SEGMENT|1091,1097|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|SIMPLE_SEGMENT|1091,1102|true|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|SIMPLE_SEGMENT|1091,1102|true|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Finding|SIMPLE_SEGMENT|1098,1102|true|false|false|C5890125|Loss (adaptation)|loss
Finding|Body Substance|SIMPLE_SEGMENT|1144,1151|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1144,1151|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1144,1151|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|1144,1155|false|false|false|C0332310|Has patient|patient has
Finding|Conceptual Entity|SIMPLE_SEGMENT|1165,1172|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1165,1172|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1165,1172|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1165,1175|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1178,1183|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1178,1183|false|false|false|C0006111|Brain Diseases|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1178,1192|false|false|false|C0751003|Brain Aneurysm|brain aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|1184,1192|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Idea or Concept|SIMPLE_SEGMENT|1201,1210|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|SIMPLE_SEGMENT|1201,1210|false|false|false|C1555324|inpatient encounter|inpatient
Finding|Conceptual Entity|SIMPLE_SEGMENT|1263,1267|false|false|false|C0868928;C1706256|Case - situation;Clinical Study Case|case
Finding|Functional Concept|SIMPLE_SEGMENT|1263,1267|false|false|false|C0868928;C1706256|Case - situation;Clinical Study Case|case
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1268,1281|false|false|false|C0016018|Fibrinolytic Agents|thrombolytics
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1314,1321|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Functional Concept|SIMPLE_SEGMENT|1336,1344|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1336,1344|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1336,1344|false|false|false|C4706767|Transfer (immobility management)|transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1360,1367|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|SIMPLE_SEGMENT|1368,1373|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1368,1379|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|SIMPLE_SEGMENT|1368,1379|false|false|false|C0150404|Taking vital signs|vital signs
Finding|Finding|SIMPLE_SEGMENT|1374,1379|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1374,1379|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1410,1414|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1410,1414|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1454,1458|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1454,1458|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|echo
Finding|Finding|SIMPLE_SEGMENT|1478,1483|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1478,1483|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|1487,1492|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1487,1498|false|false|false|C0225808|Right side of heart|right heart
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1493,1498|false|false|false|C0018787;C4037974|Chest>Heart;Heart|heart
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1493,1498|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|heart
Finding|Sign or Symptom|SIMPLE_SEGMENT|1493,1498|false|false|false|C0795691|HEART PROBLEM|heart
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|1499,1505|false|false|false|C0080194|Muscle strain|strain
Finding|Idea or Concept|SIMPLE_SEGMENT|1499,1505|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Mental Process|SIMPLE_SEGMENT|1499,1505|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Physiologic Function|SIMPLE_SEGMENT|1499,1505|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1499,1505|false|false|false|C0442694;C1510453;C1548152;C2987481|Emotional Strain;Nature of Abnormal Testing - Strain;Straining (finding);strain symptom|strain
Finding|Body Substance|SIMPLE_SEGMENT|1507,1514|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|1507,1514|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|1507,1514|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1545,1552|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|1545,1552|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1545,1552|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Gene or Genome|SIMPLE_SEGMENT|1581,1584|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|SIMPLE_SEGMENT|1581,1584|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1598,1601|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|1598,1601|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Functional Concept|SIMPLE_SEGMENT|1613,1621|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Finding|Idea or Concept|SIMPLE_SEGMENT|1613,1621|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|Transfer
Procedure|Health Care Activity|SIMPLE_SEGMENT|1613,1621|false|false|false|C4706767|Transfer (immobility management)|Transfer
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1657,1662|false|false|false|C0028429||Nasal
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1657,1662|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Organic Chemical|SIMPLE_SEGMENT|1657,1662|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1657,1662|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|Nasal
Finding|Finding|SIMPLE_SEGMENT|1657,1662|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Finding|Functional Concept|SIMPLE_SEGMENT|1657,1662|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|Nasal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1663,1670|false|false|false|C1550232|Body Parts - Cannula|Cannula
Finding|Body Substance|SIMPLE_SEGMENT|1663,1670|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Finding|Intellectual Product|SIMPLE_SEGMENT|1663,1670|false|false|false|C1546577;C1550622|Specimen Type - Cannula|Cannula
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1677,1686|false|false|false|C5885990||breathing
Finding|Finding|SIMPLE_SEGMENT|1677,1686|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|SIMPLE_SEGMENT|1677,1686|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|SIMPLE_SEGMENT|1677,1686|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|SIMPLE_SEGMENT|1677,1686|false|false|false|C1160636|respiratory system process|breathing
Finding|Finding|SIMPLE_SEGMENT|1690,1697|false|false|false|C3840786|Greatly|greatly
Finding|Finding|SIMPLE_SEGMENT|1698,1706|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|SIMPLE_SEGMENT|1698,1706|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1723,1728|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1723,1728|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1723,1733|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1723,1733|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1729,1733|true|false|false|C2598155||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1729,1733|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1729,1733|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|SIMPLE_SEGMENT|1740,1760|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Finding|Functional Concept|SIMPLE_SEGMENT|1745,1752|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1745,1752|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1745,1752|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1745,1752|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1745,1760|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1753,1760|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1753,1760|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1753,1760|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1762,1770|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|CEREBRAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1762,1779|false|false|false|C0917996|Cerebral Aneurysm|CEREBRAL ANEURYSM
Finding|Pathologic Function|SIMPLE_SEGMENT|1771,1779|false|false|false|C0002940|Aneurysm|ANEURYSM
Finding|Functional Concept|SIMPLE_SEGMENT|1782,1792|false|false|false|C0444507|Incidental|incidental
Finding|Finding|SIMPLE_SEGMENT|1782,1800|false|false|false|C0743997|Incidental Findings|incidental finding
Finding|Finding|SIMPLE_SEGMENT|1793,1800|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|SIMPLE_SEGMENT|1793,1800|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Finding|SIMPLE_SEGMENT|1848,1854|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|1848,1854|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Sign or Symptom|SIMPLE_SEGMENT|1859,1868|false|false|false|C0012833;C0042571|Dizziness;Vertigo|dizziness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1870,1874|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1870,1874|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1870,1874|false|false|false|C0362076|Problems with head|Head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1870,1874|false|false|false|C0876917|Procedure on head|Head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1870,1877|false|false|false|C0202691|CAT scan of head|Head CT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1898,1914|false|false|false|C0333559|Infarction, Lacunar|lacunar infarcts
Finding|Pathologic Function|SIMPLE_SEGMENT|1906,1914|false|false|false|C0021308|Infarction|infarcts
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1923,1936|false|false|false|C0004781;C1321510|Basal Ganglia|basal ganglia
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1929,1936|false|false|false|C0017067|Ganglia|ganglia
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|1971,1979|true|false|false|C0009924|Contrast Media|contrast
Finding|Intellectual Product|SIMPLE_SEGMENT|1983,1989|false|false|false|C1547311|Patient Condition Code - Stable|stable
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1995,2007|false|false|false|C2339173|Protuberance|protuberance
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2016,2020|false|false|false|C0022742;C0152321|Knee;Structure of genu of corpus callosum|genu
Finding|Functional Concept|SIMPLE_SEGMENT|2028,2032|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2044,2051|false|false|false|C0007272|Carotid Arteries|carotid
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2044,2058|false|false|false|C0007272;C0162859;C1305384;C4071877|Carotid Arteries;Common carotid artery;Head+Neck>Carotid artery|carotid artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2052,2058|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|2052,2058|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2092,2095|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|2092,2095|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2092,2095|false|false|false|C1609165|tocilizumab|MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2092,2095|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2092,2095|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2119,2124|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2119,2124|false|false|false|C1528558|BRCA1 protein, human|BRCA1
Finding|Gene or Genome|SIMPLE_SEGMENT|2119,2124|false|false|false|C0376571|BRCA1 gene|BRCA1
Finding|Gene or Genome|SIMPLE_SEGMENT|2119,2129|false|false|false|C0376571|BRCA1 gene|BRCA1 GENE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|2119,2129|false|false|false|C2010863|BRCA1 gene (lab test)|BRCA1 GENE
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2119,2138|false|false|false|C1511022|BRCA1 gene mutation|BRCA1 GENE MUTATION
Finding|Finding|SIMPLE_SEGMENT|2125,2129|false|false|false|C0017337;C5849123|Genes;Gross Extranodal Extension|GENE
Finding|Gene or Genome|SIMPLE_SEGMENT|2125,2129|false|false|false|C0017337;C5849123|Genes;Gross Extranodal Extension|GENE
Finding|Gene or Genome|SIMPLE_SEGMENT|2125,2138|false|false|false|C0596611;C0678941|Gene Mutant;Gene Mutation|GENE MUTATION
Finding|Genetic Function|SIMPLE_SEGMENT|2125,2138|false|false|false|C0596611;C0678941|Gene Mutant;Gene Mutation|GENE MUTATION
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|2130,2138|false|false|false|C1705285|Mutation Abnormality|MUTATION
Finding|Genetic Function|SIMPLE_SEGMENT|2130,2138|false|false|false|C0026882|Mutation|MUTATION
Finding|Intellectual Product|SIMPLE_SEGMENT|2141,2148|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|SIMPLE_SEGMENT|2141,2148|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2141,2178|false|false|false|C0024117|Chronic Obstructive Airway Disease|CHRONIC OBSTRUCTIVE PULMONARY DISEASE
Finding|Functional Concept|SIMPLE_SEGMENT|2149,2160|false|false|false|C0549186|Obstructed|OBSTRUCTIVE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2149,2178|false|false|false|C0600260|Lung Diseases, Obstructive|OBSTRUCTIVE PULMONARY DISEASE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2161,2170|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2161,2170|false|false|false|C2707265||PULMONARY
Finding|Finding|SIMPLE_SEGMENT|2161,2170|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2161,2178|false|false|false|C0024115|Lung diseases|PULMONARY DISEASE
Finding|Finding|SIMPLE_SEGMENT|2161,2178|false|false|false|C0455540|History of - respiratory disease|PULMONARY DISEASE
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2171,2178|false|true|false|C0012634|Disease|DISEASE
Drug|Organic Chemical|SIMPLE_SEGMENT|2181,2186|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|SLEEP
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2181,2186|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|SLEEP
Finding|Organism Function|SIMPLE_SEGMENT|2181,2186|false|false|false|C0037313|Sleep|SLEEP
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2181,2192|false|false|false|C0037315|Sleep Apnea Syndromes|SLEEP APNEA
Finding|Sign or Symptom|SIMPLE_SEGMENT|2187,2192|false|false|false|C0003578|Apnea|APNEA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2195,2202|false|false|false|C0009368|Colon structure (body structure)|COLONIC
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2195,2209|false|false|false|C0009376|Colonic Polyps|COLONIC POLYPS
Finding|Finding|SIMPLE_SEGMENT|2195,2209|false|false|false|C2911243|Encounter due to family history of colonic polyps|COLONIC POLYPS
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2203,2209|false|false|false|C0032584|polyps|POLYPS
Finding|Intellectual Product|SIMPLE_SEGMENT|2203,2209|false|false|false|C1546747||POLYPS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2212,2228|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2212,2235|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|SIMPLE_SEGMENT|2212,2235|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Finding|Pathologic Function|SIMPLE_SEGMENT|2229,2235|false|false|false|C0232483|Reflux|REFLUX
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|2238,2248|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|DEPRESSION
Finding|Functional Concept|SIMPLE_SEGMENT|2238,2248|false|false|false|C0460137;C1579931|Depression - motion|DEPRESSION
Finding|Sign or Symptom|SIMPLE_SEGMENT|2238,2248|false|false|false|C0460137;C1579931|Depression - motion|DEPRESSION
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2251,2263|false|false|false|C0362046|Prediabetes syndrome|PRE-DIABETES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2269,2278|false|false|false|C0018965|Hematuria|HEMATURIA
Finding|Finding|SIMPLE_SEGMENT|2281,2284|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|LOW
Finding|Intellectual Product|SIMPLE_SEGMENT|2281,2284|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|LOW
Finding|Sign or Symptom|SIMPLE_SEGMENT|2281,2294|false|true|false|C0024031|Low Back Pain|LOW BACK PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|2285,2294|false|true|false|C0004604|Back Pain|BACK PAIN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2290,2294|false|false|false|C2598155||PAIN
Finding|Functional Concept|SIMPLE_SEGMENT|2290,2294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|SIMPLE_SEGMENT|2290,2294|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2295,2309|false|false|false|C0042345|Varicosity|VARICOSE VEINS
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2304,2309|false|false|false|C0042449|Veins|VEINS
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2304,2309|false|false|false|C0398102|Procedure on vein|VEINS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2316,2323|false|false|false|C0036262|Scabies infestation|SCABIES
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2326,2340|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Finding|Finding|SIMPLE_SEGMENT|2326,2340|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2343,2355|false|false|false|C0085515|Rotator Cuff|ROTATOR CUFF
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2343,2360|false|false|false|C0263912|Rotator cuff syndrome|ROTATOR CUFF TEAR
Finding|Finding|SIMPLE_SEGMENT|2343,2360|false|false|false|C5399759|Rotator Cuff Tears|ROTATOR CUFF TEAR
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2351,2355|false|false|false|C1550244|Cuff - body part|CUFF
Finding|Pathologic Function|SIMPLE_SEGMENT|2351,2355|false|false|false|C3668885|Cuffing (morphologic abnormality)|CUFF
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|2356,2360|false|false|false|C0043246;C3203359|Laceration;Rupture|TEAR
Finding|Body Substance|SIMPLE_SEGMENT|2356,2360|false|false|false|C0039409|Tears (substance)|TEAR
Finding|Sign or Symptom|SIMPLE_SEGMENT|2363,2370|false|false|false|C0039070|Syncope|syncope
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2374,2377|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2378,2385|false|false|false|C0007272|Carotid Arteries|carotid
Finding|Idea or Concept|SIMPLE_SEGMENT|2412,2423|true|false|false|C0750502|Significant|significant
Finding|Pathologic Function|SIMPLE_SEGMENT|2427,2435|false|false|false|C1261287|Stenosis|stenosis
Procedure|Health Care Activity|SIMPLE_SEGMENT|2437,2441|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2437,2441|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2448,2451|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2448,2455|false|false|false|C0542407|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|TAH/BSO
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|2452,2455|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|2452,2455|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2452,2455|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|2458,2473|false|false|false|C0008320|Cholecystectomy procedure|CHOLECYSTECTOMY
Finding|Functional Concept|SIMPLE_SEGMENT|2479,2485|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|2479,2493|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2486,2493|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2486,2493|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2486,2493|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|2499,2505|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|2499,2513|false|false|false|C0241889|Family Medical History|Family History
Finding|Conceptual Entity|SIMPLE_SEGMENT|2506,2513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|2506,2513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|2506,2513|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|2518,2524|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|SIMPLE_SEGMENT|2518,2524|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|SIMPLE_SEGMENT|2518,2524|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|SIMPLE_SEGMENT|2518,2524|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2531,2534|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2531,2534|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2531,2534|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2559,2565|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2559,2578|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2559,2578|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|2559,2578|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2566,2578|false|false|false|C0232197|Fibrillation|fibrillation
Finding|Finding|SIMPLE_SEGMENT|2585,2593|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|2585,2593|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|2585,2593|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|2585,2598|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2585,2598|false|false|false|C0031809|Physical Examination|Physical Exam
Finding|Functional Concept|SIMPLE_SEGMENT|2594,2598|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2594,2598|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|2603,2612|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Classification|SIMPLE_SEGMENT|2647,2654|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2647,2654|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2656,2659|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2656,2659|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2656,2659|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2656,2659|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2656,2659|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|2656,2659|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2661,2666|false|false|false|C0028754|Obesity|obese
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2669,2674|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|2689,2694|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|SIMPLE_SEGMENT|2696,2705|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2706,2712|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2706,2712|false|false|false|C0036412|Scleral Diseases|sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2706,2712|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2719,2730|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2719,2730|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2719,2730|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|2719,2730|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|2719,2730|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|2719,2730|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2733,2736|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2733,2736|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Idea or Concept|SIMPLE_SEGMENT|2738,2742|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2743,2752|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2755,2759|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|2755,2759|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|2755,2759|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|SIMPLE_SEGMENT|2771,2777|false|false|false|C0332254|Supple|supple
Finding|Finding|SIMPLE_SEGMENT|2771,2782|false|false|false|C2230237|Supple neck|supple neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2778,2782|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2778,2782|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|2778,2782|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2787,2790|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2787,2790|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|2787,2790|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|2795,2798|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2801,2808|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|2801,2808|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|2825,2832|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|2846,2850|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2853,2857|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2853,2857|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2853,2857|false|false|false|C0024115|Lung diseases|LUNG
Finding|Finding|SIMPLE_SEGMENT|2853,2857|false|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|SIMPLE_SEGMENT|2859,2863|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Sign or Symptom|SIMPLE_SEGMENT|2868,2875|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|SIMPLE_SEGMENT|2877,2882|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|SIMPLE_SEGMENT|2884,2891|true|false|false|C0035508|Rhonchi|rhonchi
Finding|Functional Concept|SIMPLE_SEGMENT|2924,2927|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|2924,2927|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|SIMPLE_SEGMENT|2924,2930|true|false|false|C1524063|Use of|use of
Finding|Finding|SIMPLE_SEGMENT|2924,2948|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2931,2948|false|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2941,2948|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|2941,2948|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2951,2958|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2951,2958|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|2951,2958|false|false|false|C0941288|Abdomen problem|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3019,3027|false|false|false|C0427198|Protective muscle spasm|guarding
Finding|Sign or Symptom|SIMPLE_SEGMENT|3032,3050|true|false|false|C0019214|Hepatosplenomegaly|hepatosplenomegaly
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3053,3064|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3081,3086|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3081,3086|false|false|false|C2003888|Lower (action)|lower
Finding|Functional Concept|SIMPLE_SEGMENT|3087,3091|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3087,3091|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|SIMPLE_SEGMENT|3092,3100|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|3092,3100|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3110,3116|false|false|false|C0489801|Posterior part of right leg|R calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3112,3116|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3112,3116|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3131,3140|false|false|false|C0030247|Palpation|palpation
Drug|Food|SIMPLE_SEGMENT|3141,3147|false|false|false|C5890763||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3141,3147|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3141,3147|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|SIMPLE_SEGMENT|3155,3161|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3155,3161|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3155,3161|false|false|false|C0034107|Pulse taking|pulses
Finding|Finding|SIMPLE_SEGMENT|3193,3199|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body System|SIMPLE_SEGMENT|3221,3225|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3221,3225|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3221,3225|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3221,3225|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3221,3225|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Finding|SIMPLE_SEGMENT|3227,3231|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3227,3231|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3236,3240|false|false|false|C5575035|Well (answer to question)|well
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3254,3266|true|false|false|C0015256|Excoriation|excoriations
Finding|Finding|SIMPLE_SEGMENT|3270,3277|true|false|false|C0221198|Lesion|lesions
Finding|Sign or Symptom|SIMPLE_SEGMENT|3283,3289|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Body Substance|SIMPLE_SEGMENT|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3297,3306|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3297,3306|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Classification|SIMPLE_SEGMENT|3340,3347|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|3340,3347|false|false|false|C3812897|General medical service|GENERAL
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3349,3352|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3349,3352|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3349,3352|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|3349,3352|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3349,3352|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|SIMPLE_SEGMENT|3349,3352|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3354,3359|false|false|false|C0028754|Obesity|obese
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3362,3367|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|SIMPLE_SEGMENT|3382,3387|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Finding|Finding|SIMPLE_SEGMENT|3389,3398|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3399,3405|false|false|false|C0036410|Sclera|sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3399,3405|false|false|false|C0036412|Scleral Diseases|sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|3399,3405|false|false|false|C2228481|examination of sclera|sclera
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3412,3423|false|false|false|C0009758;C0229274|Structure of palpebral conjunctiva;conjunctiva|conjunctiva
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3412,3423|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3412,3423|false|false|false|C0009759;C0153628;C0154025|Benign neoplasm of conjunctiva;Conjunctival Diseases;Malignant neoplasm of conjunctiva|conjunctiva
Finding|Body Substance|SIMPLE_SEGMENT|3412,3423|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Finding|Intellectual Product|SIMPLE_SEGMENT|3412,3423|false|false|false|C1546576;C1550624|Specimen Type - Conjunctiva|conjunctiva
Procedure|Health Care Activity|SIMPLE_SEGMENT|3412,3423|false|false|false|C0872390;C2228431|Procedure on conjunctiva;examination of conjunctiva|conjunctiva
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3426,3429|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3426,3429|false|false|false|C0026987|Myelofibrosis|MMM
Finding|Idea or Concept|SIMPLE_SEGMENT|3431,3435|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3436,3445|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3448,3452|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|SIMPLE_SEGMENT|3448,3452|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|SIMPLE_SEGMENT|3448,3452|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Finding|Functional Concept|SIMPLE_SEGMENT|3464,3470|false|false|false|C0332254|Supple|supple
Finding|Finding|SIMPLE_SEGMENT|3464,3475|false|false|false|C2230237|Supple neck|supple neck
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3471,3475|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|SIMPLE_SEGMENT|3471,3475|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|SIMPLE_SEGMENT|3471,3475|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3480,3483|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3480,3483|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Finding|Gene or Genome|SIMPLE_SEGMENT|3480,3483|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Finding|Finding|SIMPLE_SEGMENT|3488,3491|true|false|false|C0425687|Jugular venous engorgement|JVD
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3494,3501|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|SIMPLE_SEGMENT|3494,3501|false|false|false|C1314974|Cardiac attachment|CARDIAC
Finding|Finding|SIMPLE_SEGMENT|3518,3525|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|SIMPLE_SEGMENT|3539,3543|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3546,3550|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3546,3550|false|false|false|C0024109;C4037972|Chest>Lung;Lung|LUNG
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3546,3550|false|false|false|C0024115|Lung diseases|LUNG
Finding|Finding|SIMPLE_SEGMENT|3546,3550|false|false|false|C0740941|Lung Problem|LUNG
Drug|Organic Chemical|SIMPLE_SEGMENT|3552,3556|false|false|false|C0951233|cetrimonium bromide|CTAB
Finding|Sign or Symptom|SIMPLE_SEGMENT|3561,3568|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|SIMPLE_SEGMENT|3570,3575|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|SIMPLE_SEGMENT|3577,3584|true|false|false|C0035508|Rhonchi|rhonchi
Finding|Functional Concept|SIMPLE_SEGMENT|3617,3620|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|SIMPLE_SEGMENT|3617,3620|true|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Functional Concept|SIMPLE_SEGMENT|3617,3623|true|false|false|C1524063|Use of|use of
Finding|Finding|SIMPLE_SEGMENT|3617,3641|true|false|false|C1821466|Use of accessory muscles|use of accessory muscles
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3624,3641|false|false|false|C0158784|Accessory skeletal muscle|accessory muscles
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3634,3641|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Tissue|SIMPLE_SEGMENT|3634,3641|false|false|false|C0026845;C1995013;C4083049|Muscle (organ);Muscle Tissue;Set of muscles|muscles
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3644,3651|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3644,3651|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3644,3651|false|false|false|C0941288|Abdomen problem|ABDOMEN
Finding|Finding|SIMPLE_SEGMENT|3712,3720|false|false|false|C0427198|Protective muscle spasm|guarding
Finding|Sign or Symptom|SIMPLE_SEGMENT|3725,3743|true|false|false|C0019214|Hepatosplenomegaly|hepatosplenomegaly
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3746,3757|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3774,3779|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3774,3779|false|false|false|C2003888|Lower (action)|lower
Finding|Functional Concept|SIMPLE_SEGMENT|3780,3784|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|3780,3784|false|false|false|C0582103|Medical Examination|exam
Finding|Finding|SIMPLE_SEGMENT|3785,3793|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|3785,3793|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3803,3809|false|false|false|C0489801|Posterior part of right leg|R calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3805,3809|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3805,3809|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3824,3833|false|false|false|C0030247|Palpation|palpation
Drug|Food|SIMPLE_SEGMENT|3834,3840|false|false|false|C5890763||PULSES
Finding|Physiologic Function|SIMPLE_SEGMENT|3834,3840|false|false|false|C0391850|Physiologic pulse|PULSES
Procedure|Health Care Activity|SIMPLE_SEGMENT|3834,3840|false|false|false|C0034107|Pulse taking|PULSES
Drug|Food|SIMPLE_SEGMENT|3848,3854|false|false|false|C5890763||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3848,3854|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3848,3854|false|false|false|C0034107|Pulse taking|pulses
Finding|Finding|SIMPLE_SEGMENT|3886,3892|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body System|SIMPLE_SEGMENT|3914,3918|false|false|false|C1123023;C4520765|Skin;Skin, Human|SKIN
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3914,3918|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3914,3918|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|SKIN
Finding|Body Substance|SIMPLE_SEGMENT|3914,3918|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Intellectual Product|SIMPLE_SEGMENT|3914,3918|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|SKIN
Finding|Finding|SIMPLE_SEGMENT|3920,3924|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3920,3924|false|false|false|C0687712|warming process|warm
Finding|Finding|SIMPLE_SEGMENT|3929,3933|false|false|false|C5575035|Well (answer to question)|well
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|3947,3959|true|false|false|C0015256|Excoriation|excoriations
Finding|Finding|SIMPLE_SEGMENT|3963,3970|true|false|false|C0221198|Lesion|lesions
Finding|Sign or Symptom|SIMPLE_SEGMENT|3976,3982|false|false|false|C0015230;C5779628|Exanthema;Skin rash|rashes
Finding|Body Substance|SIMPLE_SEGMENT|3987,3996|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|3987,3996|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|3987,3996|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|3987,3996|false|false|false|C0030685|Patient Discharge|DISCHARGE
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4037,4040|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4037,4040|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4066,4069|false|false|false|C0201617|Primed lymphocyte test|PLT
Drug|Antibiotic|SIMPLE_SEGMENT|4109,4114|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|4109,4114|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Drug|Organic Chemical|SIMPLE_SEGMENT|4109,4114|false|false|false|C0540173;C3275179|Mono-S;Monos|MONOS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4119,4122|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|EOS
Finding|Gene or Genome|SIMPLE_SEGMENT|4119,4122|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|EOS
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4152,4159|false|false|false|C0017725|glucose|GLUCOSE
Drug|Organic Chemical|SIMPLE_SEGMENT|4152,4159|false|false|false|C0017725|glucose|GLUCOSE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4152,4159|false|false|false|C0017725|glucose|GLUCOSE
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4152,4159|false|false|false|C5781949|Glucose^1.5H post dose glucagon|GLUCOSE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4152,4159|false|false|false|C0337438|Glucose measurement|GLUCOSE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4165,4169|false|false|false|C0041942|urea|UREA
Drug|Organic Chemical|SIMPLE_SEGMENT|4165,4169|false|false|false|C0041942|urea|UREA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4165,4169|false|false|false|C0041942|urea|UREA
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4165,4169|false|false|false|C0523961|Urea measurement|UREA
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4185,4191|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4185,4191|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4185,4191|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|SODIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4185,4191|false|false|false|C4553025|Sodium metabolic function|SODIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4185,4191|false|false|false|C0337443|Sodium measurement|SODIUM
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4197,4206|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4197,4206|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Food|SIMPLE_SEGMENT|4197,4206|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4197,4206|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4197,4206|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|POTASSIUM
Finding|Physiologic Function|SIMPLE_SEGMENT|4197,4206|false|false|false|C4553027|Potassium metabolic function|POTASSIUM
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4197,4206|false|false|false|C0202194|Potassium measurement|POTASSIUM
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4211,4219|false|false|false|C0008203;C0596019|Chlorides;chloride ion|CHLORIDE
Finding|Physiologic Function|SIMPLE_SEGMENT|4211,4219|false|false|false|C4553021|Chloride metabolic function|CHLORIDE
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4211,4219|false|false|false|C0201952|Chloride measurement|CHLORIDE
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4230,4233|false|false|false|C0007012|carbon dioxide|CO2
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4230,4233|false|false|false|C0007012|carbon dioxide|CO2
Finding|Finding|SIMPLE_SEGMENT|4230,4233|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Finding|Gene or Genome|SIMPLE_SEGMENT|4230,4233|false|false|false|C0860710;C1537986;C4284286|C2 wt Allele;MT-CO2 gene|CO2
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4237,4242|false|false|false|C0003075|Anions|ANION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4237,4246|false|false|false|C0003074|Anion Gap|ANION GAP
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4237,4246|false|false|false|C1509129|Anion gap result|ANION GAP
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4237,4246|false|false|false|C0201889;C2189246|Anion gap measurement;blood anion gap (lab test)|ANION GAP
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4243,4246|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4243,4246|false|false|false|C0061928;C2984553|GTPase-Activating Proteins;Ras GTPase-Activating Protein 1, Human|GAP
Finding|Gene or Genome|SIMPLE_SEGMENT|4243,4246|false|false|false|C1419277;C2984552|RASA1 gene;RASA1 wt Allele|GAP
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4268,4271|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4268,4271|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Finding|Conceptual Entity|SIMPLE_SEGMENT|4283,4290|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4283,4290|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|4283,4290|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|4283,4293|false|false|false|C0262926|Medical History|history of
Finding|Finding|SIMPLE_SEGMENT|4283,4311|false|false|false|C5192533|History of cerebral aneurysm|history of cerebral aneurysm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4294,4302|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4294,4311|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|4303,4311|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Conceptual Entity|SIMPLE_SEGMENT|4320,4329|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|4320,4329|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|4320,4329|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4320,4329|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Finding|SIMPLE_SEGMENT|4339,4347|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|4339,4347|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4352,4360|false|false|false|C0041834|Erythema|erythema
Drug|Antibiotic|SIMPLE_SEGMENT|4366,4372|false|false|false|C0700517|Keflex|keflex
Drug|Organic Chemical|SIMPLE_SEGMENT|4366,4372|false|false|false|C0700517|Keflex|keflex
Finding|Classification|SIMPLE_SEGMENT|4386,4394|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|4386,4394|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4386,4394|false|false|false|C5237010|Expression Negative|negative
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4424,4443|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|4424,4443|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|4437,4443|false|false|false|C0225386|Breath|breath
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4467,4476|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4467,4476|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|4467,4476|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|4467,4485|false|false|false|C0034065|Pulmonary Embolism|Pulmonary embolism
Finding|Finding|SIMPLE_SEGMENT|4477,4485|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|4477,4485|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Drug|Organic Chemical|SIMPLE_SEGMENT|4499,4506|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4499,4506|false|false|false|C0728963|Lovenox|lovenox
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|4544,4552|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|4544,4552|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4544,4552|false|false|false|C0043031|warfarin|warfarin
Finding|Body Substance|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|4556,4565|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|4556,4565|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4567,4586|false|false|false|C2707305||Shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|4567,4586|false|false|false|C0013404|Dyspnea|Shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|4580,4586|false|false|false|C0225386|Breath|breath
Finding|Functional Concept|SIMPLE_SEGMENT|4628,4632|true|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|SIMPLE_SEGMENT|4628,4636|true|false|false|C0686904|Patient need for (contextual qualifier)|need for
Finding|Functional Concept|SIMPLE_SEGMENT|4637,4649|false|false|false|C2348609|Supplement|supplemental
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4651,4657|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|4651,4657|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4651,4657|false|false|false|C0030054|oxygen|oxygen
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4651,4657|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Finding|Conceptual Entity|SIMPLE_SEGMENT|4662,4669|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|4662,4669|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|4662,4669|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|4662,4672|false|false|false|C0262926|Medical History|History of
Finding|Finding|SIMPLE_SEGMENT|4662,4690|false|false|false|C5192533|History of cerebral aneurysm|History of cerebral aneurysm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4673,4681|false|false|false|C0006104;C0228174|Brain;Cerebral hemisphere structure (body structure)|cerebral
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4673,4690|false|false|false|C0917996|Cerebral Aneurysm|cerebral aneurysm
Finding|Pathologic Function|SIMPLE_SEGMENT|4682,4690|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Body Substance|SIMPLE_SEGMENT|4720,4727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|4720,4727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|4720,4727|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Pathologic Function|SIMPLE_SEGMENT|4730,4738|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Functional Concept|SIMPLE_SEGMENT|4764,4770|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|SIMPLE_SEGMENT|4764,4770|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Gene or Genome|SIMPLE_SEGMENT|4775,4778|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4775,4778|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|4775,4778|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Finding|Pathologic Function|SIMPLE_SEGMENT|4819,4827|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Finding|SIMPLE_SEGMENT|4838,4851|false|false|false|C0518609|Consideration|consideration
Drug|Organic Chemical|SIMPLE_SEGMENT|4880,4887|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4880,4887|false|false|false|C0004057|aspirin|aspirin
Finding|Pathologic Function|SIMPLE_SEGMENT|4913,4921|false|false|false|C0002940|Aneurysm|aneurysm
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4939,4953|false|false|false|C3536711|Anti-coagulant [EPC]|anti-coagulant
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4967,4972|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4967,4972|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|SIMPLE_SEGMENT|4967,4972|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|SIMPLE_SEGMENT|4967,4972|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|SIMPLE_SEGMENT|4967,4972|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|4967,4972|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4967,4972|false|false|false|C0031765|Phototherapy|light
Finding|Pathologic Function|SIMPLE_SEGMENT|4980,4988|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Idea or Concept|SIMPLE_SEGMENT|5005,5009|false|false|false|C0035647|Risk|risk
Finding|Idea or Concept|SIMPLE_SEGMENT|5005,5012|false|false|false|C0035647|Risk|risk of
Finding|Pathologic Function|SIMPLE_SEGMENT|5014,5022|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Social Behavior|SIMPLE_SEGMENT|5030,5040|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5030,5040|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Mental Process|SIMPLE_SEGMENT|5063,5071|false|false|false|C0679006|Decision|decision
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5084,5090|false|false|false|C0399080|Fixation of dental bridge|bridge
Drug|Organic Chemical|SIMPLE_SEGMENT|5094,5102|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5094,5102|false|false|false|C0699129|Coumadin|Coumadin
Drug|Organic Chemical|SIMPLE_SEGMENT|5108,5115|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5108,5115|false|false|false|C0728963|Lovenox|lovenox
Event|Activity|SIMPLE_SEGMENT|5120,5124|false|false|false|C1948035|Hold (action)|hold
Finding|Functional Concept|SIMPLE_SEGMENT|5120,5124|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Finding|Intellectual Product|SIMPLE_SEGMENT|5120,5124|false|false|false|C1553387;C3853841|Hold - dosing instruction fragment;hold - Data Operation|hold
Drug|Organic Chemical|SIMPLE_SEGMENT|5130,5137|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5130,5137|false|false|false|C0004057|aspirin|aspirin
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5143,5146|false|false|false|C1609165|tocilizumab|MRA
Drug|Immunologic Factor|SIMPLE_SEGMENT|5143,5146|false|false|false|C1609165|tocilizumab|MRA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5143,5146|false|false|false|C1609165|tocilizumab|MRA
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5143,5146|false|false|false|C3891069|MRI-Based Angiogram|MRA
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5143,5146|false|false|false|C0243032|Magnetic Resonance Angiography|MRA
Finding|Pathologic Function|SIMPLE_SEGMENT|5194,5202|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Body Substance|SIMPLE_SEGMENT|5213,5220|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5213,5220|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5213,5220|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5241,5247|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Pathologic Function|SIMPLE_SEGMENT|5261,5269|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Functional Concept|SIMPLE_SEGMENT|5284,5290|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5284,5290|true|false|false|C4319952|Change - procedure|change
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5304,5318|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Finding|Finding|SIMPLE_SEGMENT|5304,5318|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Organic Chemical|SIMPLE_SEGMENT|5330,5342|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5330,5342|false|false|false|C0286651|atorvastatin|atorvastatin
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5350,5360|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|Depression
Finding|Functional Concept|SIMPLE_SEGMENT|5350,5360|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Sign or Symptom|SIMPLE_SEGMENT|5350,5360|false|false|false|C0460137;C1579931|Depression - motion|Depression
Finding|Idea or Concept|SIMPLE_SEGMENT|5372,5376|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5372,5376|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5372,5376|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5391,5395|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Finding|Idea or Concept|SIMPLE_SEGMENT|5407,5411|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|5407,5411|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|5407,5411|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|SIMPLE_SEGMENT|5412,5422|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5412,5422|false|false|false|C0028978|omeprazole|omeprazole
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5427,5433|false|false|false|C0004096|Asthma|Asthma
Finding|Idea or Concept|SIMPLE_SEGMENT|5438,5446|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5438,5449|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5450,5458|false|false|false|C4722408|Reactive Therapy|reactive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5450,5473|true|false|false|C3714496;C3714497|Chronic obstructive pulmonary disease of horses;Reactive airway disease|reactive airway disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5459,5465|false|false|false|C0458827;C4071894|Airway structure;Chest>Airway|airway
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5459,5473|true|false|false|C0699949|airway disease|airway disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5466,5473|true|false|false|C0012634|Disease|disease
Finding|Functional Concept|SIMPLE_SEGMENT|5477,5481|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|5477,5481|false|false|false|C0582103|Medical Examination|exam
Drug|Organic Chemical|SIMPLE_SEGMENT|5494,5503|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5494,5503|false|false|false|C0001927|albuterol|albuterol
Finding|Functional Concept|SIMPLE_SEGMENT|5504,5511|false|false|false|C4319647|Inhaler (unit of presentation)|inhaler
Finding|Idea or Concept|SIMPLE_SEGMENT|5526,5538|false|false|false|C1548597|Marketing basis - Transitional|Transitional
Finding|Physiologic Function|SIMPLE_SEGMENT|5549,5565|false|false|false|C3537050|Decreased Coagulation Activity [PE]|Anti-coagulation
Finding|Intellectual Product|SIMPLE_SEGMENT|5581,5588|false|false|false|C3260738|Outpatient Physical Therapy Improvement in Movement and Assessment Log (OPTIMAL) Survey|optimal
Finding|Conceptual Entity|SIMPLE_SEGMENT|5599,5608|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|SIMPLE_SEGMENT|5599,5608|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|SIMPLE_SEGMENT|5599,5608|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5599,5608|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Body Substance|SIMPLE_SEGMENT|5618,5625|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5618,5625|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5618,5625|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5630,5639|false|false|false|C1704760|Cigarette Dosage Form|Cigarette
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|5630,5647|false|false|false|C0239059|Cigarette smoke (substance)|Cigarette smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|5630,5647|false|false|false|C0700219|Cigarette smoking behavior|Cigarette smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|5640,5647|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|5640,5647|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Body Substance|SIMPLE_SEGMENT|5653,5660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|5653,5660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|5653,5660|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Procedure|Health Care Activity|SIMPLE_SEGMENT|5677,5686|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Social Behavior|SIMPLE_SEGMENT|5718,5731|false|false|false|C0870494|encouragement|encouragement
Finding|Idea or Concept|SIMPLE_SEGMENT|5736,5745|false|false|false|C0035201|Resources|resources
Finding|Individual Behavior|SIMPLE_SEGMENT|5757,5764|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Intellectual Product|SIMPLE_SEGMENT|5757,5764|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|smoking
Finding|Individual Behavior|SIMPLE_SEGMENT|5757,5774|false|false|false|C0085134|Cessation of smoking|smoking cessation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5757,5774|false|false|false|C1095963|Smoking cessation therapy|smoking cessation
Event|Activity|SIMPLE_SEGMENT|5765,5774|false|false|false|C1880019|Cessation|cessation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5779,5790|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5779,5790|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|5779,5790|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|5779,5803|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|5794,5803|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5822,5832|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5822,5832|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|5822,5837|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|SIMPLE_SEGMENT|5833,5837|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|SIMPLE_SEGMENT|5854,5862|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5854,5862|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|5854,5862|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|SIMPLE_SEGMENT|5854,5862|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|5854,5862|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|SIMPLE_SEGMENT|5867,5877|false|false|false|C0024027|lovastatin|Lovastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5867,5877|false|false|false|C0024027|lovastatin|Lovastatin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5884,5888|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|5884,5888|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|5884,5888|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|5884,5888|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|5899,5909|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5899,5909|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|5930,5937|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5930,5937|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|5958,5968|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5958,5968|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|5978,5981|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5978,5981|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5978,5981|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|5978,5981|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|5986,5995|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5986,5995|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|5986,6003|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5986,6003|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5996,6003|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5996,6003|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5996,6003|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|6021,6031|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|6021,6031|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|SIMPLE_SEGMENT|6038,6041|false|false|false|C1422467|CIAO3 gene|prn
Finding|Sign or Symptom|SIMPLE_SEGMENT|6043,6051|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|SIMPLE_SEGMENT|6056,6063|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6056,6063|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|6056,6063|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|6056,6065|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|6056,6065|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6056,6065|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|6056,6065|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6056,6065|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|6088,6101|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6088,6101|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|6088,6101|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6104,6112|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6115,6118|false|false|false|C0039225|Tablet Dosage Form|TAB
Finding|Body Substance|SIMPLE_SEGMENT|6132,6141|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6132,6141|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6132,6141|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6132,6141|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6132,6153|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6142,6153|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6142,6153|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|6142,6153|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|6158,6168|false|false|false|C0024027|lovastatin|Lovastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6158,6168|false|false|false|C0024027|lovastatin|Lovastatin
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6175,6179|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6175,6179|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|SIMPLE_SEGMENT|6175,6179|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|SIMPLE_SEGMENT|6175,6179|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Organic Chemical|SIMPLE_SEGMENT|6190,6203|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6190,6203|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|6190,6203|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6206,6214|false|false|false|C0026162|Minerals|minerals
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6217,6220|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|6234,6244|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6234,6244|false|false|false|C0028978|omeprazole|Omeprazole
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6254,6257|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|6254,6257|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6254,6257|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|SIMPLE_SEGMENT|6254,6257|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|6262,6272|false|false|false|C0074393|sertraline|Sertraline
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6262,6272|false|false|false|C0074393|sertraline|Sertraline
Drug|Organic Chemical|SIMPLE_SEGMENT|6293,6300|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6293,6300|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|6293,6300|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|6293,6302|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|6293,6302|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6293,6302|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|6293,6302|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6293,6302|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|6325,6335|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6325,6335|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6325,6342|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6325,6342|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6336,6342|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6336,6342|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6336,6342|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|6336,6342|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6336,6342|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Idea or Concept|SIMPLE_SEGMENT|6391,6395|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|SIMPLE_SEGMENT|6396,6403|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|SIMPLE_SEGMENT|6396,6403|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6396,6403|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|SIMPLE_SEGMENT|6404,6418|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6404,6418|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|SIMPLE_SEGMENT|6420,6424|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|SIMPLE_SEGMENT|6420,6424|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|SIMPLE_SEGMENT|6420,6424|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|SIMPLE_SEGMENT|6430,6440|false|false|false|C0206460|enoxaparin|enoxaparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6430,6440|false|false|false|C0206460|enoxaparin|enoxaparin
Finding|Idea or Concept|SIMPLE_SEGMENT|6513,6520|false|true|false|C0807726|refill|Refills
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6527,6535|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|6527,6535|false|false|false|C0028040|nicotine|Nicotine
Drug|Clinical Drug|SIMPLE_SEGMENT|6527,6541|false|false|false|C0358855|Nicotine Transdermal Patch|Nicotine Patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6536,6541|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|SIMPLE_SEGMENT|6536,6541|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6562,6570|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|6562,6570|false|false|false|C0028040|nicotine|nicotine
Drug|Organic Chemical|SIMPLE_SEGMENT|6572,6580|false|false|false|C0701369|Nicoderm|Nicoderm
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6572,6580|false|false|false|C0701369|Nicoderm|Nicoderm
Drug|Organic Chemical|SIMPLE_SEGMENT|6572,6583|false|false|false|C1170429|Nicoderm C-Q|Nicoderm CQ
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6572,6583|false|false|false|C1170429|Nicoderm C-Q|Nicoderm CQ
Finding|Functional Concept|SIMPLE_SEGMENT|6599,6604|false|false|false|C1632850;C1879355;C4048755;C4521676|Apply;Apply (administration method);Apply (instruction)|Apply
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6609,6614|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|patch
Finding|Finding|SIMPLE_SEGMENT|6609,6614|false|false|false|C0332461|Plaque (lesion)|patch
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6632,6637|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Finding|Finding|SIMPLE_SEGMENT|6632,6637|false|false|false|C0332461|Plaque (lesion)|Patch
Finding|Idea or Concept|SIMPLE_SEGMENT|6638,6645|false|false|false|C0807726|refill|Refills
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6652,6660|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|6652,6660|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6652,6660|false|false|false|C0043031|warfarin|Warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|6682,6690|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|6682,6690|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6682,6690|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|6692,6700|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6692,6700|false|false|false|C0699129|Coumadin|Coumadin
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6709,6715|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|SIMPLE_SEGMENT|6719,6727|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6722,6727|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|6722,6727|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|SIMPLE_SEGMENT|6735,6739|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|SIMPLE_SEGMENT|6735,6739|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6746,6752|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|SIMPLE_SEGMENT|6753,6760|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|SIMPLE_SEGMENT|6767,6776|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6767,6776|false|false|false|C0001927|albuterol|albuterol
Drug|Organic Chemical|SIMPLE_SEGMENT|6767,6784|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6767,6784|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|6777,6784|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|SIMPLE_SEGMENT|6777,6784|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6777,6784|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Finding|Functional Concept|SIMPLE_SEGMENT|6802,6812|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|SIMPLE_SEGMENT|6802,6812|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Gene or Genome|SIMPLE_SEGMENT|6819,6822|false|false|false|C1422467|CIAO3 gene|prn
Finding|Sign or Symptom|SIMPLE_SEGMENT|6824,6832|false|false|false|C0043144|Wheezing|wheezing
Finding|Classification|SIMPLE_SEGMENT|6838,6848|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|6838,6848|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Gene or Genome|SIMPLE_SEGMENT|6849,6852|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Finding|Intellectual Product|SIMPLE_SEGMENT|6849,6852|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|Lab
Event|Occupational Activity|SIMPLE_SEGMENT|6853,6857|false|false|false|C0043227|Work|Work
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6871,6874|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6871,6874|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6871,6874|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6884,6887|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|6884,6887|false|false|false|C0020725;C0021122|Disruptive, Impulse Control, and Conduct Disorders;Type II Mucolipidosis|ICD
Finding|Gene or Genome|SIMPLE_SEGMENT|6884,6887|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|6884,6887|false|false|false|C0870733;C5891008|GNPTAB wt Allele;International Classification of Diseases|ICD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6884,6887|false|false|false|C5575277|Icd Regimen|ICD
Finding|Intellectual Product|SIMPLE_SEGMENT|6884,6889|false|false|false|C1137111;C2346503|ICD-9;International Classification of Diseases, Ninth Revision|ICD-9
Finding|Finding|SIMPLE_SEGMENT|6910,6916|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|SIMPLE_SEGMENT|6910,6916|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|SIMPLE_SEGMENT|6910,6916|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Body Substance|SIMPLE_SEGMENT|6938,6947|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6938,6947|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6938,6947|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6938,6947|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6938,6959|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|6938,6959|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6948,6959|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|6948,6959|false|false|false|C0184758|Patient disposition|Disposition
Finding|Idea or Concept|SIMPLE_SEGMENT|6961,6965|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|6961,6965|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|6961,6965|false|false|false|C1553498|home health encounter|Home
Finding|Body Substance|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6968,6977|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|6968,6987|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6978,6987|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6978,6987|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6978,6987|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6978,6987|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6989,7006|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6997,7006|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|6997,7006|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|6997,7006|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6997,7006|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7008,7017|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7008,7017|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|7008,7017|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7008,7026|false|false|false|C0034065|Pulmonary Embolism|Pulmonary embolism
Finding|Finding|SIMPLE_SEGMENT|7018,7026|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|7018,7026|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7028,7037|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|7028,7037|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7028,7047|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|SIMPLE_SEGMENT|7028,7047|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7038,7047|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7038,7047|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7038,7047|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7038,7047|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7049,7077|false|false|false|C1510431|Superficial Thrombophlebitis|Superficial thrombophlebitis
Finding|Pathologic Function|SIMPLE_SEGMENT|7061,7077|false|false|false|C0040046|Thrombophlebitis|thrombophlebitis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7079,7096|false|false|false|C0801658||Primary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7087,7096|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7087,7096|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7087,7096|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7087,7096|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7098,7107|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7098,7107|false|false|false|C2707265||Pulmonary
Finding|Finding|SIMPLE_SEGMENT|7098,7107|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|SIMPLE_SEGMENT|7098,7116|false|false|false|C0034065|Pulmonary Embolism|Pulmonary embolism
Finding|Finding|SIMPLE_SEGMENT|7108,7116|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|7108,7116|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7118,7127|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|7118,7127|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7118,7137|false|false|false|C4255018||Secondary Diagnosis
Finding|Finding|SIMPLE_SEGMENT|7118,7137|false|false|false|C0332138|Secondary diagnosis|Secondary Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7128,7137|false|false|false|C0945731||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|7128,7137|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|7128,7137|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7128,7137|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7139,7167|false|false|false|C1510431|Superficial Thrombophlebitis|Superficial thrombophlebitis
Finding|Pathologic Function|SIMPLE_SEGMENT|7151,7167|false|false|false|C0040046|Thrombophlebitis|thrombophlebitis
Finding|Body Substance|SIMPLE_SEGMENT|7171,7180|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7171,7180|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7171,7180|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7171,7180|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7181,7190|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7181,7190|false|false|false|C0012634|Disease|Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|7181,7190|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|7192,7198|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7192,7205|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|7192,7205|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7199,7205|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7199,7205|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7207,7212|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|SIMPLE_SEGMENT|7217,7225|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7227,7249|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7227,7249|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|7236,7249|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|7236,7249|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7251,7256|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|7251,7256|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7251,7256|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|SIMPLE_SEGMENT|7251,7256|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7251,7256|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|7251,7256|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|7261,7272|false|false|false|C1704675|Interaction|interactive
Event|Activity|SIMPLE_SEGMENT|7274,7282|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|7274,7282|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|SIMPLE_SEGMENT|7274,7282|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7283,7289|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|7283,7289|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|SIMPLE_SEGMENT|7291,7301|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|SIMPLE_SEGMENT|7291,7301|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|SIMPLE_SEGMENT|7291,7301|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|SIMPLE_SEGMENT|7291,7301|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Finding|SIMPLE_SEGMENT|7304,7315|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|SIMPLE_SEGMENT|7304,7315|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Body Substance|SIMPLE_SEGMENT|7320,7329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|7320,7329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|7320,7329|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|7320,7329|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7320,7342|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7320,7342|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|7320,7342|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7330,7342|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|7330,7342|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|7344,7348|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|SIMPLE_SEGMENT|7368,7376|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|7368,7376|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7440,7449|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7440,7449|false|false|false|C2707265||pulmonary
Finding|Finding|SIMPLE_SEGMENT|7440,7449|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Finding|SIMPLE_SEGMENT|7451,7459|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|SIMPLE_SEGMENT|7451,7459|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7461,7466|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|7461,7466|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|7461,7471|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|SIMPLE_SEGMENT|7467,7471|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7467,7471|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|SIMPLE_SEGMENT|7467,7471|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7479,7484|false|false|false|C0024109|Lung|lungs
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7503,7508|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|SIMPLE_SEGMENT|7503,7508|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|7503,7513|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|SIMPLE_SEGMENT|7509,7513|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7509,7513|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|SIMPLE_SEGMENT|7509,7513|false|false|false|C0302148|Blood Clot|clot
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7546,7554|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Finding|Classification|SIMPLE_SEGMENT|7594,7604|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7594,7604|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7639,7649|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7639,7649|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Intellectual Product|SIMPLE_SEGMENT|7661,7673|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|SIMPLE_SEGMENT|7661,7673|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|SIMPLE_SEGMENT|7669,7673|false|false|false|C1947933|care activity|care
Finding|Finding|SIMPLE_SEGMENT|7669,7673|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7669,7673|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|7674,7680|false|false|false|C2348314|Doctor - Title|doctor
Finding|Finding|SIMPLE_SEGMENT|7713,7719|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|7713,7719|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Pathologic Function|SIMPLE_SEGMENT|7792,7800|false|false|false|C0002940|Aneurysm|aneurysm
Finding|Functional Concept|SIMPLE_SEGMENT|7836,7842|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Gene or Genome|SIMPLE_SEGMENT|7843,7846|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7843,7846|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|7843,7846|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7855,7860|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7855,7860|false|false|false|C0006111|Brain Diseases|brain
Finding|Gene or Genome|SIMPLE_SEGMENT|7892,7895|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7892,7895|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|SIMPLE_SEGMENT|7892,7895|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7963,7968|false|false|false|C1410088|Still|still
Finding|Idea or Concept|SIMPLE_SEGMENT|8015,8024|false|false|false|C0549178|Continuous|continued
Event|Activity|SIMPLE_SEGMENT|8025,8033|false|false|false|C0237820||recovery
Finding|Organism Function|SIMPLE_SEGMENT|8025,8033|false|false|false|C2004454|Recovery - healing process|recovery
Procedure|Health Care Activity|SIMPLE_SEGMENT|8064,8072|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8073,8085|false|false|false|C3263700||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|8073,8085|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

