 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|46,55|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|46,55|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|46,60|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|80,89|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|80,89|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|80,89|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|80,94|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|112,117|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|136,139|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|136,139|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|147,154|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|147,154|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|156,168|false|false|false|||NEUROSURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|156,168|false|false|false|C0524850|Neurosurgical Procedures|NEUROSURGERY
Disorder|Injury or Poisoning|Allergies|183,194|false|false|false|C0161486;C2876539|Poisoning by penicillin;Poisoning by, adverse effect of and underdosing of penicillins|Penicillins
Drug|Antibiotic|Allergies|183,194|false|false|false|C0030842|penicillins|Penicillins
Drug|Organic Chemical|Allergies|183,194|false|false|false|C0030842|penicillins|Penicillins
Event|Event|Allergies|183,194|false|false|false|||Penicillins
Finding|Pathologic Function|Allergies|183,194|false|false|false|C0413443|Adverse reaction to penicillins|Penicillins
Drug|Organic Chemical|Allergies|197,202|false|false|false|C0376414|Paxil|Paxil
Drug|Pharmacologic Substance|Allergies|197,202|false|false|false|C0376414|Paxil|Paxil
Drug|Organic Chemical|Allergies|205,215|false|false|false|C0085934|Wellbutrin|Wellbutrin
Drug|Pharmacologic Substance|Allergies|205,215|false|false|false|C0085934|Wellbutrin|Wellbutrin
Event|Event|Allergies|218,227|false|false|false|||Attending
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|261,271|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Chief Complaint|272,280|false|false|false|||hardware
Finding|Classification|Chief Complaint|283,288|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|289,297|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|289,297|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|301,319|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|310,319|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|310,319|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|310,319|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|310,319|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|310,319|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Injury or Poisoning|Chief Complaint|321,326|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Chief Complaint|321,326|false|false|false|||wound
Finding|Body Substance|Chief Complaint|321,326|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Chief Complaint|321,326|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Chief Complaint|321,326|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Chief Complaint|327,335|false|false|false|||revision
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|327,335|false|false|false|C0558347;C1527075|Revision procedure;Surgical revision|revision
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|340,356|false|false|false|C5453054|Hardware Removal|hardware removal
Event|Activity|Chief Complaint|349,356|false|false|false|C1883720|Removing (action)|removal
Event|Event|Chief Complaint|349,356|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|349,356|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Finding|Idea or Concept|History of Present Illness|402,406|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|402,406|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|History of Present Illness|407,410|false|false|false|||old
Finding|Finding|History of Present Illness|423,436|false|false|false|C0455610|History of surgery|prior surgery
Event|Event|History of Present Illness|429,436|false|false|false|||surgery
Finding|Finding|History of Present Illness|429,436|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|429,436|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|429,436|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|429,436|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|443,451|false|false|false|||includes
Finding|Functional Concept|History of Present Illness|452,457|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Neoplastic Process|History of Present Illness|467,489|false|false|false|C0334579|Anaplastic astrocytoma|anaplastic astrocytoma
Disorder|Neoplastic Process|History of Present Illness|478,489|false|false|false|C0004114|Astrocytoma|astrocytoma
Event|Event|History of Present Illness|478,489|false|false|false|||astrocytoma
Event|Event|History of Present Illness|495,505|false|false|false|||Craniotomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|495,505|false|false|false|C0010280|Craniotomy|Craniotomy
Event|Event|History of Present Illness|510,519|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|510,519|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Finding|Functional Concept|History of Present Illness|558,566|false|false|false|C1314939|Involvement with|involved
Finding|Conceptual Entity|History of Present Illness|567,572|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|field
Procedure|Health Care Activity|History of Present Illness|567,572|false|false|false|C1553496|field - patient encounter|field
Event|Event|History of Present Illness|573,584|false|false|false|||irradiation
Phenomenon|Natural Phenomenon or Process|History of Present Illness|573,584|false|false|false|C0851346;C1282930|Irradiation (physical force);Radiation|irradiation
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|573,584|false|false|false|C1522449|Radiation therapy (procedure)|irradiation
Event|Event|History of Present Illness|612,618|false|false|false|||cycles
Drug|Organic Chemical|History of Present Illness|622,629|false|false|false|C0876179|Temodar|Temodar
Drug|Pharmacologic Substance|History of Present Illness|622,629|false|false|false|C0876179|Temodar|Temodar
Event|Event|History of Present Illness|630,635|false|false|false|||ended
Finding|Functional Concept|History of Present Illness|646,652|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Idea or Concept|History of Present Illness|646,652|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Finding|Intellectual Product|History of Present Illness|646,652|false|false|false|C1522484;C1561503;C1705190|Precision - second;Second Suffix;metastatic qualifier|second
Event|Event|History of Present Illness|653,663|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|653,663|false|false|false|C0010280|Craniotomy|craniotomy
Disorder|Neoplastic Process|History of Present Illness|668,673|false|false|false|C0027651|Neoplasms|tumor
Event|Event|History of Present Illness|668,673|false|false|false|||tumor
Finding|Finding|History of Present Illness|668,673|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|History of Present Illness|668,673|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Disorder|Neoplastic Process|History of Present Illness|674,684|false|false|false|C1458156|Recurrent Malignant Neoplasm|recurrence
Event|Event|History of Present Illness|674,684|false|false|false|||recurrence
Finding|Pathologic Function|History of Present Illness|674,684|false|false|false|C2825055|Recurrence (disease attribute)|recurrence
Phenomenon|Phenomenon or Process|History of Present Illness|674,684|false|false|false|C0034897|Recurrence|recurrence
Anatomy|Body Location or Region|History of Present Illness|715,718|false|false|false|C5239890|area PCV|PCV
Disorder|Virus|History of Present Illness|715,718|false|false|false|C0206411|Porcine circovirus|PCV
Drug|Nucleic Acid, Nucleoside, or Nucleotide|History of Present Illness|715,718|false|false|false|C0164815|penciclovir|PCV
Drug|Pharmacologic Substance|History of Present Illness|715,718|false|false|false|C0164815|penciclovir|PCV
Event|Event|History of Present Illness|715,718|false|false|false|||PCV
Procedure|Laboratory Procedure|History of Present Illness|715,718|false|false|false|C0018935;C0070167;C1882252|Hematocrit Measurement;Procarbazine-Lomustine-Vincristine (PCV) Regimen;lomustine/procarbazine/vincristine|PCV
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|715,718|false|false|false|C0018935;C0070167;C1882252|Hematocrit Measurement;Procarbazine-Lomustine-Vincristine (PCV) Regimen;lomustine/procarbazine/vincristine|PCV
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|719,723|false|false|false|C0376161|Comb (body structure)|comb
Drug|Organic Chemical|History of Present Illness|719,723|false|false|false|C0278789|Combid|comb
Drug|Pharmacologic Substance|History of Present Illness|719,723|false|false|false|C0278789|Combid|comb
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|719,723|false|false|false|C0279325;C0280054|bleomycin/cyclophosphamide/methotrexate/vincristine protocol;bleomycin/cyclophosphamide/semustine/vincristine protocol|comb
Event|Event|History of Present Illness|724,729|false|false|false|||chemo
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|724,729|false|false|false|C0392920;C3665472|Chemotherapy;Chemotherapy Regimen|chemo
Finding|Body Substance|History of Present Illness|749,756|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|749,756|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|749,756|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|757,765|false|false|false|||presents
Finding|Idea or Concept|History of Present Illness|781,786|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|781,786|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|History of Present Illness|787,794|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|787,794|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|787,794|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|787,794|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|787,797|false|false|false|C0262926|Medical History|history of
Event|Event|History of Present Illness|798,806|false|false|false|||pruritus
Finding|Sign or Symptom|History of Present Illness|798,806|false|false|false|C0033774|Pruritus|pruritus
Anatomy|Body Location or Region|History of Present Illness|825,829|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|825,829|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|825,829|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|825,829|false|false|false|C0876917|Procedure on head|head
Event|Event|History of Present Illness|836,843|false|false|false|||reports
Event|Event|History of Present Illness|869,873|false|false|false|||look
Anatomy|Body Location or Region|History of Present Illness|892,896|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|892,896|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|892,896|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|892,896|false|false|false|C0876917|Procedure on head|head
Finding|Gene or Genome|History of Present Illness|906,909|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|914,917|false|false|false|||saw
Drug|Inorganic Chemical|History of Present Illness|923,928|false|false|false|C0025552|Metals|metal
Event|Event|History of Present Illness|929,937|false|false|false|||hardware
Finding|Finding|History of Present Illness|947,960|false|false|false|C0455610|History of surgery|prior surgery
Event|Event|History of Present Illness|953,960|false|false|false|||surgery
Finding|Finding|History of Present Illness|953,960|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|953,960|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|953,960|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|953,960|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|965,972|false|false|false|||present
Finding|Finding|History of Present Illness|965,972|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|History of Present Illness|965,972|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Body Substance|History of Present Illness|979,986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|979,986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|979,986|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1003,1012|false|false|false|||presented
Finding|Idea or Concept|History of Present Illness|1022,1027|false|false|false|C1550012|Local Remote Control State - Local|local
Event|Event|History of Present Illness|1028,1037|false|false|false|||Emergency
Finding|Finding|History of Present Illness|1028,1037|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|History of Present Illness|1028,1037|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|History of Present Illness|1028,1037|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|History of Present Illness|1028,1037|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|History of Present Illness|1028,1037|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|History of Present Illness|1028,1037|false|false|false|C1553500|emergency encounter|Emergency
Event|Event|History of Present Illness|1046,1050|false|false|false|||told
Finding|Body Substance|History of Present Illness|1075,1082|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1075,1082|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1075,1082|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1083,1089|false|false|false|||denies
Event|Event|History of Present Illness|1090,1095|false|false|false|||fever
Finding|Finding|History of Present Illness|1090,1095|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1090,1095|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1097,1103|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1097,1103|true|false|false|C0085593|Chills|chills
Attribute|Clinical Attribute|History of Present Illness|1105,1111|false|false|false|C4255480||nausea
Finding|Sign or Symptom|History of Present Illness|1105,1111|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|1105,1120|true|false|false|C0027498|Nausea and vomiting|nausea vomiting
Event|Event|History of Present Illness|1112,1120|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1112,1120|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1122,1128|false|false|false|||nuchal
Event|Event|History of Present Illness|1129,1137|false|false|false|||rigidity
Finding|Sign or Symptom|History of Present Illness|1129,1137|false|false|false|C0026837|Muscle Rigidity|rigidity
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1129,1137|false|false|false|C0700109|plastic property - rigidity|rigidity
Event|Event|History of Present Illness|1139,1147|false|false|false|||numbness
Finding|Finding|History of Present Illness|1139,1147|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1139,1147|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Finding|History of Present Illness|1139,1159|false|false|false|C3842982|Numbness or tingling|numbness or tingling
Disorder|Disease or Syndrome|History of Present Illness|1151,1159|false|false|false|C0030554|Paresthesia|tingling
Event|Event|History of Present Illness|1151,1159|false|false|false|||tingling
Finding|Sign or Symptom|History of Present Illness|1151,1159|false|false|false|C2242996|Has tingling sensation|tingling
Finding|Sign or Symptom|History of Present Illness|1151,1169|false|false|false|C2242996|Has tingling sensation|tingling sensation
Event|Event|History of Present Illness|1160,1169|false|false|false|||sensation
Finding|Finding|History of Present Illness|1160,1169|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|1160,1169|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|1160,1169|false|false|false|C2229507|sensory exam|sensation
Attribute|Clinical Attribute|History of Present Illness|1171,1177|false|false|false|C2707266||vision
Event|Event|History of Present Illness|1171,1177|false|false|false|||vision
Finding|Organism Function|History of Present Illness|1171,1177|false|false|false|C0042789|Vision|vision
Event|Event|History of Present Illness|1181,1188|false|false|false|||hearing
Finding|Finding|History of Present Illness|1181,1188|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|History of Present Illness|1181,1188|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Event|Event|History of Present Illness|1189,1196|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|1189,1196|false|false|false|C0392747|Changing|changes
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1198,1203|false|false|false|C0021853|Intestines|bowel
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1207,1214|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|1207,1214|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1207,1214|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Disease or Syndrome|History of Present Illness|1207,1227|false|false|false|C3668875|Urinary incontinence due to bladder problem|bladder incontinence
Finding|Finding|History of Present Illness|1207,1227|false|false|false|C0042024;C2188450|Urinary Incontinence;urinary incontinence by exam|bladder incontinence
Finding|Pathologic Function|History of Present Illness|1207,1227|false|false|false|C0042024;C2188450|Urinary Incontinence;urinary incontinence by exam|bladder incontinence
Disorder|Disease or Syndrome|History of Present Illness|1215,1227|false|false|false|C0021167|Incontinence|incontinence
Event|Event|History of Present Illness|1215,1227|false|false|false|||incontinence
Event|Event|History of Present Illness|1234,1240|false|false|false|||denies
Finding|Finding|History of Present Illness|1241,1244|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|History of Present Illness|1241,1244|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|History of Present Illness|1241,1250|true|false|false|C0746890|new onset|new onset
Event|Event|History of Present Illness|1245,1250|false|false|false|||onset
Event|Event|History of Present Illness|1251,1259|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1251,1259|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|History of Present Illness|1266,1273|false|false|false|||reports
Drug|Biomedical or Dental Material|History of Present Illness|1274,1282|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1274,1282|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1274,1282|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|History of Present Illness|1283,1290|false|false|false|||tremors
Finding|Sign or Symptom|History of Present Illness|1283,1290|false|false|false|C0040822|Tremor|tremors
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1294,1298|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|History of Present Illness|1294,1298|false|false|false|C5782111||arms
Disorder|Neoplastic Process|History of Present Illness|1294,1298|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Finding|Gene or Genome|History of Present Illness|1294,1298|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|History of Present Illness|1294,1298|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Disorder|Disease or Syndrome|History of Present Illness|1310,1322|false|false|false|C0020550|Hyperthyroidism|hyperthyroid
Event|Event|History of Present Illness|1310,1322|false|false|false|||hyperthyroid
Disorder|Disease or Syndrome|History of Present Illness|1323,1330|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|1323,1330|false|false|false|||disease
Drug|Biomedical or Dental Material|History of Present Illness|1335,1343|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1335,1343|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1335,1343|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Functional Concept|History of Present Illness|1344,1348|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|History of Present Illness|1344,1363|false|false|false|C0457436|Left hemiparesis|left sided weakness
Event|Event|History of Present Illness|1355,1363|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|1355,1363|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Idea or Concept|History of Present Illness|1374,1381|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1382,1389|false|false|false|||surgery
Finding|Finding|History of Present Illness|1382,1389|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|History of Present Illness|1382,1389|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|History of Present Illness|1382,1389|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1382,1389|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|History of Present Illness|1405,1413|false|false|false|||ambulate
Finding|Finding|History of Present Illness|1405,1413|false|true|false|C4036205|Ambulate|ambulate
Finding|Functional Concept|Past Medical History|1454,1459|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Neoplastic Process|Past Medical History|1469,1491|false|false|false|C0334579|Anaplastic astrocytoma|anaplastic astrocytoma
Disorder|Neoplastic Process|Past Medical History|1480,1491|false|true|false|C0004114|Astrocytoma|astrocytoma
Event|Event|Past Medical History|1480,1491|false|false|false|||astrocytoma
Event|Event|Past Medical History|1492,1502|false|false|false|||Craniotomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1492,1502|false|false|false|C0010280|Craniotomy|Craniotomy
Event|Event|Past Medical History|1525,1536|false|false|false|||irradiation
Phenomenon|Natural Phenomenon or Process|Past Medical History|1525,1536|false|false|false|C0851346;C1282930|Irradiation (physical force);Radiation|irradiation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1525,1536|false|false|false|C1522449|Radiation therapy (procedure)|irradiation
Event|Event|Past Medical History|1563,1569|false|false|false|||cycles
Drug|Organic Chemical|Past Medical History|1573,1580|false|false|false|C0876179|Temodar|Temodar
Drug|Pharmacologic Substance|Past Medical History|1573,1580|false|false|false|C0876179|Temodar|Temodar
Event|Event|Past Medical History|1581,1586|false|false|false|||ended
Event|Event|Past Medical History|1591,1601|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1591,1601|false|false|false|C0010280|Craniotomy|craniotomy
Disorder|Disease or Syndrome|Past Medical History|1658,1665|false|false|false|C0012634|Disease|disease
Event|Event|Past Medical History|1658,1665|false|false|false|||disease
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1677,1691|false|false|false|C0520483|Tubal Ligation|tubal ligation
Event|Event|Past Medical History|1683,1691|false|false|false|||ligation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1683,1691|false|false|false|C0023690|Ligation|ligation
Event|Event|Past Medical History|1692,1705|false|false|false|||tonsillectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1692,1705|false|false|false|C0040423|Tonsillectomy|tonsillectomy
Disorder|Disease or Syndrome|Past Medical History|1707,1717|false|false|false|C0006277;C0149514|Acute bronchitis;Bronchitis|bronchitis
Event|Event|Past Medical History|1707,1717|false|false|false|||bronchitis
Disorder|Mental or Behavioral Dysfunction|Past Medical History|1719,1729|false|false|false|C0011570;C0011581;C0344315;C0812393|Cancer patients and suicide and depression;Depressed mood;Depressive disorder;Mental Depression|depression
Event|Event|Past Medical History|1719,1729|false|false|false|||depression
Finding|Functional Concept|Past Medical History|1719,1729|false|false|false|C0460137;C1579931|Depression - motion|depression
Finding|Sign or Symptom|Past Medical History|1719,1729|false|false|false|C0460137;C1579931|Depression - motion|depression
Event|Event|Past Medical History|1731,1739|false|false|false|||seizures
Finding|Sign or Symptom|Past Medical History|1731,1739|false|false|false|C0036572|Seizures|seizures
Event|Event|General Exam|1856,1859|false|false|false|||Gen
Finding|Classification|General Exam|1856,1859|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1856,1859|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1868,1879|false|false|false|||comfortable
Finding|Finding|General Exam|1868,1879|false|false|false|C5546696|Feeling comfortable|comfortable
Disorder|Disease or Syndrome|General Exam|1881,1884|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1881,1884|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1881,1884|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1881,1884|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1881,1884|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|1881,1884|false|false|false|||NAD
Finding|Finding|General Exam|1881,1884|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1886,1891|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|1893,1899|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|1920,1924|false|false|false|||EOMs
Finding|Functional Concept|General Exam|1920,1924|false|false|false|C0241886|Extraocular|EOMs
Event|Event|General Exam|1926,1932|false|false|false|||intact
Finding|Finding|General Exam|1926,1932|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Location or Region|General Exam|1933,1937|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|1933,1937|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|1933,1937|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|1939,1945|false|false|false|||Supple
Finding|Functional Concept|General Exam|1939,1945|false|false|false|C0332254|Supple|Supple
Event|Event|General Exam|1955,1959|false|false|false|||Warm
Finding|Finding|General Exam|1955,1959|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1955,1959|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1964,1968|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1969,1977|false|false|false|||perfused
Anatomy|Body Part, Organ, or Organ Component|General Exam|1979,1983|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|General Exam|1979,1983|false|false|false|C5782111||arms
Disorder|Neoplastic Process|General Exam|1979,1983|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|General Exam|1979,1983|false|false|false|||arms
Finding|Gene or Genome|General Exam|1979,1983|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|General Exam|1979,1983|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|General Exam|1984,1989|false|false|false|||hands
Event|Event|General Exam|1990,1999|false|false|false|||tremulous
Finding|Sign or Symptom|General Exam|1990,1999|false|false|false|C0234369|Trembling|tremulous
Finding|Body Substance|General Exam|2002,2009|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|2002,2009|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|2002,2009|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|2010,2016|false|false|false|||states
Drug|Biomedical or Dental Material|General Exam|2029,2037|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|2029,2037|false|false|false|||baseline
Finding|Idea or Concept|General Exam|2029,2037|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|General Exam|2045,2057|false|false|false|C0020550|Hyperthyroidism|hyperthyroid
Disorder|Disease or Syndrome|General Exam|2058,2065|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|2058,2065|false|false|false|||disease
Finding|Mental Process|General Exam|2074,2080|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|2074,2087|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|2074,2087|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|2081,2087|false|false|false|C5889824||status
Event|Event|General Exam|2081,2087|false|false|false|||status
Finding|Idea or Concept|General Exam|2081,2087|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|2089,2094|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|2099,2104|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|2099,2104|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|2099,2104|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|2099,2104|false|false|false|||alert
Finding|Finding|General Exam|2099,2104|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|2099,2104|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|2099,2104|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|2106,2117|false|false|false|||cooperative
Event|Event|General Exam|2123,2127|false|false|false|||exam
Finding|Functional Concept|General Exam|2123,2127|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|2123,2127|false|false|false|C0582103|Medical Examination|exam
Event|Event|General Exam|2129,2135|false|false|false|||normal
Event|Event|General Exam|2136,2142|false|false|false|||affect
Finding|Mental Process|General Exam|2136,2142|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|2136,2142|false|false|false|C2237113|assessment of affect|affect
Event|Event|General Exam|2144,2155|false|false|false|||Orientation
Finding|Mental Process|General Exam|2144,2155|false|false|false|C0029266|Mental Orientation|Orientation
Event|Event|General Exam|2157,2165|false|false|false|||Oriented
Finding|Finding|General Exam|2157,2165|false|false|false|C1961028|Oriented to place|Oriented
Finding|Finding|General Exam|2157,2175|false|false|false|C1961030|Oriented to person|Oriented to person
Attribute|Clinical Attribute|General Exam|2169,2175|false|false|false|C5890614||person
Event|Event|General Exam|2169,2175|false|false|false|||person
Finding|Intellectual Product|General Exam|2169,2175|false|false|false|C1522390|Person Info|person
Event|Activity|General Exam|2177,2182|false|false|false|C1882509|put - instruction imperative|place
Event|Event|General Exam|2177,2182|false|false|false|||place
Finding|Functional Concept|General Exam|2177,2182|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|2177,2182|false|false|false|C1533810||place
Event|Event|General Exam|2194,2200|false|false|false|||Recall
Event|Governmental or Regulatory Activity|General Exam|2194,2200|false|false|false|C1705180|Recall (activity)|Recall
Finding|Mental Process|General Exam|2194,2200|false|false|false|C0034770|Mental Recall|Recall
Event|Event|General Exam|2206,2213|false|false|false|||objects
Procedure|Therapeutic or Preventive Procedure|General Exam|2217,2226|false|false|false|C0886384|5 minutes Office visit|5 minutes
Event|Event|General Exam|2219,2226|false|false|false|||minutes
Attribute|Clinical Attribute|General Exam|2228,2236|false|false|false|C2706915||Language
Event|Event|General Exam|2228,2236|false|false|false|||Language
Finding|Intellectual Product|General Exam|2228,2236|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|2238,2244|false|false|false|||Speech
Finding|Organism Function|General Exam|2238,2244|false|false|false|C0037817|Speech|Speech
Procedure|Diagnostic Procedure|General Exam|2238,2244|false|false|false|C0846595|Speech assessment|Speech
Finding|Idea or Concept|General Exam|2257,2261|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|2262,2275|false|false|false|||comprehension
Finding|Mental Process|General Exam|2262,2275|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|2280,2290|false|false|false|||repetition
Finding|Finding|General Exam|2280,2290|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|2280,2290|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|2292,2298|false|false|false|||Naming
Finding|Mental Process|General Exam|2292,2298|false|false|false|C0233735|Naming (function)|Naming
Event|Event|General Exam|2299,2305|false|false|false|||intact
Finding|Finding|General Exam|2299,2305|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Mental or Behavioral Dysfunction|General Exam|2310,2320|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|2310,2320|false|false|false|||dysarthria
Event|Event|General Exam|2335,2341|false|false|false|||errors
Anatomy|Body Part, Organ, or Organ Component|General Exam|2344,2351|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|2344,2358|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|2344,2358|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|2352,2358|false|false|false|C0027740|Nerve|Nerves
Event|Event|General Exam|2367,2373|false|false|false|||tested
Anatomy|Body Part, Organ, or Organ Component|General Exam|2378,2384|false|false|false|C0034121|Pupil|Pupils
Event|Event|General Exam|2393,2398|false|false|false|||round
Event|Event|General Exam|2403,2411|false|false|false|||reactive
Procedure|Therapeutic or Preventive Procedure|General Exam|2403,2411|false|false|false|C4722408|Reactive Therapy|reactive
Finding|Finding|General Exam|2403,2420|false|false|false|C4068744|Reactive to light|reactive to light
Drug|Amino Acid, Peptide, or Protein|General Exam|2415,2420|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2415,2420|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|2415,2420|false|false|false|||light
Finding|Finding|General Exam|2415,2420|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2415,2420|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2415,2420|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2415,2420|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2415,2420|false|false|false|C0031765|Phototherapy|light
Finding|Functional Concept|General Exam|2446,2452|false|false|false|C0234621|Visual|Visual
Event|Event|General Exam|2453,2459|false|false|false|||fields
Event|Event|General Exam|2464,2468|false|false|false|||full
Event|Event|General Exam|2472,2485|false|false|false|||confrontation
Finding|Finding|General Exam|2472,2485|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|2472,2485|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|2472,2485|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Finding|Functional Concept|General Exam|2500,2511|false|false|false|C0241886|Extraocular|Extraocular
Procedure|Diagnostic Procedure|General Exam|2500,2521|false|false|false|C2228439|examination of extraocular movements|Extraocular movements
Event|Event|General Exam|2512,2521|false|false|false|||movements
Finding|Organism Function|General Exam|2512,2521|false|false|false|C0026649|Movement|movements
Event|Event|General Exam|2522,2528|false|false|false|||intact
Finding|Finding|General Exam|2522,2528|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|2549,2558|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|2549,2558|false|false|false|||nystagmus
Anatomy|Body Part, Organ, or Organ Component|General Exam|2563,2566|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|2563,2566|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|2568,2574|false|false|false|C0015450|Face|Facial
Event|Event|General Exam|2575,2583|false|false|false|||strength
Finding|Idea or Concept|General Exam|2575,2583|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|2588,2597|false|false|false|||sensation
Finding|Finding|General Exam|2588,2597|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2588,2597|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2588,2597|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|2598,2604|false|false|false|||intact
Finding|Finding|General Exam|2598,2604|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2609,2618|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|2609,2618|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|2609,2618|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2620,2624|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|2620,2624|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|2620,2624|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Event|Event|General Exam|2626,2633|false|false|false|||Hearing
Finding|Finding|General Exam|2626,2633|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|2626,2633|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|2634,2640|false|false|false|||intact
Finding|Finding|General Exam|2634,2640|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|2644,2649|false|false|false|||voice
Finding|Idea or Concept|General Exam|2644,2649|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Intellectual Product|General Exam|2644,2649|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Finding|Organism Function|General Exam|2644,2649|false|false|false|C0042939;C1547570;C4281800|Authorization Mode - Voice;Voice;Voice G-code|voice
Anatomy|Body Part, Organ, or Organ Component|General Exam|2658,2665|false|false|false|C0700374|Palate|Palatal
Event|Event|General Exam|2666,2675|false|false|false|||elevation
Procedure|Therapeutic or Preventive Procedure|General Exam|2666,2675|false|false|false|C0439775|Elevation procedure|elevation
Event|Event|General Exam|2676,2687|false|false|false|||symmetrical
Finding|Finding|General Exam|2676,2687|false|false|false|C0332516|Symmetrical|symmetrical
Anatomy|Body Part, Organ, or Organ Component|General Exam|2693,2712|false|false|false|C0224153|Structure of sternocleidomastoid muscle|Sternocleidomastoid
Anatomy|Body Part, Organ, or Organ Component|General Exam|2717,2726|false|false|false|C0224361|Structure of trapezius muscle|trapezius
Event|Event|General Exam|2727,2733|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|2752,2758|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|2752,2758|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Procedure|Health Care Activity|General Exam|2752,2758|false|false|false|C0872394|Procedure on tongue|Tongue
Finding|Finding|General Exam|2752,2766|false|false|false|C3693372|tongue midline|Tongue midline
Anatomy|Cell Component|General Exam|2759,2766|false|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|2775,2789|false|false|false|||fasciculations
Finding|Sign or Symptom|General Exam|2775,2789|true|false|false|C0015644|Muscular fasciculation|fasciculations
Event|Event|General Exam|2792,2797|false|false|false|||Motor
Finding|Functional Concept|General Exam|2792,2797|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|2806,2810|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|2806,2810|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|2806,2810|false|false|false|||bulk
Event|Event|General Exam|2815,2819|false|false|false|||tone
Finding|Finding|General Exam|2836,2844|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|General Exam|2836,2844|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Disorder|Disease or Syndrome|General Exam|2836,2854|true|false|false|C0013384|Dyskinetic syndrome|abnormal movements
Finding|Finding|General Exam|2836,2854|true|false|false|C0558189|Abnormal movement|abnormal movements
Event|Event|General Exam|2845,2854|false|false|false|||movements
Finding|Organism Function|General Exam|2845,2854|true|false|false|C0026649|Movement|movements
Event|Event|General Exam|2856,2863|false|false|false|||tremors
Finding|Sign or Symptom|General Exam|2856,2863|false|false|false|C0040822|Tremor|tremors
Finding|Idea or Concept|General Exam|2865,2873|false|false|false|C0808080|Strength (attribute)|Strength
Finding|Social Behavior|General Exam|2879,2884|false|false|false|C0032863|Power (Psychology)|power
Finding|Functional Concept|General Exam|2892,2897|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Event|Event|General Exam|2906,2910|false|false|false|||left
Finding|Functional Concept|General Exam|2906,2910|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Pathologic Function|General Exam|2915,2929|false|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|2924,2929|false|false|false|||drift
Event|Event|General Exam|2931,2940|false|false|false|||Sensation
Finding|Finding|General Exam|2931,2940|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Finding|Organ or Tissue Function|General Exam|2931,2940|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|Sensation
Procedure|Health Care Activity|General Exam|2931,2940|false|false|false|C2229507|sensory exam|Sensation
Event|Event|General Exam|2942,2948|false|false|false|||Intact
Finding|Finding|General Exam|2942,2948|false|false|false|C1554187|Gender Status - Intact|Intact
Drug|Amino Acid, Peptide, or Protein|General Exam|2952,2957|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|2952,2957|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|2952,2957|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|2952,2957|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|2952,2957|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|2952,2957|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|2952,2957|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|2952,2963|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|2958,2963|false|false|false|||touch
Finding|Mental Process|General Exam|2958,2963|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|2958,2963|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|2958,2963|false|false|false|C0152054|Therapeutic Touch|touch
Anatomy|Body Part, Organ, or Organ Component|General Exam|2978,2982|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|Toes
Event|Event|General Exam|2983,2992|false|false|false|||downgoing
Event|Event|General Exam|3006,3018|false|false|false|||Coordination
Finding|Functional Concept|General Exam|3006,3018|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|3006,3018|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|3006,3018|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|General Exam|3020,3026|false|false|false|||normal
Anatomy|Body Part, Organ, or Organ Component|General Exam|3030,3036|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Anatomy|Body Part, Organ, or Organ Component|General Exam|3042,3048|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Event|Event|General Exam|3056,3067|false|false|false|||alternating
Finding|Functional Concept|General Exam|3056,3067|false|false|false|C0332270|Alternating|alternating
Event|Event|General Exam|3068,3077|false|false|false|||movements
Finding|Organism Function|General Exam|3068,3077|false|false|false|C0026649|Movement|movements
Anatomy|Body Part, Organ, or Organ Component|General Exam|3079,3083|false|false|false|C0018870|Heel|heel
Anatomy|Body Location or Region|General Exam|3087,3091|false|false|false|C0230444|Shin|shin
Attribute|Clinical Attribute|General Exam|3114,3121|false|false|false|C0881943||CT Head
Procedure|Diagnostic Procedure|General Exam|3114,3121|false|false|false|C0202691|CAT scan of head|CT Head
Anatomy|Body Location or Region|General Exam|3117,3121|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Anatomy|Body Part, Organ, or Organ Component|General Exam|3117,3121|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|Head
Disorder|Disease or Syndrome|General Exam|3117,3121|false|false|false|C0362076|Problems with head|Head
Event|Event|General Exam|3117,3121|false|false|false|||Head
Procedure|Therapeutic or Preventive Procedure|General Exam|3117,3121|false|false|false|C0876917|Procedure on head|Head
Event|Event|General Exam|3128,3136|false|false|false|||evidence
Finding|Idea or Concept|General Exam|3128,3136|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|3128,3139|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|General Exam|3140,3147|true|false|false|C0000833|Abscess|abscess
Finding|Intellectual Product|General Exam|3140,3147|true|false|false|C1546533||abscess
Finding|Finding|General Exam|3140,3157|true|false|false|C4014106|Abscess formation|abscess formation
Event|Event|General Exam|3148,3157|false|false|false|||formation
Finding|Functional Concept|General Exam|3148,3157|true|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|General Exam|3148,3157|true|false|false|C0220781|Anabolism|formation
Finding|Intellectual Product|General Exam|3163,3169|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Attribute|Clinical Attribute|General Exam|3170,3180|false|false|false|C0550215||appearance
Event|Event|General Exam|3170,3180|false|false|false|||appearance
Procedure|Health Care Activity|General Exam|3170,3180|false|false|false|C2051406|patient appearance regarding mental status exam|appearance
Event|Event|General Exam|3198,3205|false|false|false|||changes
Finding|Functional Concept|General Exam|3198,3205|false|false|false|C0392747|Changing|changes
Drug|Organic Chemical|General Exam|3206,3213|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|General Exam|3206,3213|false|false|false|||related
Finding|Finding|General Exam|3206,3213|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|General Exam|3206,3213|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|General Exam|3217,3222|false|false|false|||right
Finding|Functional Concept|General Exam|3217,3222|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Finding|Finding|General Exam|3232,3236|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|General Exam|3232,3236|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|General Exam|3232,3236|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Event|Event|General Exam|3237,3246|false|false|false|||resection
Procedure|Therapeutic or Preventive Procedure|General Exam|3237,3246|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Disorder|Disease or Syndrome|General Exam|3261,3277|false|false|false|C0014068|Encephalomalacia|encephalomalacia
Event|Event|General Exam|3261,3277|false|false|false|||encephalomalacia
Attribute|Clinical Attribute|General Exam|3282,3287|false|false|false|C1717255||edema
Event|Event|General Exam|3282,3287|false|false|false|||edema
Finding|Pathologic Function|General Exam|3282,3287|false|false|false|C0013604|Edema|edema
Event|Event|General Exam|3302,3314|false|false|false|||distribution
Finding|Cell Function|General Exam|3302,3314|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Finding|Functional Concept|General Exam|3302,3314|false|false|false|C1704711;C5779816|Distribution;Distribution [PK]|distribution
Event|Event|General Exam|3325,3329|false|false|false|||exam
Finding|Functional Concept|General Exam|3325,3329|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|3325,3329|false|false|false|C0582103|Medical Examination|exam
Finding|Body Substance|Hospital Course|3358,3365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|3358,3365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|3358,3365|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|3366,3375|false|false|false|||presented
Event|Event|Hospital Course|3405,3415|false|false|false|||complaints
Finding|Finding|Hospital Course|3405,3415|false|false|false|C5441521|Complaint (finding)|complaints
Finding|Sign or Symptom|Hospital Course|3420,3425|false|false|false|C0033774|Pruritus|itchy
Anatomy|Body Location or Region|Hospital Course|3426,3430|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|3426,3430|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|3426,3430|false|false|false|C0362076|Problems with head|head
Event|Event|Hospital Course|3426,3430|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3426,3430|false|false|false|C0876917|Procedure on head|head
Event|Event|Hospital Course|3443,3451|false|false|false|||hardware
Event|Event|Hospital Course|3462,3470|false|false|false|||admitted
Anatomy|Anatomical Structure|Hospital Course|3478,3483|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|3489,3500|false|false|false|||observation
Finding|Finding|Hospital Course|3489,3500|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Finding|Idea or Concept|Hospital Course|3489,3500|false|false|false|C0478530;C1548358;C1554188;C5890437|Examination and observation for unspecified reason;Observation (finding)|observation
Procedure|Diagnostic Procedure|Hospital Course|3489,3500|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Health Care Activity|Hospital Course|3489,3500|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Procedure|Research Activity|Hospital Course|3489,3500|false|false|false|C0302523;C0700325;C1964257|Observation - diagnostic procedure;Observation in research;Patient observation|observation
Event|Event|Hospital Course|3519,3527|false|false|false|||planning
Finding|Functional Concept|Hospital Course|3519,3527|false|false|false|C0032074;C1301732|Planned|planning
Finding|Mental Process|Hospital Course|3519,3527|false|false|false|C0032074;C1301732|Planned|planning
Event|Event|Hospital Course|3546,3551|false|false|false|||taken
Disorder|Injury or Poisoning|Hospital Course|3566,3571|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Finding|Body Substance|Hospital Course|3566,3571|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Hospital Course|3566,3571|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Hospital Course|3566,3571|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Event|Event|Hospital Course|3572,3580|false|false|false|||revision
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3572,3580|false|false|false|C0558347;C1527075|Revision procedure;Surgical revision|revision
Event|Activity|Hospital Course|3585,3592|false|false|false|C1883720|Removing (action)|removal
Event|Event|Hospital Course|3585,3592|false|false|false|||removal
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3585,3592|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|removal
Event|Event|Hospital Course|3609,3617|false|false|false|||hardware
Event|Event|Hospital Course|3624,3633|false|false|false|||tolerated
Attribute|Clinical Attribute|Hospital Course|3638,3647|false|false|false|C0945766||procedure
Event|Event|Hospital Course|3638,3647|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|3638,3647|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|3638,3647|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3638,3647|false|false|false|C0184661|Interventional procedure|procedure
Finding|Finding|Hospital Course|3648,3652|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|3661,3672|false|false|false|||transferred
Event|Event|Hospital Course|3712,3723|false|false|false|||transferred
Anatomy|Anatomical Structure|Hospital Course|3731,3736|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|Hospital Course|3750,3760|false|false|false|||management
Event|Occupational Activity|Hospital Course|3750,3760|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|3750,3760|false|false|false|C0376636|Disease Management|management
Event|Event|Hospital Course|3774,3780|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|3774,3780|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|Hospital Course|3814,3820|false|false|false|||deemed
Event|Activity|Hospital Course|3821,3824|false|false|false|C2349186|Fit (action)|fit
Event|Event|Hospital Course|3821,3824|false|false|false|||fit
Finding|Finding|Hospital Course|3821,3824|false|false|false|C0036572;C0424576;C4553125;C5703308|Fit and well;Fit by Myeloma Frailty Index;Prosthesis fit;Seizures|fit
Finding|Sign or Symptom|Hospital Course|3821,3824|false|false|false|C0036572;C0424576;C4553125;C5703308|Fit and well;Fit by Myeloma Frailty Index;Prosthesis fit;Seizures|fit
Procedure|Laboratory Procedure|Hospital Course|3821,3824|false|false|false|C2700166|Fecal Immunochemical Test|fit
Event|Event|Hospital Course|3829,3838|false|false|false|||discharge
Finding|Body Substance|Hospital Course|3829,3838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|3829,3838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|3829,3838|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|3829,3838|false|false|false|C0030685|Patient Discharge|discharge
Attribute|Clinical Attribute|Hospital Course|3853,3865|false|false|false|C3263700||instructions
Event|Event|Hospital Course|3853,3865|false|false|false|||instructions
Finding|Intellectual Product|Hospital Course|3853,3865|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|instructions
Finding|Finding|Hospital Course|3871,3876|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|3871,3876|false|false|false|C0587267;C3810854|Close;Closed|close
Event|Event|Hospital Course|3877,3883|false|false|false|||follow
Finding|Functional Concept|Hospital Course|3877,3883|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|3877,3883|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|3877,3886|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|Hospital Course|3877,3886|false|false|false|C1522577|follow-up|follow-up
Event|Event|Hospital Course|3884,3886|false|false|false|||up
Anatomy|Body Location or Region|Hospital Course|3894,3902|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Hospital Course|3894,3902|false|false|false|C0332803|Surgical wound|incision
Event|Event|Hospital Course|3894,3902|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Hospital Course|3894,3902|false|false|false|C0184898|Surgical incisions|incision
Attribute|Clinical Attribute|Hospital Course|3908,3919|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|3908,3919|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|3908,3919|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|3908,3919|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|3908,3932|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Hospital Course|3923,3932|false|false|false|||Admission
Procedure|Health Care Activity|Hospital Course|3923,3932|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Hazardous or Poisonous Substance|Hospital Course|3934,3946|false|false|false|C0004482|azathioprine|azathioprine
Drug|Organic Chemical|Hospital Course|3934,3946|false|false|false|C0004482|azathioprine|azathioprine
Drug|Pharmacologic Substance|Hospital Course|3934,3946|false|false|false|C0004482|azathioprine|azathioprine
Event|Event|Hospital Course|3934,3946|false|false|false|||azathioprine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|3948,3955|false|false|false|C0678171|Pentasa|Pentasa
Drug|Pharmacologic Substance|Hospital Course|3948,3955|false|false|false|C0678171|Pentasa|Pentasa
Event|Event|Hospital Course|3948,3955|false|false|false|||Pentasa
Drug|Organic Chemical|Hospital Course|3957,3967|false|false|false|C0076829|topiramate|topiramate
Drug|Pharmacologic Substance|Hospital Course|3957,3967|false|false|false|C0076829|topiramate|topiramate
Event|Event|Hospital Course|3957,3967|false|false|false|||topiramate
Procedure|Laboratory Procedure|Hospital Course|3957,3967|false|false|false|C0519827|Topiramate measurement|topiramate
Drug|Organic Chemical|Hospital Course|3969,3979|false|false|false|C0002333|alprazolam|alprazolam
Drug|Pharmacologic Substance|Hospital Course|3969,3979|false|false|false|C0002333|alprazolam|alprazolam
Event|Event|Hospital Course|3969,3979|false|false|false|||alprazolam
Drug|Organic Chemical|Hospital Course|3981,3991|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|3981,3991|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|3981,3991|false|false|false|||omeprazole
Drug|Organic Chemical|Hospital Course|3993,4001|false|false|false|C0078839|zolpidem|zolpidem
Drug|Pharmacologic Substance|Hospital Course|3993,4001|false|false|false|C0078839|zolpidem|zolpidem
Event|Event|Hospital Course|3993,4001|false|false|false|||zolpidem
Drug|Organic Chemical|Hospital Course|4003,4014|false|false|false|C0078569|venlafaxine|venlafaxine
Drug|Pharmacologic Substance|Hospital Course|4003,4014|false|false|false|C0078569|venlafaxine|venlafaxine
Event|Event|Hospital Course|4003,4014|false|false|false|||venlafaxine
Drug|Organic Chemical|Hospital Course|4003,4018|false|false|false|C0771200|venlafaxine hydrochloride|venlafaxine hcl
Drug|Pharmacologic Substance|Hospital Course|4003,4018|false|false|false|C0771200|venlafaxine hydrochloride|venlafaxine hcl
Drug|Organic Chemical|Hospital Course|4003,4021|false|false|false|C2918046|Venlafaxine Hydrochloride ER|venlafaxine hcl er
Drug|Pharmacologic Substance|Hospital Course|4003,4021|false|false|false|C2918046|Venlafaxine Hydrochloride ER|venlafaxine hcl er
Disorder|Neoplastic Process|Hospital Course|4015,4018|false|false|false|C0023443|Hairy Cell Leukemia|hcl
Drug|Immunologic Factor|Hospital Course|4015,4018|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|hcl
Drug|Inorganic Chemical|Hospital Course|4015,4018|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|hcl
Drug|Pharmacologic Substance|Hospital Course|4015,4018|false|false|false|C0443985;C1512523|Flinders medical centre-7 marker;hydrochloride|hcl
Event|Event|Hospital Course|4015,4018|false|false|false|||hcl
Event|Event|Hospital Course|4026,4041|false|false|false|||popylthiouracil
Drug|Organic Chemical|Hospital Course|4043,4055|false|false|false|C0033405|promethazine|promethazine
Drug|Pharmacologic Substance|Hospital Course|4043,4055|false|false|false|C0033405|promethazine|promethazine
Event|Event|Hospital Course|4043,4055|false|false|false|||promethazine
Finding|Body Substance|Hospital Course|4057,4064|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|4057,4064|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|4057,4064|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|Hospital Course|4079,4084|false|false|false|||doses
Finding|Finding|Hospital Course|4093,4097|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|4093,4097|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|4093,4097|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Hospital Course|4105,4109|false|false|false|||exam
Finding|Functional Concept|Hospital Course|4105,4109|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|4105,4109|false|false|false|C0582103|Medical Examination|exam
Event|Event|Hospital Course|4114,4123|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|4114,4123|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|4114,4123|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|4114,4123|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|4114,4123|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|4114,4135|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|4124,4135|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|4124,4135|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|4124,4135|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|4124,4135|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|4140,4153|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|4140,4153|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|4140,4153|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|4140,4153|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|4161,4167|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|4177,4184|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|Hospital Course|4177,4184|false|false|false|||Tablets
Event|Event|Hospital Course|4212,4218|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|4223,4227|false|false|false|C2598155||pain
Event|Event|Hospital Course|4223,4227|false|false|false|||pain
Finding|Functional Concept|Hospital Course|4223,4227|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|4223,4227|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Hospital Course|4234,4246|false|false|false|C0004482|azathioprine|azathioprine
Drug|Organic Chemical|Hospital Course|4234,4246|false|false|false|C0004482|azathioprine|azathioprine
Drug|Pharmacologic Substance|Hospital Course|4234,4246|false|false|false|C0004482|azathioprine|azathioprine
Event|Event|Hospital Course|4234,4246|false|false|false|||azathioprine
Drug|Biomedical or Dental Material|Hospital Course|4253,4259|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|4273,4279|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|4273,4279|false|false|false|||Tablet
Drug|Organic Chemical|Hospital Course|4304,4314|false|false|false|C0002333|alprazolam|alprazolam
Drug|Pharmacologic Substance|Hospital Course|4304,4314|false|false|false|C0002333|alprazolam|alprazolam
Event|Event|Hospital Course|4304,4314|false|false|false|||alprazolam
Drug|Biomedical or Dental Material|Hospital Course|4320,4326|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|4327,4330|false|false|false|||Sig
Drug|Biomedical or Dental Material|Hospital Course|4336,4342|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|4346,4349|false|false|false|||TID
Finding|Finding|Hospital Course|4351,4358|false|false|false|C4035626|3 times|3 times
Disorder|Disease or Syndrome|Hospital Course|4353,4358|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|4353,4358|false|false|false|||times
Finding|Idea or Concept|Hospital Course|4361,4364|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4361,4364|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|4370,4376|false|false|false|||needed
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4381,4388|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|4381,4388|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|4381,4388|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Organic Chemical|Hospital Course|4395,4407|false|false|false|C0033405|promethazine|promethazine
Drug|Pharmacologic Substance|Hospital Course|4395,4407|false|false|false|C0033405|promethazine|promethazine
Event|Event|Hospital Course|4395,4407|false|false|false|||promethazine
Drug|Biomedical or Dental Material|Hospital Course|4414,4420|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|4434,4440|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|4434,4440|false|false|false|||Tablet
Event|Event|Hospital Course|4468,4474|false|false|false|||needed
Attribute|Clinical Attribute|Hospital Course|4479,4485|false|false|false|C4255480||nausea
Event|Event|Hospital Course|4479,4485|false|false|false|||nausea
Finding|Sign or Symptom|Hospital Course|4479,4485|false|false|false|C0027497|Nausea|nausea
Drug|Organic Chemical|Hospital Course|4492,4502|false|false|false|C0028978|omeprazole|omeprazole
Drug|Pharmacologic Substance|Hospital Course|4492,4502|false|false|false|C0028978|omeprazole|omeprazole
Event|Event|Hospital Course|4492,4502|false|false|false|||omeprazole
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4509,4516|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4509,4516|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4509,4516|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|4518,4525|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|4518,4533|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|4526,4533|false|false|false|||Release
Finding|Functional Concept|Hospital Course|4526,4533|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|4526,4533|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4526,4533|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Event|Event|Hospital Course|4540,4543|false|false|false|||Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4554,4561|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4554,4561|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4554,4561|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Attribute|Clinical Attribute|Hospital Course|4563,4570|false|false|false|C1545665|Views delayed|Delayed
Drug|Biomedical or Dental Material|Hospital Course|4563,4578|false|false|false|C1707664|Delayed Release Dosage Form|Delayed Release
Event|Event|Hospital Course|4571,4578|false|false|false|||Release
Finding|Functional Concept|Hospital Course|4571,4578|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|4571,4578|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4571,4578|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Antibiotic|Hospital Course|4608,4618|false|false|false|C0007716|cephalexin|cephalexin
Drug|Organic Chemical|Hospital Course|4608,4618|false|false|false|C0007716|cephalexin|cephalexin
Event|Event|Hospital Course|4608,4618|false|false|false|||cephalexin
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4626,4633|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4626,4633|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4626,4633|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4647,4654|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4647,4654|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4647,4654|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Intellectual Product|Hospital Course|4663,4668|false|false|false|C1720374|Every - dosing instruction fragment|every
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4701,4708|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4701,4708|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4701,4708|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Finding|Idea or Concept|Hospital Course|4713,4720|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|4728,4736|false|false|false|C1692318|docusate|docusate
Drug|Pharmacologic Substance|Hospital Course|4728,4736|false|false|false|C1692318|docusate|docusate
Event|Event|Hospital Course|4728,4736|false|false|false|||docusate
Drug|Organic Chemical|Hospital Course|4728,4743|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Pharmacologic Substance|Hospital Course|4728,4743|false|false|false|C0243237|docusate sodium|docusate sodium
Drug|Biologically Active Substance|Hospital Course|4737,4743|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Element, Ion, or Isotope|Hospital Course|4737,4743|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Drug|Pharmacologic Substance|Hospital Course|4737,4743|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|sodium
Event|Event|Hospital Course|4737,4743|false|false|false|||sodium
Finding|Physiologic Function|Hospital Course|4737,4743|false|false|false|C4553025|Sodium metabolic function|sodium
Procedure|Laboratory Procedure|Hospital Course|4737,4743|false|false|false|C0337443|Sodium measurement|sodium
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4751,4758|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4751,4758|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4751,4758|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4772,4779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4772,4779|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4772,4779|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Disorder|Mental or Behavioral Dysfunction|Hospital Course|4783,4786|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|4783,4786|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|4783,4786|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|4783,4786|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|4783,4786|false|false|false|C1332410|BID gene|BID
Disorder|Disease or Syndrome|Hospital Course|4791,4796|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|4799,4802|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|4799,4802|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|4810,4818|false|false|false|C0078839|zolpidem|zolpidem
Drug|Pharmacologic Substance|Hospital Course|4810,4818|false|false|false|C0078839|zolpidem|zolpidem
Drug|Biomedical or Dental Material|Hospital Course|4824,4830|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|4844,4850|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|4844,4850|false|false|false|||Tablet
Event|Event|Hospital Course|4874,4880|false|false|false|||needed
Drug|Organic Chemical|Hospital Course|4889,4894|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|4889,4894|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Event|Event|Hospital Course|4889,4894|false|false|false|||sleep
Finding|Organism Function|Hospital Course|4889,4894|false|false|false|C0037313|Sleep|sleep
Drug|Organic Chemical|Hospital Course|4901,4911|false|false|false|C0127615|mesalamine|mesalamine
Drug|Pharmacologic Substance|Hospital Course|4901,4911|false|false|false|C0127615|mesalamine|mesalamine
Event|Event|Hospital Course|4901,4911|false|false|false|||mesalamine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4919,4926|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4919,4926|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4919,4926|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4919,4944|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Hospital Course|4928,4936|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|4928,4936|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|4937,4944|false|false|false|||Release
Finding|Functional Concept|Hospital Course|4937,4944|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|4937,4944|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4937,4944|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|4959,4966|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|4959,4966|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4959,4966|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|4959,4984|false|false|false|C0991505|Extended Release Oral Capsule|Capsule, Extended Release
Finding|Finding|Hospital Course|4968,4976|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|4968,4976|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|4977,4984|false|false|false|||Release
Finding|Functional Concept|Hospital Course|4977,4984|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|4977,4984|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|4977,4984|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Finding|Hospital Course|4993,5000|false|false|false|C4264481|4 times|4 times
Disorder|Disease or Syndrome|Hospital Course|4995,5000|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5003,5006|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5003,5006|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5015,5025|false|false|false|C0076829|topiramate|topiramate
Drug|Pharmacologic Substance|Hospital Course|5015,5025|false|false|false|C0076829|topiramate|topiramate
Event|Event|Hospital Course|5015,5025|false|false|false|||topiramate
Procedure|Laboratory Procedure|Hospital Course|5015,5025|false|false|false|C0519827|Topiramate measurement|topiramate
Drug|Biomedical or Dental Material|Hospital Course|5033,5039|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5053,5059|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|5060,5062|false|false|false|||PO
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5063,5066|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5063,5066|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5063,5066|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5063,5066|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5063,5066|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5068,5075|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|5070,5075|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|Hospital Course|5070,5075|false|false|false|||times
Finding|Idea or Concept|Hospital Course|5079,5082|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5079,5082|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|5091,5102|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5091,5102|false|false|false|C0082607|fluticasone|fluticasone
Drug|Pharmacologic Substance|Hospital Course|5091,5113|false|false|false|C0939232|fluticasone / salmeterol|fluticasone-salmeterol
Drug|Organic Chemical|Hospital Course|5103,5113|false|false|false|C0073992|salmeterol|salmeterol
Drug|Pharmacologic Substance|Hospital Course|5103,5113|false|false|false|C0073992|salmeterol|salmeterol
Event|Event|Hospital Course|5103,5113|false|false|false|||salmeterol
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5130,5134|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5130,5134|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5140,5146|false|false|false|C1550509|Participation Type - device|Device
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5147,5150|false|false|false|C0262329|Short insular gyrus|Sig
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5147,5150|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Drug|Immunologic Factor|Hospital Course|5147,5150|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Finding|Receptor|Hospital Course|5147,5150|false|false|false|C0034789|Receptors, Antigen, B-Cell|Sig
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5161,5165|false|false|false|C1556138|Disc - Body Part|Disk
Drug|Biomedical or Dental Material|Hospital Course|5161,5165|false|false|false|C0993608|Disk Drug Form|Disk
Finding|Functional Concept|Hospital Course|5171,5177|false|false|false|C1550509|Participation Type - device|Device
Event|Event|Hospital Course|5178,5188|false|false|false|||Inhalation
Finding|Functional Concept|Hospital Course|5178,5188|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Finding|Organism Function|Hospital Course|5178,5188|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|Inhalation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5189,5192|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5189,5192|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|5189,5192|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|5189,5192|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|5189,5192|false|false|false|C1332410|BID gene|BID
Finding|Finding|Hospital Course|5194,5201|false|false|false|C4035627|2 times|2 times
Disorder|Disease or Syndrome|Hospital Course|5196,5201|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Finding|Idea or Concept|Hospital Course|5204,5207|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5204,5207|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Hospital Course|5216,5232|false|false|false|C0033511|propylthiouracil|propylthiouracil
Drug|Pharmacologic Substance|Hospital Course|5216,5232|false|false|false|C0033511|propylthiouracil|propylthiouracil
Event|Event|Hospital Course|5216,5232|false|false|false|||propylthiouracil
Drug|Biomedical or Dental Material|Hospital Course|5239,5245|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5259,5265|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Organic Chemical|Hospital Course|5297,5308|false|false|false|C0078569|venlafaxine|venlafaxine
Drug|Pharmacologic Substance|Hospital Course|5297,5308|false|false|false|C0078569|venlafaxine|venlafaxine
Event|Event|Hospital Course|5297,5308|false|false|false|||venlafaxine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5315,5322|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5315,5322|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5315,5322|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5315,5341|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Hospital Course|5324,5327|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Hospital Course|5324,5327|false|false|false|||Ext
Finding|Gene or Genome|Hospital Course|5324,5327|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Hospital Course|5328,5335|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5328,5335|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5328,5335|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5328,5335|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5356,5363|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5356,5363|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5356,5363|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5356,5382|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Hospital Course|5365,5368|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Hospital Course|5365,5368|false|false|false|||Ext
Finding|Gene or Genome|Hospital Course|5365,5368|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Hospital Course|5369,5376|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5369,5376|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5369,5376|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5369,5376|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|5407,5418|false|false|false|C0078569|venlafaxine|venlafaxine
Drug|Pharmacologic Substance|Hospital Course|5407,5418|false|false|false|C0078569|venlafaxine|venlafaxine
Event|Event|Hospital Course|5407,5418|false|false|false|||venlafaxine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5425,5432|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5425,5432|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5425,5432|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5425,5451|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Hospital Course|5434,5437|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Hospital Course|5434,5437|false|false|false|||Ext
Finding|Gene or Genome|Hospital Course|5434,5437|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Hospital Course|5438,5445|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5438,5445|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5438,5445|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5438,5445|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5466,5473|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Anatomy|Cell Component|Hospital Course|5466,5473|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5466,5473|false|false|false|C0006935|capsule (pharmacologic)|Capsule
Drug|Biomedical or Dental Material|Hospital Course|5466,5492|false|false|false|C1337463|CAPSULE, EXT RELEASE 24 HR|Capsule, Ext Release 24 hr
Disorder|Congenital Abnormality|Hospital Course|5475,5478|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|Hospital Course|5475,5478|false|false|false|||Ext
Finding|Gene or Genome|Hospital Course|5475,5478|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|Hospital Course|5479,5486|false|false|false|||Release
Finding|Functional Concept|Hospital Course|5479,5486|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|5479,5486|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5479,5486|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|5517,5528|false|false|false|C0020264|hydrocodone|hydrocodone
Drug|Pharmacologic Substance|Hospital Course|5517,5528|false|false|false|C0020264|hydrocodone|hydrocodone
Drug|Organic Chemical|Hospital Course|5529,5542|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|5529,5542|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|5529,5542|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|5529,5542|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|5550,5556|false|false|false|C0039225|Tablet Dosage Form|Tablet
Drug|Biomedical or Dental Material|Hospital Course|5566,5573|false|false|false|C0039225|Tablet Dosage Form|Tablets
Event|Event|Hospital Course|5566,5573|false|false|false|||Tablets
Event|Event|Hospital Course|5601,5607|false|false|false|||needed
Finding|Sign or Symptom|Hospital Course|5612,5621|false|true|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|Hospital Course|5617,5621|false|false|false|C2598155||pain
Event|Event|Hospital Course|5617,5621|false|false|false|||pain
Finding|Functional Concept|Hospital Course|5617,5621|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|5617,5621|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Biomedical or Dental Material|Hospital Course|5632,5638|false|false|false|C0039225|Tablet Dosage Form|Tablet
Finding|Idea or Concept|Hospital Course|5643,5650|false|false|false|C0807726|refill|Refills
Event|Event|Hospital Course|5658,5667|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5658,5667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5658,5667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5658,5667|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5658,5667|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|5658,5679|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|5658,5679|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|5668,5679|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|5668,5679|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|5668,5679|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|5681,5685|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|5681,5685|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|5681,5685|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|5681,5685|false|false|false|C1553498|home health encounter|Home
Event|Event|Hospital Course|5688,5697|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|5688,5697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|5688,5697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|5688,5697|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|5688,5697|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|5688,5707|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|5698,5707|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|5698,5707|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|5698,5707|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|5698,5707|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|5698,5707|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Injury or Poisoning|Hospital Course|5709,5717|false|false|false|C0274281|Injury due to exposure to external cause|exposure
Event|Event|Hospital Course|5709,5717|false|false|false|||exposure
Finding|Finding|Hospital Course|5709,5717|false|false|false|C2220266|exposure history|exposure
Phenomenon|Phenomenon or Process|Hospital Course|5709,5717|false|false|false|C0728853|Accident due to exposure to weather conditions|exposure
Event|Event|Hospital Course|5721,5731|false|false|false|||craniotomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5721,5731|false|false|false|C0010280|Craniotomy|craniotomy
Event|Event|Hospital Course|5732,5740|false|false|false|||hardware
Disorder|Disease or Syndrome|Hospital Course|5745,5754|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Hospital Course|5745,5754|false|false|false|||infection
Finding|Pathologic Function|Hospital Course|5745,5754|false|false|false|C3714514|Infection|infection
Finding|Mental Process|Discharge Condition|5779,5785|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|5779,5792|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|5779,5792|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|5786,5792|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|5786,5792|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|5794,5799|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|5794,5799|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|5804,5812|false|false|false|||coherent
Finding|Finding|Discharge Condition|5804,5812|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|5814,5819|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|5814,5836|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|5814,5836|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|5823,5836|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|5823,5836|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|5823,5836|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|5838,5843|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|5838,5843|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|5838,5843|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|5838,5843|false|false|false|||Alert
Finding|Finding|Discharge Condition|5838,5843|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|5838,5843|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|5838,5843|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|5848,5859|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|5848,5859|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|5861,5869|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|5861,5869|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|5861,5869|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|5870,5876|false|false|false|C5889824||Status
Event|Event|Discharge Condition|5870,5876|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|5870,5876|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|5878,5888|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|5878,5888|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|5878,5888|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|5878,5888|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|5878,5888|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|5891,5902|false|false|false|||Independent
Finding|Finding|Discharge Condition|5891,5902|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|5891,5902|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Event|Event|Discharge Instructions|5939,5945|false|false|false|||friend
Finding|Idea or Concept|Discharge Instructions|5939,5945|false|false|false|C1546502|Relationship - Friend|friend
Finding|Classification|Discharge Instructions|5946,5952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|5946,5952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|5946,5952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|5946,5952|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Discharge Instructions|5960,5965|false|false|false|||check
Anatomy|Body Location or Region|Discharge Instructions|5971,5979|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5971,5979|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5971,5979|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5971,5979|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5991,5996|false|false|false|||signs
Finding|Finding|Discharge Instructions|5991,5996|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|5991,5996|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|6000,6009|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|6000,6009|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|6000,6009|false|false|false|C3714514|Infection|infection
Event|Event|Discharge Instructions|6012,6016|false|false|false|||Take
Attribute|Clinical Attribute|Discharge Instructions|6022,6026|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6022,6026|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6022,6026|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6022,6026|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|6022,6035|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|6022,6035|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|6022,6035|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|6027,6035|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6027,6035|false|false|false|||medicine
Event|Event|Discharge Instructions|6039,6049|false|false|false|||prescribed
Event|Event|Discharge Instructions|6052,6060|false|false|false|||Exercise
Finding|Daily or Recreational Activity|Discharge Instructions|6052,6060|false|false|false|C0015259|Exercise|Exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6052,6060|false|false|false|C1522704|Exercise Pain Management|Exercise
Event|Event|Discharge Instructions|6071,6078|false|false|false|||limited
Event|Event|Discharge Instructions|6082,6089|false|false|false|||walking
Finding|Daily or Recreational Activity|Discharge Instructions|6082,6089|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Finding|Discharge Instructions|6082,6089|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Finding|Sign or Symptom|Discharge Instructions|6082,6089|false|true|false|C0080331;C2346415;C2368355|Walking (function);history of recreational walking;walking - neurological symptom|walking
Event|Activity|Discharge Instructions|6094,6101|true|false|false|C0206244|Lifting|lifting
Event|Event|Discharge Instructions|6094,6101|false|false|false|||lifting
Event|Event|Discharge Instructions|6103,6112|false|false|false|||straining
Finding|Physiologic Function|Discharge Instructions|6103,6112|true|false|false|C0442694|Straining (finding)|straining
Disorder|Disease or Syndrome|Discharge Instructions|6128,6135|false|false|false|C0011119|Decompression Sickness|bending
Event|Event|Discharge Instructions|6128,6135|false|false|false|||bending
Finding|Finding|Discharge Instructions|6128,6135|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Finding|Physiologic Function|Discharge Instructions|6128,6135|false|false|false|C0700231;C2584296|Bending - Changing basic body position;Does bend|bending
Event|Event|Discharge Instructions|6146,6150|false|false|false|||wash
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6156,6160|false|false|false|C0018494|Hair|hair
Finding|Body Substance|Discharge Instructions|6156,6160|false|false|false|C0444095;C1546660|Hair Specimen;Hair Specimen Code|hair
Finding|Intellectual Product|Discharge Instructions|6156,6160|false|false|false|C0444095;C1546660|Hair Specimen;Hair Specimen Code|hair
Anatomy|Body Space or Junction|Discharge Instructions|6172,6179|false|false|false|C0502420|Suture Joint|sutures
Event|Event|Discharge Instructions|6206,6213|false|false|false|||removed
Event|Event|Discharge Instructions|6217,6225|false|false|false|||Increase
Event|Event|Discharge Instructions|6231,6237|false|false|false|||intake
Finding|Functional Concept|Discharge Instructions|6231,6237|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Discharge Instructions|6231,6237|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Drug|Substance|Discharge Instructions|6241,6247|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|6241,6247|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|6241,6247|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6241,6247|false|false|false|C0016286|Fluid Therapy|fluids
Anatomy|Tissue|Discharge Instructions|6252,6257|false|false|false|C1304649|Tissue fiber|fiber
Drug|Organic Chemical|Discharge Instructions|6252,6257|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Pharmacologic Substance|Discharge Instructions|6252,6257|false|false|false|C0225326;C1321801|Fiber brand of calcium polycarbophil;fiber|fiber
Drug|Hazardous or Poisonous Substance|Discharge Instructions|6262,6270|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|6262,6270|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|6271,6275|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6271,6275|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6271,6275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6271,6275|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|6277,6285|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6277,6285|false|false|false|||medicine
Event|Event|Discharge Instructions|6290,6295|false|false|false|||cause
Event|Event|Discharge Instructions|6296,6308|false|false|false|||constipation
Finding|Sign or Symptom|Discharge Instructions|6296,6308|false|false|false|C0009806|Constipation|constipation
Event|Event|Discharge Instructions|6323,6332|false|false|false|||recommend
Event|Event|Discharge Instructions|6333,6339|false|false|false|||taking
Drug|Pharmacologic Substance|Discharge Instructions|6344,6360|false|false|false|C0013231|Drugs, Non-Prescription|over the counter
Drug|Hazardous or Poisonous Substance|Discharge Instructions|6353,6360|false|false|false|C0702263|Counter brand of Terbufos|counter
Drug|Organic Chemical|Discharge Instructions|6353,6360|false|false|false|C0702263|Counter brand of Terbufos|counter
Finding|Body Substance|Discharge Instructions|6361,6366|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|6361,6375|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|6361,6375|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|6367,6375|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|6385,6393|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Discharge Instructions|6385,6393|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Discharge Instructions|6395,6401|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|6395,6401|false|false|false|C0282139|Colace|Colace
Drug|Hazardous or Poisonous Substance|Discharge Instructions|6417,6425|false|false|false|C0027415|Narcotics|narcotic
Drug|Pharmacologic Substance|Discharge Instructions|6417,6425|false|false|false|C0027415|Narcotics|narcotic
Attribute|Clinical Attribute|Discharge Instructions|6426,6430|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6426,6430|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6426,6430|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6426,6430|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|6431,6441|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|6431,6441|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|6431,6441|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|6451,6459|false|false|false|||directed
Event|Event|Discharge Instructions|6468,6474|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|6468,6474|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|6483,6487|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|6493,6510|false|false|false|C0003209|Anti-Inflammatory Agents|anti-inflammatory
Drug|Pharmacologic Substance|Discharge Instructions|6511,6520|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|6511,6520|false|false|false|||medicines
Drug|Organic Chemical|Discharge Instructions|6529,6535|false|false|false|C0699203|Motrin|Motrin
Drug|Pharmacologic Substance|Discharge Instructions|6529,6535|false|false|false|C0699203|Motrin|Motrin
Drug|Organic Chemical|Discharge Instructions|6537,6544|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Discharge Instructions|6537,6544|false|false|false|C0004057|aspirin|Aspirin
Event|Event|Discharge Instructions|6537,6544|false|false|false|||Aspirin
Drug|Organic Chemical|Discharge Instructions|6546,6551|false|false|false|C0593507|Advil|Advil
Drug|Pharmacologic Substance|Discharge Instructions|6546,6551|false|false|false|C0593507|Advil|Advil
Event|Event|Discharge Instructions|6546,6551|false|false|false|||Advil
Finding|Gene or Genome|Discharge Instructions|6546,6551|false|false|false|C1422473|AVIL gene|Advil
Drug|Organic Chemical|Discharge Instructions|6558,6567|false|false|false|C0020740|ibuprofen|Ibuprofen
Drug|Pharmacologic Substance|Discharge Instructions|6558,6567|false|false|false|C0020740|ibuprofen|Ibuprofen
Finding|Idea or Concept|Discharge Instructions|6568,6571|false|false|false|C1548556|Etc.|etc
Event|Event|Discharge Instructions|6574,6575|false|false|false|||
Attribute|Clinical Attribute|Discharge Instructions|6575,6584|false|false|false|C1382187|Clearance of substance|Clearance
Event|Event|Discharge Instructions|6575,6584|false|false|false|||Clearance
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|6575,6584|false|false|false|C2825073|Clearance [PK]|Clearance
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6575,6584|false|false|false|C4554548|Clearance procedure|Clearance
Event|Event|Discharge Instructions|6588,6593|false|false|false|||drive
Event|Event|Discharge Instructions|6598,6604|false|false|false|||return
Event|Occupational Activity|Discharge Instructions|6608,6612|false|false|false|C0043227|Work|work
Event|Event|Discharge Instructions|6621,6630|false|false|false|||addressed
Finding|Idea or Concept|Discharge Instructions|6655,6661|false|false|false|C1549636|Address type - Office|office
Procedure|Health Care Activity|Discharge Instructions|6655,6667|false|false|false|C0028900|Office Visits|office visit
Event|Event|Discharge Instructions|6662,6667|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|6662,6667|false|false|false|C0545082|Visit|visit
Event|Event|Discharge Instructions|6670,6674|false|false|false|||Make
Finding|Functional Concept|Discharge Instructions|6670,6674|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Finding|Intellectual Product|Discharge Instructions|6670,6674|false|false|false|C0947322;C1881534|Make - Instruction Imperative;Manufacturer Name|Make
Event|Event|Discharge Instructions|6675,6679|false|false|false|||sure
Finding|Intellectual Product|Discharge Instructions|6675,6679|false|false|false|C4724437|SURE Test|sure
Event|Event|Discharge Instructions|6683,6691|false|false|false|||continue
Finding|Idea or Concept|Discharge Instructions|6683,6691|false|false|false|C0549178|Continuous|continue
Event|Event|Discharge Instructions|6695,6698|false|false|false|||use
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6704,6724|false|false|false|C0454512|Incentive spirometry|incentive spirometer
Finding|Finding|Discharge Instructions|6732,6739|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|6735,6739|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|6735,6739|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|6735,6739|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|6762,6772|false|false|false|||instructed
Event|Event|Discharge Instructions|6783,6787|false|false|false|||CALL
Finding|Functional Concept|Discharge Instructions|6783,6787|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Gene or Genome|Discharge Instructions|6783,6787|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Intellectual Product|Discharge Instructions|6783,6787|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Finding|Mental Process|Discharge Instructions|6783,6787|false|false|false|C0679006;C1413393;C1720420;C1947967|CHL1 gene;Call (Instruction);Call - dosing instruction fragment;Decision|CALL
Attribute|Clinical Attribute|Discharge Instructions|6793,6800|false|false|false|C5444295||SURGEON
Event|Event|Discharge Instructions|6793,6800|false|false|false|||SURGEON
Event|Event|Discharge Instructions|6820,6830|false|false|false|||EXPERIENCE
Finding|Mental Process|Discharge Instructions|6820,6830|false|false|false|C0237607;C0596545|Experience;Experience (Practice)|EXPERIENCE
Event|Event|Discharge Instructions|6831,6834|false|false|false|||ANY
Finding|Finding|Discharge Instructions|6855,6858|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Idea or Concept|Discharge Instructions|6855,6858|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|New
Finding|Finding|Discharge Instructions|6855,6864|false|false|false|C0746890|new onset|New onset
Event|Event|Discharge Instructions|6859,6864|false|false|false|||onset
Event|Event|Discharge Instructions|6868,6875|false|false|false|||tremors
Finding|Sign or Symptom|Discharge Instructions|6868,6875|false|false|false|C0040822|Tremor|tremors
Event|Event|Discharge Instructions|6879,6887|false|false|false|||seizures
Finding|Sign or Symptom|Discharge Instructions|6879,6887|false|false|false|C0036572|Seizures|seizures
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|6894,6903|true|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|6894,6903|false|false|false|||confusion
Finding|Finding|Discharge Instructions|6894,6903|true|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Discharge Instructions|6907,6913|false|false|false|||change
Finding|Functional Concept|Discharge Instructions|6907,6913|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6907,6913|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|6907,6916|false|false|false|C0392747|Changing|change in
Attribute|Clinical Attribute|Discharge Instructions|6907,6930|false|false|false|C5774124||change in mental status
Finding|Finding|Discharge Instructions|6907,6930|false|false|false|C0856054|Mental status changes|change in mental status
Finding|Mental Process|Discharge Instructions|6917,6923|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Discharge Instructions|6917,6930|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Discharge Instructions|6917,6930|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Discharge Instructions|6924,6930|false|false|false|C5889824||status
Event|Event|Discharge Instructions|6924,6930|false|false|false|||status
Finding|Idea or Concept|Discharge Instructions|6924,6930|false|false|false|C1546481|What subject filter - Status|status
Event|Event|Discharge Instructions|6938,6946|false|false|false|||numbness
Finding|Finding|Discharge Instructions|6938,6946|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Discharge Instructions|6938,6946|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|Discharge Instructions|6948,6956|false|false|false|C0030554|Paresthesia|tingling
Event|Event|Discharge Instructions|6948,6956|false|false|false|||tingling
Finding|Sign or Symptom|Discharge Instructions|6948,6956|false|false|false|C2242996|Has tingling sensation|tingling
Event|Event|Discharge Instructions|6958,6966|false|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|6958,6966|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6975,6986|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Attribute|Clinical Attribute|Discharge Instructions|6989,6993|false|false|false|C2598155||Pain
Event|Event|Discharge Instructions|6989,6993|false|false|false|||Pain
Finding|Functional Concept|Discharge Instructions|6989,6993|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Discharge Instructions|6989,6993|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Event|Event|Discharge Instructions|6997,7005|false|false|false|||headache
Finding|Sign or Symptom|Discharge Instructions|6997,7005|false|false|false|C0018681|Headache|headache
Event|Event|Discharge Instructions|7026,7036|false|false|false|||increasing
Event|Event|Discharge Instructions|7046,7054|false|false|false|||relieved
Attribute|Clinical Attribute|Discharge Instructions|7058,7062|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|7058,7062|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7058,7062|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|7063,7073|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Discharge Instructions|7063,7073|false|false|false|||medication
Finding|Intellectual Product|Discharge Instructions|7063,7073|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Discharge Instructions|7080,7085|false|false|false|||signs
Finding|Finding|Discharge Instructions|7080,7085|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Discharge Instructions|7080,7085|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|Discharge Instructions|7089,7098|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|7089,7098|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|7089,7098|false|false|false|C3714514|Infection|infection
Disorder|Injury or Poisoning|Discharge Instructions|7106,7111|false|false|false|C0043250;C0043251;C3263723|Traumatic Wound;Traumatic injury;Wounds and Injuries|wound
Event|Event|Discharge Instructions|7106,7111|false|false|false|||wound
Finding|Body Substance|Discharge Instructions|7106,7111|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Functional Concept|Discharge Instructions|7106,7111|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Finding|Intellectual Product|Discharge Instructions|7106,7111|false|false|false|C1547965;C1549529;C1550680|Route of Administration - Wound;Specimen Type - Wound|wound
Anatomy|Body Location or Region|Discharge Instructions|7112,7116|false|false|false|C1515974|Anatomic Site|site
Finding|Intellectual Product|Discharge Instructions|7112,7116|false|false|false|C1546778||site
Disorder|Disease or Syndrome|Discharge Instructions|7118,7125|false|false|false|C0041834|Erythema|redness
Event|Event|Discharge Instructions|7118,7125|false|false|false|||redness
Finding|Finding|Discharge Instructions|7118,7125|false|false|false|C0332575|Redness|redness
Event|Event|Discharge Instructions|7127,7135|false|false|false|||swelling
Finding|Finding|Discharge Instructions|7127,7135|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|7127,7135|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|Discharge Instructions|7138,7148|false|false|false|||tenderness
Finding|Mental Process|Discharge Instructions|7138,7148|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|Discharge Instructions|7138,7148|false|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|Discharge Instructions|7153,7161|false|false|false|||drainage
Finding|Body Substance|Discharge Instructions|7153,7161|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|Discharge Instructions|7153,7161|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7153,7161|false|false|false|C0013103|Drainage procedure|drainage
Finding|Finding|Discharge Instructions|7164,7169|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Finding|Sign or Symptom|Discharge Instructions|7164,7169|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|Fever
Event|Event|Discharge Instructions|7186,7191|false|false|false|||equal
Finding|Intellectual Product|Discharge Instructions|7186,7191|false|false|false|C1549782|Relational Operator - Equal|equal
Procedure|Health Care Activity|Discharge Instructions|7206,7214|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|7215,7227|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|7215,7227|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|7215,7227|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

