 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|153,161|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|185,194|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|185,194|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|197,219|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|205,209|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|205,209|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|205,219|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|222,231|false|false|false|C1999232|Attending (action)|Attending
Attribute|Clinical Attribute|Chief Complaint|257,267|false|false|false|C2979880||subjective
Finding|Finding|Chief Complaint|257,267|false|false|false|C2266644|subjective (symptom)|subjective
Finding|Sign or Symptom|Chief Complaint|268,274|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|Chief Complaint|276,284|false|false|false|C0023380|Lethargy|lethargy
Finding|Finding|Chief Complaint|290,296|false|false|false|C4554530|Bloody|bloody
Drug|Substance|Chief Complaint|297,302|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Chief Complaint|297,302|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Conceptual Entity|Chief Complaint|303,309|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Chief Complaint|303,309|false|false|false|C3251815|Measurement of fluid output|output
Finding|Classification|Chief Complaint|313,318|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|319,327|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|319,327|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|331,349|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|340,349|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|340,349|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|340,349|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|340,349|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Gene or Genome|Chief Complaint|364,369|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Anatomy|Body Part, Organ, or Organ Component|Chief Complaint|370,376|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|Chief Complaint|377,382|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Chief Complaint|377,382|false|false|false|C1546638|Fluid Specimen Code|fluid
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|407,420|false|false|false|C0556030|Repositioning (procedure)|repositioning
Drug|Substance|Chief Complaint|433,438|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Chief Complaint|433,438|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Health Care Activity|Chief Complaint|443,452|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|443,452|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|Chief Complaint|459,469|false|false|false|C1524062|Additional|additional
Drug|Substance|Chief Complaint|471,476|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Chief Complaint|471,476|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|Chief Complaint|484,491|false|false|false|C1883720|Removing (action)|Removal
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|484,491|false|false|false|C0015252;C0185115;C0728940|Excision;Extraction;removal technique|Removal
Drug|Substance|Chief Complaint|516,521|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Chief Complaint|516,521|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Finding|History of Present Illness|578,581|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|PMH
Disorder|Disease or Syndrome|History of Present Illness|585,597|false|false|false|C0020538|Hypertensive disease|hypertension
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|602,609|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|602,609|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|602,609|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|History of Present Illness|611,617|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Finding|History of Present Illness|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|History of Present Illness|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|History of Present Illness|619,623|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|History of Present Illness|619,629|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|History of Present Illness|619,629|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|History of Present Illness|624,629|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|History of Present Illness|624,629|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|History of Present Illness|630,659|false|false|false|C1512751|Invasive Urothelial Carcinoma|invasive urothelial carcinoma
Disorder|Neoplastic Process|History of Present Illness|639,659|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|History of Present Illness|650,659|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Finding|History of Present Illness|660,664|false|false|false|C1711132|pT2b TNM Finding|pT2b
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|671,674|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|671,678|false|false|false|C0542407|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|TAH/BSO
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|History of Present Illness|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|History of Present Illness|675,678|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Chemical Viewed Structurally|History of Present Illness|680,687|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|680,698|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|688,698|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|701,706|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|History of Present Illness|701,714|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|701,714|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Finding|Functional Concept|History of Present Illness|719,734|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|History of Present Illness|736,745|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|History of Present Illness|736,745|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|750,756|false|false|false|C0030797|Pelvis|pelvic
Disorder|Disease or Syndrome|History of Present Illness|750,773|false|false|false|C1697454|Pelvic fluid collection|pelvic fluid collection
Drug|Substance|History of Present Illness|757,762|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|757,762|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|History of Present Illness|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|History of Present Illness|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|History of Present Illness|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|History of Present Illness|763,773|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|History of Present Illness|789,794|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|789,794|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Health Care Activity|History of Present Illness|796,805|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|796,805|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Sign or Symptom|History of Present Illness|851,858|false|false|false|C0231218|Malaise|malaise
Finding|Idea or Concept|History of Present Illness|865,868|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|865,868|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Sign or Symptom|History of Present Illness|872,878|false|false|false|C0015967|Fever|fevers
Finding|Body Substance|History of Present Illness|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|883,890|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Substance|History of Present Illness|915,920|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|915,920|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|915,930|false|false|false|C3495845|Drain placement|drain placement
Procedure|Health Care Activity|History of Present Illness|921,930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|921,930|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Finding|Functional Concept|History of Present Illness|936,951|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|History of Present Illness|936,968|false|false|false|C4285843|Intra-abdominal fluid collection|intra-abdominal fluid collection
Drug|Substance|History of Present Illness|952,957|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|History of Present Illness|952,957|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|History of Present Illness|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|History of Present Illness|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|History of Present Illness|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|History of Present Illness|958,968|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|History of Present Illness|973,982|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|History of Present Illness|973,982|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|History of Present Illness|984,991|false|false|true|C0039869;C4319827|Thought|thought
Finding|Mental Process|History of Present Illness|984,991|false|false|true|C0039869;C4319827|Thought|thought
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1021,1024|false|false|false|C0404079|Total abdominal hysterectomy|TAH
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1021,1028|false|false|false|C0542407|Total abdominal hysterectomy with bilateral salpingo-oophorectomy|TAH/BSO
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|History of Present Illness|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|History of Present Illness|1025,1028|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Chemical Viewed Structurally|History of Present Illness|1030,1037|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1030,1048|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1038,1048|false|false|false|C0010651|Cystectomy|cystectomy
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1053,1059|false|false|false|C0030797|Pelvis|pelvic
Finding|Body Substance|History of Present Illness|1061,1066|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1061,1071|false|false|false|C0024204|lymph nodes|lymph node
Procedure|Diagnostic Procedure|History of Present Illness|1061,1078|false|false|false|C0193842|Biopsy of lymph node|lymph node biopsy
Finding|Finding|History of Present Illness|1072,1078|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Finding|Intellectual Product|History of Present Illness|1072,1078|false|false|false|C0220797;C1546569|biopsy characteristics|biopsy
Procedure|Diagnostic Procedure|History of Present Illness|1072,1078|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Procedure|Health Care Activity|History of Present Illness|1072,1078|false|false|false|C0005558;C1548825;C3668914|Biopsy;Biopsy Procedures on the Pharynx, Adenoids, and Tonsils;Consent Type - biopsy|biopsy
Attribute|Clinical Attribute|History of Present Illness|1085,1094|false|false|false|C0945766||procedure
Event|Occupational Activity|History of Present Illness|1085,1094|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|History of Present Illness|1085,1094|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1085,1094|false|false|false|C0184661|Interventional procedure|procedure
Finding|Sign or Symptom|History of Present Illness|1162,1169|false|false|false|C0231218|Malaise|malaise
Finding|Idea or Concept|History of Present Illness|1176,1179|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|1176,1179|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|History of Present Illness|1184,1189|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1184,1189|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1192,1198|false|false|false|C0424790|Rigor - Temperature-associated observation|rigors
Finding|Finding|History of Present Illness|1213,1220|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|History of Present Illness|1216,1220|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1216,1220|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1216,1220|false|false|false|C1553498|home health encounter|home
Finding|Body Substance|History of Present Illness|1242,1250|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|History of Present Illness|1242,1250|false|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1242,1250|false|false|false|C0013103|Drainage procedure|drainage
Finding|Functional Concept|History of Present Illness|1260,1275|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|History of Present Illness|1276,1281|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|1276,1281|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Anatomical Structure|History of Present Illness|1302,1310|false|false|false|C0559495|Urological stoma|urostomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1302,1310|false|false|false|C0856443|Urostomy procedure|urostomy
Finding|Conceptual Entity|History of Present Illness|1311,1317|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|History of Present Illness|1311,1317|false|false|false|C3251815|Measurement of fluid output|output
Finding|Finding|History of Present Illness|1327,1336|false|false|false|C0442739||unchanged
Finding|Intellectual Product|History of Present Illness|1365,1369|false|false|false|C1547225|Mild Severity of Illness Code|mild
Anatomy|Body Location or Region|History of Present Illness|1370,1373|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Finding|Sign or Symptom|History of Present Illness|1370,1378|false|false|false|C0238551|Left lower quadrant pain|LLQ pain
Attribute|Clinical Attribute|History of Present Illness|1374,1378|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1374,1378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1374,1378|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|1391,1399|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1391,1399|true|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|History of Present Illness|1401,1406|false|false|false|C0018932|Hematochezia|BRBPR
Disorder|Disease or Syndrome|History of Present Illness|1408,1412|true|false|false|C5779629|Eruption of skin (disorder)|rash
Finding|Pathologic Function|History of Present Illness|1408,1412|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|1408,1412|true|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Drug|Organic Chemical|History of Present Illness|1414,1419|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1414,1419|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|History of Present Illness|1414,1419|false|false|false|C0010200|Coughing|cough
Finding|Sign or Symptom|History of Present Illness|1422,1430|false|false|false|C0018681|Headache|headache
Anatomy|Body Location or Region|History of Present Illness|1432,1436|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|History of Present Illness|1432,1436|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|History of Present Illness|1432,1436|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Finding|Sign or Symptom|History of Present Illness|1432,1446|false|false|false|C0151315|Neck stiffness|neck stiffness
Finding|Sign or Symptom|History of Present Illness|1437,1446|false|false|false|C0427008|Stiffness|stiffness
Drug|Substance|History of Present Illness|1518,1523|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|History of Present Illness|1518,1523|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Biomedical or Dental Material|History of Present Illness|1524,1531|false|false|false|C1706355|Culture Dose Form|culture
Finding|Functional Concept|History of Present Illness|1524,1531|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|History of Present Illness|1524,1531|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|History of Present Illness|1524,1531|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Drug|Antibiotic|History of Present Illness|1552,1557|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|History of Present Illness|1552,1557|false|false|false|C0250482|Zosyn|zosyn
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1562,1572|false|false|false|C0042313|vancomycin|vancomycin
Drug|Antibiotic|History of Present Illness|1562,1572|false|false|false|C0042313|vancomycin|vancomycin
Procedure|Laboratory Procedure|History of Present Illness|1562,1572|false|false|false|C0489941|Vancomycin measurement|vancomycin
Drug|Organic Chemical|History of Present Illness|1589,1602|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|History of Present Illness|1589,1602|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Procedure|Laboratory Procedure|History of Present Illness|1589,1602|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Event|Occupational Activity|History of Present Illness|1644,1654|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|History of Present Illness|1644,1654|false|false|false|C0376636|Disease Management|management
Disorder|Disease or Syndrome|Past Medical History|1685,1697|false|false|false|C0020538|Hypertensive disease|Hypertension
Disorder|Disease or Syndrome|Past Medical History|1707,1710|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1707,1710|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|Past Medical History|1707,1710|false|false|false|C1870042|ACP2 protein, human|lap
Finding|Finding|Past Medical History|1707,1710|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|Past Medical History|1707,1710|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|Past Medical History|1707,1710|false|false|false|C0031150|Laparoscopy|lap
Finding|Functional Concept|Past Medical History|1726,1730|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Past Medical History|1726,1735|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1726,1735|false|false|false|C0230432;C4281599|Structure of left knee;Structure of left knee region|left knee
Anatomy|Body Location or Region|Past Medical History|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|Past Medical History|1731,1735|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|Past Medical History|1731,1735|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|Past Medical History|1731,1747|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1731,1747|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Finding|Functional Concept|Past Medical History|1736,1747|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|1736,1747|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1736,1747|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1757,1768|false|false|false|C0022983|Laminectomy|laminectomy
Attribute|Clinical Attribute|Past Medical History|1781,1784|false|false|false|C1114365||age
Drug|Biologically Active Substance|Past Medical History|1781,1784|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Past Medical History|1781,1784|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1794,1801|false|false|false|C0005682|Urinary Bladder|Bladder
Disorder|Neoplastic Process|Past Medical History|1794,1801|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|Bladder
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1794,1801|false|false|false|C0872388|Procedures on bladder|Bladder
Disorder|Neoplastic Process|Past Medical History|1794,1808|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|Bladder Cancer
Disorder|Neoplastic Process|Past Medical History|1802,1808|false|false|false|C0006826|Malignant Neoplasms|Cancer
Finding|Finding|Past Medical History|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Past Medical History|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Past Medical History|1809,1813|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Past Medical History|1809,1819|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Intellectual Product|Past Medical History|1809,1819|false|false|false|C0205082;C4554016|Enneking High Surgical Grade;Severe (severity modifier)|high grade
Finding|Classification|Past Medical History|1814,1819|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Past Medical History|1814,1819|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Anatomy|Cell Component|Past Medical History|1820,1823|false|false|false|C1167383|membrane attack complex location|TCC
Disorder|Disease or Syndrome|Past Medical History|1820,1823|false|false|false|C1861305|TARSAL-CARPAL COALITION SYNDROME|TCC
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Biologically Active Substance|Past Medical History|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Organic Chemical|Past Medical History|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Drug|Pharmacologic Substance|Past Medical History|1820,1823|false|false|false|C0077072;C5552697|Membrane Attack Complex;triclocarban|TCC
Finding|Intellectual Product|Past Medical History|1846,1850|false|false|false|C1720594|Then - dosing instruction fragment|then
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1856,1862|false|false|false|C0030797|Pelvis|pelvic
Procedure|Diagnostic Procedure|Past Medical History|1856,1866|false|false|false|C0203201|Magnetic Resonance Imaging (MRI) of Pelvis|pelvic MRI
Finding|Gene or Genome|Past Medical History|1863,1866|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Past Medical History|1863,1866|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Past Medical History|1863,1866|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Disorder|Neoplastic Process|Past Medical History|1869,1877|false|false|false|C1269955|Tumor Cell Invasion|invasion
Finding|Pathologic Function|Past Medical History|1869,1877|false|false|false|C2699153|Cell Invasion|invasion
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1883,1890|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Past Medical History|1883,1890|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1883,1890|false|false|false|C0872388|Procedures on bladder|bladder
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1883,1895|false|false|false|C0458421|Wall of bladder|bladder wall
Disorder|Disease or Syndrome|Past Medical History|1910,1914|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|Past Medical History|1910,1921|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Past Medical History|1910,1921|false|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|Past Medical History|1915,1921|false|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|Past Medical History|1915,1921|false|false|false|C1547928|Tissue Specimen Code|tissue
Disorder|Disease or Syndrome|Past Medical History|1926,1934|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1935,1942|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|1935,1942|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|1935,1942|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|1935,1942|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1935,1947|false|false|false|C0447612|Vaginal wall|vaginal wall
Finding|Functional Concept|Past Medical History|1955,1962|false|false|false|C0332305|With staging|staging
Finding|Finding|Past Medical History|1972,1984|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1972,1984|false|false|false|C0020699|Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1989,2011|false|false|false|C0278321|Bilateral oophorectomy|bilateral oophorectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1999,2011|false|false|false|C0029936|Ovariectomy|oophorectomy
Finding|Gene or Genome|Past Medical History|2016,2021|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|Past Medical History|2016,2028|false|false|false|C0151994|Enlarged uterus|large uterus
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2022,2028|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Anatomy|Tissue|Past Medical History|2022,2028|false|false|false|C0042149;C1519876;C4266525|Mouse Uterus;Pelvis>Uterus;Uterus|uterus
Disorder|Disease or Syndrome|Past Medical History|2022,2028|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Disorder|Neoplastic Process|Past Medical History|2022,2028|false|false|false|C0042131;C0496919|Neoplasm of uncertain or unknown behavior of uterus;Uterine Diseases|uterus
Procedure|Diagnostic Procedure|Past Medical History|2022,2028|false|false|false|C0869889|examination of uterus|uterus
Disorder|Neoplastic Process|Past Medical History|2032,2039|false|false|false|C0023267|Fibroid Tumor|fibroid
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2062,2068|false|false|false|C0030797|Pelvis|pelvic
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2062,2079|false|false|false|C0729595|Pelvic lymph node group|pelvic lymph node
Finding|Body Substance|Past Medical History|2069,2074|false|false|false|C0024202|Lymph|lymph
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2069,2079|false|false|false|C0024204|lymph nodes|lymph node
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2080,2089|false|false|false|C0015252;C0728940|Excision;removal technique|resection
Drug|Chemical Viewed Structurally|Past Medical History|2096,2103|false|false|false|C0302912|Radicals (chemistry)|radical
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2096,2114|false|false|false|C0194401|Complete cystectomy|radical cystectomy
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2104,2114|false|false|false|C0010651|Cystectomy|cystectomy
Disorder|Disease or Syndrome|Past Medical History|2119,2127|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2128,2139|false|false|false|C0195130|Vaginectomy|vaginectomy
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2145,2152|false|false|false|C0042232|Vagina|vaginal
Drug|Biomedical or Dental Material|Past Medical History|2145,2152|false|false|false|C1272941|Vaginal Dosage Form|vaginal
Finding|Finding|Past Medical History|2145,2152|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Finding|Functional Concept|Past Medical History|2145,2152|false|false|false|C1522570;C4521343|Vaginal (intended site);Vaginal Route of Administration|vaginal
Procedure|Machine Activity|Past Medical History|2154,2168|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2154,2168|false|false|false|C0020912;C0524865|Optical Image Reconstruction;Reconstructive Surgical Procedures|reconstruction
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2174,2179|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|Past Medical History|2174,2187|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2174,2187|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Event|Activity|Past Medical History|2188,2196|false|false|false|C1706214|Creation|creation
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2188,2196|false|false|false|C0441513|Surgical construction|creation
Finding|Finding|Past Medical History|2225,2235|false|false|false|C0004610|Bacteremia|bacteremia
Finding|Functional Concept|Past Medical History|2240,2251|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Organism Function|Past Medical History|2240,2251|false|false|false|C0018271;C0243107;C0678723;C1527148|Development;Growth and Development function;biological development;development aspects|development
Finding|Functional Concept|Past Medical History|2255,2270|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Drug|Substance|Past Medical History|2272,2277|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Past Medical History|2272,2277|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Past Medical History|2278,2288|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Past Medical History|2278,2288|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Past Medical History|2278,2288|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Past Medical History|2278,2288|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|Past Medical History|2297,2302|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Past Medical History|2297,2302|false|false|false|C1546604|Drain Specimen Code|drain
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2297,2312|false|false|false|C3495845|Drain placement|drain placement
Procedure|Health Care Activity|Past Medical History|2303,2312|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2303,2312|false|false|false|C0021107;C0441587;C1533810|Clinical act of insertion;Implantation procedure|placement
Anatomy|Body Location or Region|Past Medical History|2337,2340|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Past Medical History|2337,2340|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Past Medical History|2337,2340|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Organic Chemical|Past Medical History|2351,2358|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Past Medical History|2351,2358|false|false|false|C0728963|Lovenox|lovenox
Finding|Classification|Family Medical History|2400,2408|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Finding|Finding|Family Medical History|2400,2408|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|Negative
Lab|Laboratory or Test Result|Family Medical History|2400,2408|false|false|false|C5237010|Expression Negative|Negative
Finding|Finding|Family Medical History|2400,2412|false|false|false|C0205160|Negative|Negative for
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2413,2420|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Family Medical History|2413,2420|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2413,2420|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Family Medical History|2413,2423|false|true|false|C0005684|Malignant neoplasm of urinary bladder|bladder CA
Procedure|Health Care Activity|General Exam|2443,2452|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Functional Concept|General Exam|2453,2457|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2453,2457|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|General Exam|2476,2481|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|General Exam|2476,2487|false|false|false|C0488614;C0518766|Vital signs|Vital Signs
Procedure|Health Care Activity|General Exam|2476,2487|false|false|false|C0150404|Taking vital signs|Vital Signs
Finding|Finding|General Exam|2482,2487|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Functional Concept|General Exam|2482,2487|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|Signs
Finding|Individual Behavior|General Exam|2509,2514|false|false|false|C0600261|Telling untruths|Lying
Finding|Classification|General Exam|2530,2537|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|2530,2537|false|false|false|C3812897|General medical service|General
Attribute|Clinical Attribute|General Exam|2539,2544|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|2539,2544|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|2539,2544|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|General Exam|2539,2544|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|2539,2544|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2539,2544|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2559,2564|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|2565,2573|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2565,2573|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|2577,2582|false|false|false|C1512338|HEENT|HEENT
Finding|Finding|General Exam|2592,2601|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2603,2606|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|2603,2606|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|2608,2618|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|2619,2624|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Organ or Tissue Function|General Exam|2651,2659|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|2651,2666|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Finding|Finding|General Exam|2660,2666|false|false|false|C0018808|Heart murmur|murmur
Finding|Finding|General Exam|2667,2671|false|false|false|C0232267|Pericardial friction rub|RUBS
Finding|Finding|General Exam|2676,2680|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2693,2698|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|2700,2705|false|false|false|C1550016|Remote control command - Clear|Clear
Procedure|Diagnostic Procedure|General Exam|2709,2721|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|General Exam|2738,2745|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|General Exam|2747,2752|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|General Exam|2755,2762|false|false|false|C0035508|Rhonchi|rhonchi
Anatomy|Body Location or Region|General Exam|2766,2773|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2766,2773|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|2766,2773|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2775,2779|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|2808,2813|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|2808,2820|false|false|false|C0232693|Bowel sounds|bowel sounds
Phenomenon|Natural Phenomenon or Process|General Exam|2814,2820|false|false|false|C0037709||sounds
Finding|Finding|General Exam|2821,2828|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|2821,2828|false|false|false|C0150312;C0449450|Present;Presentation|present
Anatomy|Body Part, Organ, or Organ Component|General Exam|2832,2837|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|General Exam|2832,2845|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|General Exam|2832,2845|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Drug|Substance|General Exam|2846,2851|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|2846,2851|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Location or Region|General Exam|2855,2858|false|false|false|C0230178|Structure of right lower quadrant of abdomen|RLQ
Drug|Substance|General Exam|2873,2878|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|2873,2878|false|false|false|C1546604|Drain Specimen Code|drain
Anatomy|Body Location or Region|General Exam|2882,2885|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Finding|Gene or Genome|General Exam|2901,2905|false|false|false|C1864650|GNAS-AS1 gene|sang
Drug|Substance|General Exam|2906,2911|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|2906,2911|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Congenital Abnormality|General Exam|2931,2934|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|2931,2934|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|2936,2940|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2936,2940|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2942,2946|false|false|false|C5575035|Well (answer to question)|well
Attribute|Clinical Attribute|General Exam|2971,2976|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|2971,2976|false|false|false|C0013604|Edema|edema
Finding|Gene or Genome|General Exam|2991,2994|false|false|false|C1539110|CNDP2 gene|CN2
Finding|Finding|General Exam|3006,3012|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|3021,3036|false|false|false|C0278454|All extremities|all extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3025,3036|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Body Substance|General Exam|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3053,3062|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3053,3062|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Functional Concept|General Exam|3063,3067|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3063,3067|false|false|false|C0582103|Medical Examination|EXAM
Drug|Food|General Exam|3087,3092|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|Vital
Attribute|Clinical Attribute|General Exam|3087,3098|false|false|false|C0488614;C0518766|Vital signs|Vital signs
Procedure|Health Care Activity|General Exam|3087,3098|false|false|false|C0150404|Taking vital signs|Vital signs
Finding|Finding|General Exam|3093,3098|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|General Exam|3093,3098|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Classification|General Exam|3130,3137|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3130,3137|false|false|false|C3812897|General medical service|General
Anatomy|Body Location or Region|General Exam|3147,3152|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3154,3160|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3154,3160|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|3154,3160|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|3161,3170|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Location or Region|General Exam|3172,3176|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3172,3176|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3172,3176|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|General Exam|3178,3184|false|false|false|C0332254|Supple|supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3187,3192|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|3194,3199|false|false|false|C1550016|Remote control command - Clear|Clear
Procedure|Diagnostic Procedure|General Exam|3203,3215|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|General Exam|3232,3239|true|false|false|C0043144|Wheezing|wheezes
Finding|Finding|General Exam|3241,3246|false|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Finding|Finding|General Exam|3249,3256|false|false|false|C0035508|Rhonchi|rhonchi
Disorder|Disease or Syndrome|General Exam|3260,3268|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Procedure|Diagnostic Procedure|General Exam|3269,3281|false|false|false|C0004339|Auscultation|auscultation
Event|Activity|General Exam|3296,3300|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|3296,3300|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|3305,3311|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3305,3311|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|General Exam|3336,3339|false|false|false|C0694547|SYSTOLIC EJECTION MURMUR|SEM
Anatomy|Body Location or Region|General Exam|3341,3348|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|3341,3348|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|3341,3348|false|false|false|C0941288|Abdomen problem|Abdomen
Anatomy|Body Part, Organ, or Organ Component|General Exam|3355,3360|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|General Exam|3355,3368|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|General Exam|3355,3368|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Finding|Idea or Concept|General Exam|3378,3383|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Body Substance|General Exam|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|General Exam|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|General Exam|3391,3396|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Location or Region|General Exam|3408,3411|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|General Exam|3412,3417|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|3412,3417|false|false|false|C1546604|Drain Specimen Code|drain
Event|Activity|General Exam|3421,3426|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|3421,3426|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|3421,3426|false|false|false|C1533810||place
Finding|Body Substance|General Exam|3436,3456|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|General Exam|3451,3456|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|3451,3456|false|false|false|C1546638|Fluid Specimen Code|fluid
Disorder|Congenital Abnormality|General Exam|3460,3463|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|3460,3463|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|3465,3469|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3465,3469|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3471,3475|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|3489,3495|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3489,3495|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3489,3495|false|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|3500,3508|true|false|false|C0149651|Clubbing|clubbing
Finding|Sign or Symptom|General Exam|3510,3518|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|3523,3528|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|3523,3528|false|false|false|C0013604|Edema|edema
Procedure|Health Care Activity|General Exam|3552,3561|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|3562,3566|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3596,3601|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3596,3601|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3602,3605|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3613,3616|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3613,3616|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3613,3616|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3623,3626|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3623,3626|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3623,3626|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3623,3626|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3632,3635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3632,3635|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3643,3646|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3643,3646|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3643,3646|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3643,3646|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3650,3653|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3650,3653|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3650,3653|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3650,3653|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3650,3653|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3659,3663|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3691,3694|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3711,3716|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3711,3716|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3729,3735|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3741,3746|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3752,3755|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|3752,3755|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3859,3864|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3859,3864|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3869,3872|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|3869,3872|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3894,3899|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3894,3899|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|3900,3903|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|General Exam|3900,3903|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|General Exam|3900,3903|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Congenital Abnormality|General Exam|3913,3916|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Disorder|Disease or Syndrome|General Exam|3913,3916|false|false|false|C0002636;C0220724|Amniotic Band Syndrome;CONSTRICTING BANDS, CONGENITAL|Abs
Finding|Gene or Genome|General Exam|3913,3916|false|false|false|C1425698;C4723885|DDX41 gene;DDX41 wt Allele|Abs
Drug|Amino Acid, Peptide, or Protein|General Exam|3917,3920|false|false|false|C0389252|RET protein, human|Ret
Finding|Gene or Genome|General Exam|3917,3920|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Finding|Receptor|General Exam|3917,3920|false|false|false|C0389252;C0694890;C0813143;C1704885|Oncogene RET;RET gene;RET protein, human;RET wt Allele|Ret
Disorder|Disease or Syndrome|General Exam|3938,3943|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3938,3943|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3938,3951|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3938,3951|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3938,3951|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3944,3951|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3944,3951|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3944,3951|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|3944,3951|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3944,3951|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|3997,4001|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|3997,4001|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|3997,4001|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4026,4031|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4026,4031|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4032,4035|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4032,4035|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4032,4035|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|General Exam|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4032,4035|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4032,4035|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4038,4041|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4038,4041|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4038,4041|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|General Exam|4038,4041|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4044,4051|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4044,4051|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4079,4084|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4079,4084|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4085,4091|false|false|false|C0023764|lipase|Lipase
Drug|Enzyme|General Exam|4085,4091|false|false|false|C0023764|lipase|Lipase
Drug|Pharmacologic Substance|General Exam|4085,4091|false|false|false|C0023764|lipase|Lipase
Procedure|Laboratory Procedure|General Exam|4085,4091|false|false|false|C0373670|Lipase measurement|Lipase
Disorder|Disease or Syndrome|General Exam|4106,4111|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4106,4111|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4106,4119|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4112,4119|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Finding|Gene or Genome|General Exam|4112,4119|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4112,4119|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4112,4119|false|false|false|C0201838|Albumin measurement|Albumin
Drug|Biologically Active Substance|General Exam|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|General Exam|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|General Exam|4125,4129|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|General Exam|4125,4129|false|false|false|C0337439|Iron measurement|Iron
Disorder|Disease or Syndrome|General Exam|4145,4150|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4145,4150|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|4189,4192|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|4189,4192|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Disorder|Disease or Syndrome|General Exam|4210,4215|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4210,4215|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4210,4223|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|4216,4223|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|4216,4223|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Procedure|Laboratory Procedure|General Exam|4216,4223|false|false|false|C0202115|Lactic acid measurement|Lactate
Finding|Body Substance|General Exam|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4229,4238|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4229,4238|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|General Exam|4239,4243|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4273,4278|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4273,4278|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4279,4282|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4287,4290|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4287,4290|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4287,4290|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4297,4300|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4297,4300|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4297,4300|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4297,4300|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4306,4309|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4306,4309|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4317,4320|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4317,4320|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4317,4320|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4317,4320|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4324,4327|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4324,4327|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4324,4327|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4324,4327|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4324,4327|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4333,4337|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4365,4368|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4385,4390|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4385,4390|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4395,4398|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4395,4398|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4420,4425|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4420,4425|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4426,4429|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4446,4451|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4446,4451|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4446,4459|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4446,4459|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4446,4459|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4452,4459|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4452,4459|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4452,4459|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4452,4459|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4452,4459|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4502,4506|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4502,4506|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4502,4506|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4531,4536|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4531,4536|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4531,4544|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4537,4544|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|General Exam|4537,4544|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4537,4544|false|false|false|C0201925|Calcium measurement|Calcium
Finding|Functional Concept|General Exam|4567,4579|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Finding|Intellectual Product|General Exam|4567,4579|false|false|false|C0025953;C1571921;C4049106|Microbiological;Microbiology - Laboratory Class;Microbiology Diagnostic Service Section ID|MICROBIOLOGY
Procedure|Laboratory Procedure|General Exam|4567,4579|false|false|false|C0085672|Microbiology procedure|MICROBIOLOGY
Disorder|Disease or Syndrome|General Exam|4595,4600|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|4595,4600|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Procedure|Laboratory Procedure|General Exam|4595,4609|false|true|false|C0200949|Blood culture|Blood cultures
Finding|Idea or Concept|General Exam|4601,4609|false|false|false|C0010453|Culture (Anthropological)|cultures
Finding|Idea or Concept|General Exam|4613,4620|false|false|false|C1691786;C1704475|Pending - Allergy Clinical Status;Pending - referral status|pending
Anatomy|Body Part, Organ, or Organ Component|General Exam|4634,4640|false|false|false|C0030797|Pelvis|pelvic
Disorder|Injury or Poisoning|General Exam|4641,4651|false|false|false|C1720922|Respiratory Aspiration|aspiration
Finding|Finding|General Exam|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Organ or Tissue Function|General Exam|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Finding|Pathologic Function|General Exam|4641,4651|false|false|false|C0220787;C0700198;C2712334|Aspiration into respiratory tract;Endotracheal aspiration;Pulmonary aspiration|aspiration
Procedure|Therapeutic or Preventive Procedure|General Exam|4641,4651|false|false|false|C0349707||aspiration
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4655,4665|false|false|false|C0061856|Gram's stain|GRAM STAIN
Drug|Organic Chemical|General Exam|4655,4665|false|false|false|C0061856|Gram's stain|GRAM STAIN
Procedure|Laboratory Procedure|General Exam|4655,4665|false|false|false|C0200966|Bacterial stain, routine|GRAM STAIN
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4660,4665|false|false|false|C0038128|Stains|STAIN
Procedure|Laboratory Procedure|General Exam|4660,4665|false|false|false|C0487602|Staining method|STAIN
Finding|Idea or Concept|General Exam|4667,4672|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Conceptual Entity|General Exam|4705,4710|false|false|false|C1521738;C2346620;C2349184|Field;Force Field;Knowledge Field|FIELD
Procedure|Health Care Activity|General Exam|4705,4710|false|false|false|C1553496|field - patient encounter|FIELD
Anatomy|Cell|General Exam|4734,4744|false|false|false|C0023516|Leukocytes|LEUKOCYTES
Finding|Body Substance|General Exam|4734,4744|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Intellectual Product|General Exam|4734,4744|false|false|false|C1547962;C1550647|Specimen Type - Leukocytes|LEUKOCYTES
Finding|Finding|General Exam|4756,4775|false|false|false|C2924473|Microorganisms seen|MICROORGANISMS SEEN
Drug|Substance|General Exam|4781,4786|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|FLUID
Finding|Intellectual Product|General Exam|4781,4786|false|false|false|C1546638|Fluid Specimen Code|FLUID
Drug|Biomedical or Dental Material|General Exam|4787,4794|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|4787,4794|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4787,4794|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4787,4794|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Idea or Concept|General Exam|4796,4801|false|false|false|C1546485|Diagnosis Type - Final|Final
Finding|Finding|General Exam|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4813,4819|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4813,4819|true|false|false|C2911660|Growth action|GROWTH
Procedure|Laboratory Procedure|General Exam|4825,4842|false|false|false|C1273935|Anaerobic microbial culture|ANAEROBIC CULTURE
Drug|Biomedical or Dental Material|General Exam|4835,4842|false|false|false|C1706355|Culture Dose Form|CULTURE
Finding|Functional Concept|General Exam|4835,4842|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Finding|Idea or Concept|General Exam|4835,4842|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|CULTURE
Procedure|Laboratory Procedure|General Exam|4835,4842|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|CULTURE
Finding|Finding|General Exam|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organ or Tissue Function|General Exam|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Organism Function|General Exam|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Finding|Physiologic Function|General Exam|4864,4870|true|false|false|C0018270;C0220844;C1457898;C1621966|Growth;Growth & development aspects;Tissue Growth;growth aspects|GROWTH
Phenomenon|Phenomenon or Process|General Exam|4864,4870|true|false|false|C2911660|Growth action|GROWTH
Finding|Finding|General Exam|4884,4891|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4884,4891|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Attribute|Clinical Attribute|General Exam|4912,4918|false|false|false|C1644645||CT ABD
Anatomy|Body Location or Region|General Exam|4915,4918|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|4915,4918|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Anatomy|Body Location or Region|General Exam|4919,4922|false|false|false|C0449203|PEL (body structure)|PEL
Disorder|Disease or Syndrome|General Exam|4919,4922|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|PEL
Disorder|Neoplastic Process|General Exam|4919,4922|false|false|false|C1292753;C1394210;C4520841|Pel crisis;Primary Effusion Lymphoma;Pure Erythroid Leukemia|PEL
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|4926,4934|false|false|false|C0009924|Contrast Media|CONTRAST
Finding|Intellectual Product|General Exam|4943,4951|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Finding|Finding|General Exam|4952,4960|false|false|false|C0392756|Reduced|decrease
Finding|Functional Concept|General Exam|4976,4981|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Drug|Substance|General Exam|4993,4998|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|4993,4998|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|General Exam|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5000,5010|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|General Exam|5077,5085|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Finding|Functional Concept|General Exam|5086,5094|false|false|false|C5445118|Approach (contact)|approach
Finding|Intellectual Product|General Exam|5103,5111|false|false|false|C1546572||catheter
Finding|Finding|General Exam|5112,5121|false|false|false|C0442739||unchanged
Finding|Conceptual Entity|General Exam|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5185,5195|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5229,5237|false|false|false|C1552654|Parameterized Data Type - Interval|Interval
Finding|Functional Concept|General Exam|5238,5246|false|false|false|C0442805|Increase|increase
Finding|Finding|General Exam|5238,5254|false|false|false|C1268652|increase in size|increase in size
Finding|Functional Concept|General Exam|5262,5266|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5267,5273|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|General Exam|5274,5279|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|5274,5279|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|General Exam|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5281,5291|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Event|Activity|General Exam|5388,5399|false|false|false|C2349975|Enhance (action)|enhancement
Procedure|Therapeutic or Preventive Procedure|General Exam|5388,5399|false|false|false|C1627358|Refractive surgery enhancement|enhancement
Disorder|Disease or Syndrome|General Exam|5426,5435|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|General Exam|5426,5435|false|false|false|C3714514|Infection|infection
Finding|Finding|General Exam|5444,5447|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|General Exam|5444,5447|true|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|General Exam|5448,5453|true|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|5448,5453|true|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|General Exam|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5454,5464|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Amino Acid, Peptide, or Protein|General Exam|5481,5484|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Finding|Gene or Genome|General Exam|5481,5484|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|5481,5484|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|5485,5488|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|5485,5488|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Anatomy|Body Part, Organ, or Organ Component|General Exam|5491,5497|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Anatomy|Body Space or Junction|General Exam|5491,5497|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|PELVIS
Disorder|Neoplastic Process|General Exam|5491,5497|false|false|false|C0153663|Malignant neoplasm of pelvis|PELVIS
Finding|Finding|General Exam|5491,5497|false|false|false|C0812455|Pelvis problem|PELVIS
Finding|Finding|General Exam|5505,5513|false|false|false|C0392756|Reduced|Decrease
Finding|Functional Concept|General Exam|5525,5530|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|5525,5545|false|false|false|C0230178|Structure of right lower quadrant of abdomen|right lower quadrant
Anatomy|Body Location or Region|General Exam|5531,5536|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|5531,5536|false|false|false|C2003888|Lower (action)|lower
Drug|Substance|General Exam|5546,5551|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|5546,5551|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|General Exam|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5552,5562|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5574,5586|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Drug|Substance|General Exam|5587,5592|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|General Exam|5587,5592|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Finding|General Exam|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|General Exam|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|General Exam|5618,5622|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Activity|General Exam|5623,5634|false|false|false|C0599946|Attenuation|attenuation
Finding|Functional Concept|General Exam|5651,5655|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|General Exam|5651,5655|false|false|false|C0582103|Medical Examination|exam
Finding|Idea or Concept|General Exam|5656,5666|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|General Exam|5656,5671|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|General Exam|5672,5677|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|General Exam|5672,5677|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Pharmacologic Substance|General Exam|5672,5686|false|false|false|C0456388|Blood product|blood products
Disorder|Disease or Syndrome|General Exam|5704,5713|false|false|false|C0020452|Hyperemia|hyperemia
Finding|Finding|General Exam|5723,5729|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5723,5729|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|General Exam|5723,5742|false|false|false|C4050249|Likely Inflammatory Activity|likely inflammatory
Finding|Functional Concept|General Exam|5730,5742|false|true|false|C0333348|Inflammatory|inflammatory
Finding|Idea or Concept|General Exam|5756,5764|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|5756,5767|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|5769,5777|false|false|false|C0009924|Contrast Media|contrast
Disorder|Injury or Poisoning|General Exam|5778,5791|false|false|false|C0015379|Extravasation of Diagnostic and Therapeutic Materials|extravasation
Finding|Pathologic Function|General Exam|5778,5791|false|false|false|C0015376|Extravasation|extravasation
Finding|Gene or Genome|General Exam|5806,5811|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Intellectual Product|General Exam|5812,5818|false|false|false|C1547311|Patient Condition Code - Stable|stable
Drug|Substance|General Exam|5819,5824|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|5819,5824|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|General Exam|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|5825,5835|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Finding|General Exam|5843,5846|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|5843,5846|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Functional Concept|General Exam|5847,5851|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|5853,5860|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|5853,5860|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|5853,5860|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|General Exam|5862,5868|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|5862,5868|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|5862,5868|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|5862,5868|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Intellectual Product|General Exam|5874,5878|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Activity|General Exam|5897,5908|false|false|false|C2349975|Enhance (action)|enhancement
Procedure|Therapeutic or Preventive Procedure|General Exam|5897,5908|false|false|false|C1627358|Refractive surgery enhancement|enhancement
Disorder|Disease or Syndrome|General Exam|5911,5920|false|true|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|General Exam|5911,5920|false|true|false|C3714514|Infection|infection
Finding|Finding|General Exam|5954,5960|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|5954,5960|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|General Exam|5961,5965|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|General Exam|5971,5979|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|General Exam|5971,5979|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Finding|General Exam|5983,5989|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|5983,5989|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Functional Concept|General Exam|5990,5995|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Disease or Syndrome|General Exam|5997,6018|false|false|false|C0268804|Hydroureteronephrosis|hydroureteronephrosis
Finding|Functional Concept|General Exam|6033,6037|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Intellectual Product|General Exam|6050,6056|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|General Exam|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Gene or Genome|General Exam|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Intellectual Product|General Exam|6071,6075|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|Mass
Finding|Finding|General Exam|6071,6082|false|false|false|C4086564|Mass Effect|Mass effect
Anatomy|Body Space or Junction|General Exam|6089,6100|false|false|false|C0500470|Anatomical anastomosis|anastomosis
Disorder|Acquired Abnormality|General Exam|6089,6100|false|false|false|C0332853|Anastomosis|anastomosis
Procedure|Therapeutic or Preventive Procedure|General Exam|6089,6100|false|false|false|C0677554||anastomosis
Attribute|Clinical Attribute|General Exam|6109,6115|false|false|false|C4522154|Distal Resection Margin|distal
Anatomy|Body Part, Organ, or Organ Component|General Exam|6116,6123|false|false|false|C0041951|Ureter|ureters
Anatomy|Anatomical Structure|General Exam|6129,6139|false|false|false|C3898148|Neobladder|neobladder
Disorder|Disease or Syndrome|General Exam|6179,6193|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Attribute|Clinical Attribute|General Exam|6215,6220|false|false|false|C1717255||edema
Finding|Pathologic Function|General Exam|6215,6220|false|false|false|C0013604|Edema|edema
Finding|Functional Concept|General Exam|6261,6271|false|false|false|C0015127|Etiology aspects|etiologies
Finding|Pathologic Function|General Exam|6282,6290|false|false|false|C1261287|Stenosis|stenosis
Disorder|Neoplastic Process|General Exam|6292,6297|false|false|false|C0027651|Neoplasms|tumor
Finding|Finding|General Exam|6292,6297|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Intellectual Product|General Exam|6292,6297|false|false|false|C1578706;C3273930|Tumor Mass|tumor
Finding|Functional Concept|General Exam|6299,6311|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Finding|Pathologic Function|General Exam|6299,6311|false|false|false|C0332448;C1523986;C3669041|Infiltration;Infiltration Route of Administration;Spread by direct extension|infiltration
Procedure|Therapeutic or Preventive Procedure|General Exam|6299,6311|false|false|false|C0702249|Infiltration (procedure)|infiltration
Anatomy|Body Location or Region|General Exam|6341,6348|false|false|false|C0205054|Hepatic|hepatic
Finding|Finding|General Exam|6341,6355|false|false|false|C0577053|Lesion of liver|hepatic lesion
Finding|Finding|General Exam|6349,6355|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|6349,6355|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|General Exam|6369,6378|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|General Exam|6369,6378|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Event|Governmental or Regulatory Activity|General Exam|6387,6391|false|false|false|C1510751|Academic Research Enhancement Awards|area
Procedure|Diagnostic Procedure|General Exam|6436,6450|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|INTERVENTIONAL
Procedure|Therapeutic or Preventive Procedure|General Exam|6436,6450|false|false|false|C0184661;C2183254|Interventional procedure;interventional (invasive) radiology|INTERVENTIONAL
Procedure|Therapeutic or Preventive Procedure|General Exam|6436,6460|false|false|false|C0184661|Interventional procedure|INTERVENTIONAL PROCEDURE
Attribute|Clinical Attribute|General Exam|6451,6460|false|false|false|C0945766||PROCEDURE
Event|Occupational Activity|General Exam|6451,6460|false|false|false|C1546467|Act Class - procedure|PROCEDURE
Finding|Functional Concept|General Exam|6451,6460|false|false|false|C2700391|Procedure (set of actions)|PROCEDURE
Procedure|Therapeutic or Preventive Procedure|General Exam|6451,6460|false|false|false|C0184661|Interventional procedure|PROCEDURE
Drug|Organic Chemical|General Exam|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Pharmacologic Substance|General Exam|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Drug|Vitamin|General Exam|6470,6478|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|Complete
Finding|Functional Concept|General Exam|6470,6478|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Finding|Idea or Concept|General Exam|6470,6478|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|Complete
Finding|Finding|General Exam|6479,6487|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Finding|Pathologic Function|General Exam|6479,6487|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Phenomenon|Phenomenon or Process|General Exam|6479,6487|false|false|false|C0332521|Collapse (morphologic abnormality)|collapse
Finding|Body Substance|General Exam|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6492,6499|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|General Exam|6492,6503|false|false|false|C0332310|Has patient|patient has
Finding|Functional Concept|General Exam|6521,6525|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|6527,6532|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|6527,6532|false|false|false|C2003888|Lower (action)|lower
Finding|Conceptual Entity|General Exam|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|6543,6553|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|6560,6568|false|false|false|C1546572||catheter
Finding|Conceptual Entity|General Exam|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|6579,6589|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Finding|General Exam|6608,6621|false|false|false|C4489118|Near complete|Near complete
Drug|Organic Chemical|General Exam|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|General Exam|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|General Exam|6613,6621|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|General Exam|6613,6621|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|6613,6621|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Finding|General Exam|6622,6630|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Finding|Pathologic Function|General Exam|6622,6630|false|false|false|C0036974;C0344329;C2210463|Collapse (finding);Shock|collapse
Phenomenon|Phenomenon or Process|General Exam|6622,6630|false|false|false|C0332521|Collapse (morphologic abnormality)|collapse
Finding|Body Substance|General Exam|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6638,6645|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Conceptual Entity|General Exam|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|6669,6679|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Anatomy|Body Part, Organ, or Organ Component|General Exam|6691,6697|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|General Exam|6691,6697|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|General Exam|6691,6697|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|General Exam|6691,6697|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Intellectual Product|General Exam|6712,6720|false|false|false|C1546572||catheter
Event|Activity|General Exam|6724,6729|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|General Exam|6724,6729|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|General Exam|6724,6729|false|false|false|C1533810||place
Finding|Functional Concept|General Exam|6736,6740|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Location or Region|General Exam|6736,6755|false|false|false|C0230180|Structure of left lower quadrant of abdomen|Left lower quadrant
Anatomy|Body Location or Region|General Exam|6741,6746|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|6741,6746|false|false|false|C2003888|Lower (action)|lower
Attribute|Clinical Attribute|General Exam|6760,6764|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|General Exam|6765,6771|false|false|false|C0030797|Pelvis|pelvic
Finding|Idea or Concept|General Exam|6787,6792|false|false|false|C1552828|Table Frame - above|above
Attribute|Clinical Attribute|General Exam|6802,6810|false|false|true|C2926606||findings
Finding|Functional Concept|General Exam|6802,6810|false|false|true|C2607943|findings aspects|findings
Finding|Body Substance|General Exam|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6853,6860|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6873,6881|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Attribute|Clinical Attribute|General Exam|6873,6888|false|false|false|C0449440;C5890498|Clinical status|clinical status
Attribute|Clinical Attribute|General Exam|6882,6888|false|false|false|C5889824||status
Finding|Idea or Concept|General Exam|6882,6888|false|false|false|C1546481|What subject filter - Status|status
Finding|Mental Process|General Exam|6894,6902|false|false|false|C0679006|Decision|decision
Finding|Conceptual Entity|General Exam|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|General Exam|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|General Exam|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|General Exam|6934,6944|true|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Body Substance|General Exam|6945,6953|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Finding|Sign or Symptom|General Exam|6945,6953|true|false|false|C0012621;C2926602|Body Fluid Discharge;Body Substance Discharge|drainage
Procedure|Therapeutic or Preventive Procedure|General Exam|6945,6953|true|false|false|C0013103|Drainage procedure|drainage
Finding|Finding|General Exam|6962,6966|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|General Exam|6962,6966|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|General Exam|6962,6966|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|General Exam|6973,6979|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Finding|Intellectual Product|General Exam|6973,6979|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|Severe
Disorder|Disease or Syndrome|General Exam|6980,7004|false|false|false|C0521622|Bilateral hydronephrosis|bilateral hydronephrosis
Disorder|Disease or Syndrome|General Exam|6990,7004|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Procedure|Health Care Activity|General Exam|7018,7030|false|false|false|C0031809|Physical Examination|examinations
Finding|Idea or Concept|General Exam|7033,7047|false|false|false|C0034866|Recommendation|RECOMMENDATION
Finding|Mental Process|General Exam|7056,7067|false|false|false|C0546816|Persistence|persistence
Finding|Finding|General Exam|7071,7077|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|General Exam|7071,7077|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|General Exam|7071,7092|false|false|false|C0237061|Severe hydronephrosis|severe hydronephrosis
Disorder|Disease or Syndrome|General Exam|7078,7092|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Finding|Functional Concept|General Exam|7095,7107|false|false|false|C1522243|Percutaneous Route of Drug Administration|percutaneous
Finding|Finding|General Exam|7109,7120|false|false|false|C0481713|Has nephrostomy|nephrostomy
Procedure|Therapeutic or Preventive Procedure|General Exam|7109,7120|false|false|false|C0278314|Nephrostomy (procedure)|nephrostomy
Finding|Intellectual Product|General Exam|7121,7126|false|false|false|C1547937||tubes
Finding|Intellectual Product|Hospital Course|7176,7181|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|BRIEF
Finding|Intellectual Product|Hospital Course|7182,7189|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|SUMMARY
Finding|Idea or Concept|Hospital Course|7210,7214|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|7210,7214|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Conceptual Entity|Hospital Course|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|7232,7239|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|7232,7242|false|false|false|C0262926|Medical History|history of
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7243,7250|false|false|false|C0005682|Urinary Bladder|bladder
Disorder|Neoplastic Process|Hospital Course|7243,7250|false|false|false|C0154017;C0154091;C0496930|Benign neoplasm of bladder;Carcinoma in situ of bladder;Neoplasm of uncertain or unknown behavior of bladder|bladder
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7243,7250|false|false|false|C0872388|Procedures on bladder|bladder
Disorder|Neoplastic Process|Hospital Course|7243,7257|false|false|false|C0005684;C0005695;C0699885|Bladder Neoplasm;Carcinoma of bladder;Malignant neoplasm of urinary bladder|bladder cancer
Disorder|Neoplastic Process|Hospital Course|7251,7257|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7263,7273|false|false|false|C0010651|Cystectomy|cystectomy
Finding|Finding|Hospital Course|7275,7287|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7275,7287|false|false|false|C0020699|Hysterectomy|hysterectomy
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|Hospital Course|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|Hospital Course|7293,7296|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7306,7311|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|Hospital Course|7306,7319|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7306,7319|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Finding|Finding|Hospital Course|7328,7342|false|false|false|C0241311|post operative (finding)|post operative
Anatomy|Body Location or Region|Hospital Course|7374,7377|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7374,7377|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7374,7377|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Disease or Syndrome|Hospital Course|7382,7387|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7394,7400|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|Hospital Course|7401,7406|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|7401,7406|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Hospital Course|7426,7429|false|false|false|C0230180|Structure of left lower quadrant of abdomen|LLQ
Drug|Substance|Hospital Course|7430,7435|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|7430,7435|false|false|false|C1546604|Drain Specimen Code|drain
Attribute|Clinical Attribute|Hospital Course|7452,7462|false|false|false|C2979880||subjective
Finding|Finding|Hospital Course|7452,7462|false|false|false|C2266644|subjective (symptom)|subjective
Finding|Sign or Symptom|Hospital Course|7463,7469|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|Hospital Course|7471,7479|false|false|false|C0023380|Lethargy|lethargy
Finding|Finding|Hospital Course|7485,7491|false|false|false|C4554530|Bloody|bloody
Drug|Substance|Hospital Course|7492,7497|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|7492,7497|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Conceptual Entity|Hospital Course|7498,7504|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|7498,7504|false|false|false|C3251815|Measurement of fluid output|output
Finding|Idea or Concept|Hospital Course|7529,7538|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|Hospital Course|7539,7545|false|false|false|C0002871|Anemia|anemia
Finding|Functional Concept|Hospital Course|7594,7602|false|false|false|C0442805|Increase|increase
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Biologically Active Substance|Hospital Course|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Organic Chemical|Hospital Course|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Drug|Pharmacologic Substance|Hospital Course|7606,7616|false|false|false|C0008721;C0019046|Hemoglobin;chrysarobin|hemoglobin
Finding|Finding|Hospital Course|7606,7616|false|false|false|C1561562|Hemoglobin finding|hemoglobin
Procedure|Laboratory Procedure|Hospital Course|7606,7616|false|false|false|C0518015|Hemoglobin measurement|hemoglobin
Finding|Finding|Hospital Course|7650,7657|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|7650,7657|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Intellectual Product|Hospital Course|7669,7677|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Finding|Functional Concept|Hospital Course|7678,7686|false|false|false|C0442805|Increase|increase
Finding|Finding|Hospital Course|7678,7694|false|false|false|C1268652|increase in size|increase in size
Finding|Functional Concept|Hospital Course|7701,7705|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Hospital Course|7706,7715|false|false|false|C0000726|Abdomen|abdominal
Finding|Body Substance|Hospital Course|7706,7721|false|false|false|C2699330|Abdominal Fluid|abdominal fluid
Drug|Substance|Hospital Course|7716,7721|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|7716,7721|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|7722,7732|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Mental Process|Hospital Course|7734,7742|false|false|false|C0679006|Decision|Decision
Event|Activity|Hospital Course|7755,7760|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|7755,7760|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|7755,7760|false|false|false|C1533810||place
Drug|Substance|Hospital Course|7764,7769|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|7764,7769|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|Hospital Course|7778,7783|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|Hospital Course|7778,7783|false|false|false|C1546638|Fluid Specimen Code|Fluid
Finding|Classification|Hospital Course|7807,7815|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7807,7815|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7807,7815|false|false|false|C5237010|Expression Negative|negative
Finding|Idea or Concept|Hospital Course|7816,7824|false|true|false|C0010453|Culture (Anthropological)|cultures
Finding|Classification|Hospital Course|7827,7835|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|7827,7835|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|7827,7835|false|false|false|C5237010|Expression Negative|negative
Anatomy|Cell|Hospital Course|7836,7851|false|false|false|C0334227|Tumor cells, malignant|malignant cells
Anatomy|Cell|Hospital Course|7846,7851|false|false|false|C0007634|Cells|cells
Finding|Idea or Concept|Hospital Course|7856,7864|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|7856,7867|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7868,7877|false|false|false|C0229889|Lymphatic vessel|lymphatic
Finding|Finding|Hospital Course|7868,7877|true|false|false|C0740775|Lymphatic problem|lymphatic
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7881,7888|false|false|false|C0042027|Urinary tract|urinary
Drug|Substance|Hospital Course|7890,7895|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|7890,7895|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Finding|Hospital Course|7902,7905|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|7902,7905|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|Hospital Course|7906,7911|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|7906,7911|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|Hospital Course|7948,7953|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|7948,7953|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|7955,7965|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|7970,7980|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Drug|Substance|Hospital Course|8000,8005|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|8000,8005|false|false|false|C1546604|Drain Specimen Code|drain
Disorder|Disease or Syndrome|Hospital Course|8010,8015|false|false|false|C1410088|Still|still
Finding|Body Substance|Hospital Course|8026,8046|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|Hospital Course|8041,8046|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8041,8046|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Sign or Symptom|Hospital Course|8107,8113|false|false|false|C0015967|Fever|fevers
Disorder|Disease or Syndrome|Hospital Course|8115,8127|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|8115,8127|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Drug|Substance|Hospital Course|8132,8137|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8132,8137|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Antibiotic|Hospital Course|8174,8185|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Conceptual Entity|Hospital Course|8216,8224|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|Hospital Course|8231,8240|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|Hospital Course|8231,8240|false|false|false|C1120106|ertapenem|ertapenem
Finding|Body Substance|Hospital Course|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8244,8253|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8244,8253|false|false|false|C0030685|Patient Discharge|discharge
Finding|Functional Concept|Hospital Course|8278,8284|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|8278,8284|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Disorder|Neoplastic Process|Hospital Course|8285,8288|false|false|false|C0334463|Malignant Fibrous Histiocytoma|ups
Finding|Gene or Genome|Hospital Course|8285,8288|false|false|false|C1415597|HMBS gene|ups
Finding|Finding|Hospital Course|8293,8300|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|8293,8300|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Idea or Concept|Hospital Course|8321,8333|false|false|false|C1548597|Marketing basis - Transitional|transitional
Finding|Intellectual Product|Hospital Course|8346,8351|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8375,8381|false|false|false|C0030797|Pelvis|Pelvic
Drug|Substance|Hospital Course|8382,8387|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8382,8387|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Body Substance|Hospital Course|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|8401,8408|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Disorder|Disease or Syndrome|Hospital Course|8426,8434|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Drug|Substance|Hospital Course|8436,8441|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|8436,8441|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Body Substance|Hospital Course|8454,8474|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|Hospital Course|8469,8474|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8469,8474|false|false|false|C1546638|Fluid Specimen Code|fluid
Attribute|Clinical Attribute|Hospital Course|8476,8486|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|Hospital Course|8476,8486|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|Hospital Course|8479,8486|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|8479,8486|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|8479,8486|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8487,8493|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|8487,8493|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|8487,8493|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|8487,8493|false|false|false|C0812455|Pelvis problem|pelvis
Finding|Functional Concept|Hospital Course|8514,8518|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Substance|Hospital Course|8519,8524|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8519,8524|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|8525,8535|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Mental Process|Hospital Course|8541,8549|false|false|false|C0679006|Decision|decision
Event|Activity|Hospital Course|8563,8568|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|8563,8568|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|8563,8568|false|false|false|C1533810||place
Drug|Substance|Hospital Course|8571,8576|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|8571,8576|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|Hospital Course|8590,8595|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8590,8595|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Classification|Hospital Course|8600,8608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|8600,8608|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|8600,8608|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|8600,8612|false|false|false|C0205160|Negative|negative for
Anatomy|Cell|Hospital Course|8624,8629|false|false|false|C0007634|Cells|cells
Drug|Substance|Hospital Course|8635,8640|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8635,8640|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Biologically Active Substance|Hospital Course|8654,8667|false|false|false|C0041004|Triglycerides|triglycerides
Drug|Organic Chemical|Hospital Course|8654,8667|false|false|false|C0041004|Triglycerides|triglycerides
Finding|Physiologic Function|Hospital Course|8654,8667|false|false|false|C4554056|Triglycerides metabolic function|triglycerides
Procedure|Laboratory Procedure|Hospital Course|8654,8667|false|false|false|C0202236|Triglycerides measurement|triglycerides
Drug|Substance|Hospital Course|8688,8693|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8688,8693|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|8694,8704|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|8694,8704|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|8694,8704|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|8694,8704|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Body Substance|Hospital Course|8716,8721|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Functional Concept|Hospital Course|8716,8721|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Finding|Intellectual Product|Hospital Course|8716,8721|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|urine
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8726,8735|false|false|false|C0229889|Lymphatic vessel|lymphatic
Finding|Finding|Hospital Course|8726,8735|false|false|false|C0740775|Lymphatic problem|lymphatic
Drug|Substance|Hospital Course|8736,8741|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8736,8741|false|false|false|C1546638|Fluid Specimen Code|fluid
Drug|Substance|Hospital Course|8743,8748|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|Fluid
Finding|Intellectual Product|Hospital Course|8743,8748|false|false|false|C1546638|Fluid Specimen Code|Fluid
Drug|Biomedical or Dental Material|Hospital Course|8750,8757|false|false|false|C1706355|Culture Dose Form|culture
Finding|Functional Concept|Hospital Course|8750,8757|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Finding|Idea or Concept|Hospital Course|8750,8757|false|false|false|C0010453;C0220814|Cultural aspects;Culture (Anthropological)|culture
Procedure|Laboratory Procedure|Hospital Course|8750,8757|false|false|false|C0430400;C2242979|Laboratory culture;Microbial culture (procedure)|culture
Finding|Classification|Hospital Course|8762,8770|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|8762,8770|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|8762,8770|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|8762,8774|false|false|false|C0205160|Negative|negative for
Finding|Functional Concept|Hospital Course|8775,8783|false|false|false|C1510439|bacteria aspects|bacteria
Finding|Intellectual Product|Hospital Course|8788,8796|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Finding|Finding|Hospital Course|8797,8804|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|8797,8804|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Finding|Hospital Course|8810,8813|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|8810,8813|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Substance|Hospital Course|8825,8830|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8825,8830|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|8831,8841|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|8846,8856|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Drug|Substance|Hospital Course|8876,8881|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|8876,8881|false|false|false|C1546604|Drain Specimen Code|drain
Drug|Substance|Hospital Course|8912,8917|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8912,8917|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|8918,8928|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Drug|Substance|Hospital Course|8949,8954|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|8949,8954|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Body Substance|Hospital Course|8967,8987|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|Hospital Course|8982,8987|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|8982,8987|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Body Substance|Hospital Course|9012,9032|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|Hospital Course|9027,9032|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9027,9032|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Location or Region|Hospital Course|9042,9047|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|9042,9047|false|false|false|C2003888|Lower (action)|lower
Event|Activity|Hospital Course|9048,9052|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|9048,9052|false|false|false|C1549480|Amount type - Rate|rate
Procedure|Health Care Activity|Hospital Course|9068,9077|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Substance|Hospital Course|9083,9088|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|9083,9088|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Functional Concept|Hospital Course|9093,9097|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Activity|Hospital Course|9101,9106|false|false|false|C1882509|put - instruction imperative|place
Finding|Functional Concept|Hospital Course|9101,9106|false|false|false|C1704765|Place - dosing instruction imperative|place
Procedure|Health Care Activity|Hospital Course|9101,9106|false|false|false|C1533810||place
Drug|Substance|Hospital Course|9114,9119|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9114,9119|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|9121,9131|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|9121,9131|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|9121,9131|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|9121,9131|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Finding|Hospital Course|9135,9142|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|9135,9142|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Intellectual Product|Hospital Course|9151,9161|false|false|false|C4554154|Completely - dosing instruction fragment|completely
Finding|Finding|Hospital Course|9162,9171|false|true|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Finding|Functional Concept|Hospital Course|9162,9171|false|true|false|C0344329;C0392748|Collapse (finding);Collapsed|collapsed
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9173,9176|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9173,9176|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9173,9176|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9173,9176|false|false|false|C1332410|BID gene|BID
Finding|Idea or Concept|Hospital Course|9182,9190|false|true|false|C0010453|Culture (Anthropological)|cultures
Drug|Substance|Hospital Course|9214,9219|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9214,9219|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|9220,9230|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Cell or Molecular Dysfunction|Hospital Course|9242,9250|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|9242,9250|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|9242,9250|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|9242,9254|false|false|false|C1446409|Positive|positive for
Finding|Finding|Hospital Course|9255,9259|false|false|false|C2355591|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|MSSA
Drug|Organic Chemical|Hospital Course|9289,9292|false|true|false|C0939812|Ruta graveolens preparation|rue
Drug|Pharmacologic Substance|Hospital Course|9289,9292|false|true|false|C0939812|Ruta graveolens preparation|rue
Finding|Functional Concept|Hospital Course|9294,9309|false|false|false|C1512911|Intraabdominal Route of Administration|intra-abdominal
Disorder|Disease or Syndrome|Hospital Course|9294,9319|false|false|false|C1112209|Abdominal Infection|intra-abdominal infection
Disorder|Disease or Syndrome|Hospital Course|9310,9319|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|9310,9319|false|false|false|C3714514|Infection|infection
Finding|Body Substance|Hospital Course|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9332,9339|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|9346,9351|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|9346,9351|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Disorder|Disease or Syndrome|Hospital Course|9366,9378|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|9366,9378|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Finding|Conceptual Entity|Hospital Course|9404,9412|false|false|false|C2827424|Spectrum|spectrum
Drug|Antibiotic|Hospital Course|9413,9424|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Drug|Organic Chemical|Hospital Course|9448,9454|false|false|false|C0699678|Flagyl|flagyl
Drug|Pharmacologic Substance|Hospital Course|9448,9454|false|false|false|C0699678|Flagyl|flagyl
Drug|Antibiotic|Hospital Course|9492,9497|false|false|false|C0250482|Zosyn|zosyn
Drug|Organic Chemical|Hospital Course|9492,9497|false|false|false|C0250482|Zosyn|zosyn
Finding|Body Substance|Hospital Course|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9502,9511|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9502,9511|false|false|false|C0030685|Patient Discharge|discharge
Drug|Antibiotic|Hospital Course|9528,9537|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|Hospital Course|9528,9537|false|false|false|C1120106|ertapenem|ertapenem
Finding|Idea or Concept|Hospital Course|9570,9575|false|false|false|C1546485|Diagnosis Type - Final|final
Finding|Conceptual Entity|Hospital Course|9586,9595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|9586,9595|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|9586,9595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9586,9595|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Drug|Substance|Hospital Course|9616,9621|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|9616,9621|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|9623,9633|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|9634,9641|false|false|false|C0392747|Changing|changes
Finding|Functional Concept|Hospital Course|9645,9651|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Finding|Finding|Hospital Course|9652,9659|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|9652,9659|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Finding|Classification|Hospital Course|9663,9673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|9663,9673|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|Hospital Course|9674,9679|false|false|false|C1874451|Basis|basis
Finding|Functional Concept|Hospital Course|9674,9679|false|false|false|C1527178|Basis - conceptual entity|basis
Finding|Finding|Hospital Course|9700,9708|false|false|false|C0277797|Apyrexial|afebrile
Disorder|Disease or Syndrome|Hospital Course|9714,9726|false|false|false|C0023518|Leukocytosis|leukocytosis
Finding|Finding|Hospital Course|9714,9726|false|false|false|C0750426|Blood leukocyte number above reference range|leukocytosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9740,9749|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Hospital Course|9740,9749|false|false|false|C2707265||Pulmonary
Finding|Finding|Hospital Course|9740,9749|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Finding|Pathologic Function|Hospital Course|9740,9758|false|false|false|C0034065|Pulmonary Embolism|Pulmonary embolism
Finding|Finding|Hospital Course|9750,9758|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|Hospital Course|9750,9758|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Finding|Hospital Course|9760,9766|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|9760,9766|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Mental Process|Hospital Course|9784,9791|false|false|false|C0542559|contextual factors|setting
Anatomy|Body Location or Region|Hospital Course|9827,9830|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|9827,9830|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|9827,9830|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Organic Chemical|Hospital Course|9850,9857|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9850,9857|false|false|false|C0728963|Lovenox|lovenox
Drug|Biologically Active Substance|Hospital Course|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|9885,9892|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9893,9896|false|false|false|C0017040|Gamma-glutamyl transferase|ggt
Drug|Enzyme|Hospital Course|9893,9896|false|false|false|C0017040|Gamma-glutamyl transferase|ggt
Finding|Gene or Genome|Hospital Course|9893,9896|false|false|false|C1415053;C1415054|GGT1 gene;GGT2P gene|ggt
Procedure|Laboratory Procedure|Hospital Course|9893,9896|false|false|false|C0202035|Gamma glutamyl transferase measurement|ggt
Finding|Functional Concept|Hospital Course|9915,9925|false|false|false|C0025664;C2700391|Methods aspects;Procedure (set of actions)|procedures
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9915,9925|false|false|false|C0184661|Interventional procedure|procedures
Drug|Organic Chemical|Hospital Course|9956,9963|false|false|false|C0728963|Lovenox|lovenox
Drug|Pharmacologic Substance|Hospital Course|9956,9963|false|false|false|C0728963|Lovenox|lovenox
Anatomy|Body Location or Region|Hospital Course|9973,9978|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|9973,9978|false|false|false|C2003888|Lower (action)|lower
Attribute|Clinical Attribute|Hospital Course|9988,9994|false|false|false|C0944911||weight
Finding|Finding|Hospital Course|9988,9994|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|9988,9994|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|9988,9994|false|false|false|C1305866|Weighing patient|weight
Finding|Body Substance|Hospital Course|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10021,10030|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10021,10030|false|false|false|C0030685|Patient Discharge|discharge
Finding|Intellectual Product|Hospital Course|10035,10040|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Injury or Poisoning|Hospital Course|10035,10053|false|false|false|C2609414|Acute kidney injury|Acute renal injury
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10041,10046|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|10041,10046|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Injury or Poisoning|Hospital Course|10041,10053|false|false|false|C0160420|Injury of kidney|renal injury
Disorder|Injury or Poisoning|Hospital Course|10047,10053|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Disorder|Disease or Syndrome|Hospital Course|10055,10058|false|false|false|C5239292|Solitary Cutaneous Reticulohistiocytosis|SCr
Finding|Finding|Hospital Course|10055,10058|false|false|false|C1539487;C4050416|FBXL20 gene;Stringent Complete Response|SCr
Finding|Gene or Genome|Hospital Course|10055,10058|false|false|false|C1539487;C4050416|FBXL20 gene;Stringent Complete Response|SCr
Drug|Biomedical or Dental Material|Hospital Course|10092,10100|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|10092,10100|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|10136,10142|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10136,10142|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|10159,10167|false|false|false|C0042075|Urologic Diseases|uropathy
Finding|Gene or Genome|Hospital Course|10172,10177|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|Hospital Course|10185,10190|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|10185,10190|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Idea or Concept|Hospital Course|10241,10249|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Hospital Course|10260,10265|false|false|false|C1546485|Diagnosis Type - Final|final
Disorder|Disease or Syndrome|Hospital Course|10278,10292|false|false|false|C0020295|Hydronephrosis|Hydronephrosis
Finding|Intellectual Product|Hospital Course|10321,10329|false|false|false|C1552654|Parameterized Data Type - Interval|interval
Finding|Finding|Hospital Course|10330,10337|false|false|false|C0740845|Imaging problem|imaging
Procedure|Diagnostic Procedure|Hospital Course|10330,10337|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|imaging
Procedure|Research Activity|Hospital Course|10350,10357|false|false|false|C0947630|Scientific Study|studies
Finding|Body Substance|Hospital Course|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10365,10372|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|Hospital Course|10375,10378|false|false|false|C1114365||age
Drug|Biologically Active Substance|Hospital Course|10375,10378|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Hospital Course|10375,10378|false|false|false|C0162574|Glycation End Products, Advanced|age
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10389,10396|false|false|false|C0042027|Urinary tract|urinary
Finding|Conceptual Entity|Hospital Course|10398,10404|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Hospital Course|10398,10404|false|false|false|C3251815|Measurement of fluid output|output
Drug|Biologically Active Substance|Hospital Course|10415,10425|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|10415,10425|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|Hospital Course|10415,10425|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|10415,10425|false|false|false|C0201975|Creatinine measurement|creatinine
Phenomenon|Biologic Function|Hospital Course|10415,10435|false|false|false|C0812399|Creatinine clearance|creatinine clearance
Procedure|Laboratory Procedure|Hospital Course|10415,10435|false|false|false|C0373595|Creatinine renal clearance measurement|creatinine clearance
Attribute|Clinical Attribute|Hospital Course|10426,10435|false|false|false|C1382187|Clearance of substance|clearance
Phenomenon|Natural Phenomenon or Process|Hospital Course|10426,10435|false|false|false|C2825073|Clearance [PK]|clearance
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10426,10435|false|false|false|C4554548|Clearance procedure|clearance
Finding|Idea or Concept|Hospital Course|10444,10455|false|false|false|C0750502|Significant|significant
Drug|Inorganic Chemical|Hospital Course|10457,10468|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Drug|Pharmacologic Substance|Hospital Course|10457,10468|false|false|false|C0013832;C3536863|Electrolyte [EPC];Electrolytes|electrolyte
Disorder|Congenital Abnormality|Hospital Course|10469,10482|false|false|false|C0000768|Congenital Abnormality|abnormalities
Finding|Functional Concept|Hospital Course|10469,10482|false|false|false|C0000769|teratologic|abnormalities
Finding|Body Substance|Hospital Course|10484,10491|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10484,10491|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10484,10491|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Finding|Hospital Course|10492,10498|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10492,10498|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Procedure|Health Care Activity|Hospital Course|10537,10549|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10537,10549|false|false|false|C0184661;C0886296;C1273869|Intervention regimes;Interventional procedure;Nursing interventions|intervention
Finding|Finding|Hospital Course|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|10558,10562|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|Hospital Course|10564,10567|false|false|false|C0449201|PER (body structure)|Per
Disorder|Disease or Syndrome|Hospital Course|10564,10567|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Per
Finding|Functional Concept|Hospital Course|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Gene or Genome|Hospital Course|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Intellectual Product|Hospital Course|10564,10567|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Procedure|Health Care Activity|Hospital Course|10577,10584|false|false|false|C0009818|Consultation|consult
Finding|Intellectual Product|Hospital Course|10593,10599|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Body Substance|Hospital Course|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|10604,10613|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|10604,10613|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|10618,10629|false|false|false|C0034866|Recommendation|recommended
Finding|Classification|Hospital Course|10631,10641|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|10631,10641|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Procedure|Health Care Activity|Hospital Course|10650,10658|false|false|false|C1522577|follow-up|followup
Disorder|Disease or Syndrome|Hospital Course|10663,10669|false|false|false|C0002871|Anemia|Anemia
Finding|Finding|Hospital Course|10671,10677|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10671,10677|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|Hospital Course|10680,10691|false|true|false|C3811910|combination - answer to question|combination
Disorder|Disease or Syndrome|Hospital Course|10695,10701|false|false|false|C0002871|Anemia|anemia
Disorder|Disease or Syndrome|Hospital Course|10695,10725|false|false|false|C0002873|Anemia of chronic disease|anemia of chronic inflammation
Finding|Intellectual Product|Hospital Course|10705,10712|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|10705,10712|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Pathologic Function|Hospital Course|10705,10725|false|false|false|C0021376|Chronic inflammation|chronic inflammation
Finding|Pathologic Function|Hospital Course|10713,10725|false|false|false|C0021368|Inflammation|inflammation
Finding|Intellectual Product|Hospital Course|10731,10736|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Hospital Course|10731,10747|false|false|false|C0333276|Acute hemorrhage|acute blood loss
Disorder|Disease or Syndrome|Hospital Course|10737,10742|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|10737,10742|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|10737,10747|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|Hospital Course|10737,10747|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Finding|Hospital Course|10743,10747|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Hospital Course|10755,10763|false|false|false|C0751437|Adenohypophyseal Diseases|anterior
Anatomy|Body Location or Region|Hospital Course|10764,10773|false|false|false|C0000726|Abdomen|abdominal
Finding|Finding|Hospital Course|10764,10779|false|false|false|C2266645|abdominal drain in place|abdominal drain
Drug|Substance|Hospital Course|10774,10779|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Hospital Course|10774,10779|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Body Substance|Hospital Course|10789,10809|false|false|false|C4518404|Serosanguinous fluid|serosanguinous fluid
Drug|Substance|Hospital Course|10804,10809|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|10804,10809|false|false|false|C1546638|Fluid Specimen Code|fluid
Lab|Laboratory or Test Result|Hospital Course|10811,10815|false|false|false|C0587081|Laboratory test finding|Labs
Finding|Idea or Concept|Hospital Course|10820,10830|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|10820,10835|false|false|false|C0332290|Consistent with|consistent with
Finding|Cell Function|Hospital Course|10836,10845|false|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Finding|Hospital Course|10836,10845|false|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Pathologic Function|Hospital Course|10836,10845|false|true|false|C0019054;C1553188;C2937287;C2945560|Hemolysis (biological function);Hemolysis (disorder);Hemolysis (finding)|hemolysis
Finding|Finding|Hospital Course|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|Hospital Course|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|Hospital Course|10890,10898|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Body Substance|Hospital Course|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10900,10907|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10929,10932|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|10929,10932|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Hospital Course|10929,10932|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|10929,10932|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Pathologic Function|Hospital Course|10944,10947|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10944,10947|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Finding|Idea or Concept|Hospital Course|10952,10966|false|false|false|C0034866|Recommendation|recommendation
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10982,10985|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Hospital Course|10982,10985|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Hospital Course|10982,10985|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Hospital Course|10982,10985|false|false|false|C0019029|Hemoglobin concentration|Hgb
Finding|Body Substance|Hospital Course|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10991,10998|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11032,11038|false|false|false|C1550462|Observation Interpretation - better|better
Disorder|Disease or Syndrome|Hospital Course|11051,11056|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|11051,11056|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|11068,11079|false|false|false|C0020621|Hypokalemia|Hypokalemia
Anatomy|Body Space or Junction|Hospital Course|11119,11123|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|11119,11123|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|11119,11123|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|11119,11123|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Inorganic Chemical|Hospital Course|11124,11127|false|false|false|C0032825|potassium chloride|KCl
Drug|Pharmacologic Substance|Hospital Course|11124,11127|false|false|false|C0032825|potassium chloride|KCl
Finding|Gene or Genome|Hospital Course|11129,11132|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Intellectual Product|Hospital Course|11136,11143|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|11136,11143|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Finding|Finding|Hospital Course|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|11178,11182|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Disorder|Neoplastic Process|Hospital Course|11178,11209|false|false|false|C5556496|Urothelial Carcinoma, High Grade|high-grade urothelial carcinoma
Finding|Classification|Hospital Course|11183,11188|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Hospital Course|11183,11188|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|Hospital Course|11189,11209|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|Hospital Course|11200,11209|false|false|false|C0007097|Carcinoma|carcinoma
Attribute|Clinical Attribute|Hospital Course|11225,11229|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11231,11241|false|false|false|C0225358;C4551532|Bladder Detrusor Muscle;Muscle layer|muscularis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11231,11249|false|false|false|C0225358|Bladder Detrusor Muscle|muscularis propria
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11254,11264|false|false|false|C0010651|Cystectomy|cystectomy
Finding|Finding|Hospital Course|11266,11278|false|false|false|C1548863|Consent Type - Hysterectomy|hysterectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11266,11278|false|false|false|C0020699|Hysterectomy|hysterectomy
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Hazardous or Poisonous Substance|Hospital Course|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Drug|Pharmacologic Substance|Hospital Course|11284,11287|false|false|false|C0054252|Buthionine Sulfoximine|BSO
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11297,11302|false|false|false|C0020885|ileum|ileal
Disorder|Acquired Abnormality|Hospital Course|11297,11310|false|false|false|C0441253|Structure of ileal conduit|ileal conduit
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11297,11310|false|false|false|C0348002|Ileal conduit procedure|ileal conduit
Finding|Finding|Hospital Course|11319,11333|false|false|false|C0241311|post operative (finding)|post operative
Anatomy|Body Location or Region|Hospital Course|11365,11368|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|11365,11368|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|11365,11368|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Disease or Syndrome|Hospital Course|11374,11379|false|false|false|C1258215;C4019039|Ileus;Intestinal obstruction co-occurrent and due to decreased peristalsis|ileus
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11385,11391|false|false|false|C0030797|Pelvis|pelvic
Drug|Substance|Hospital Course|11392,11397|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|11392,11397|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Body Substance|Hospital Course|11412,11419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|11412,11419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|11412,11419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|11446,11450|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|Hospital Course|11446,11450|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|11446,11450|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|11446,11450|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11455,11460|false|false|false|C0392920;C3665472|Chemotherapy;Chemotherapy Regimen|chemo
Phenomenon|Natural Phenomenon or Process|Hospital Course|11465,11474|false|false|false|C0034519;C0851346|Electromagnetic Radiation;Radiation|radiation
Procedure|Research Activity|Hospital Course|11465,11474|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11465,11474|false|false|false|C1522449;C1524020;C1524021|Radiation Ionizing Radiotherapy;Radiation therapy (procedure);Radiotherapy Research|radiation
Procedure|Diagnostic Procedure|Hospital Course|11480,11483|false|false|false|C0032743;C0040398|Positron-Emission Tomography;Tomography, Emission-Computed|PET
Procedure|Diagnostic Procedure|Hospital Course|11480,11488|false|false|false|C0032743|Positron-Emission Tomography|PET scan
Procedure|Diagnostic Procedure|Hospital Course|11484,11488|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Finding|Hospital Course|11511,11515|false|false|false|C4321394|Foci|foci
Finding|Functional Concept|Hospital Course|11519,11529|false|false|false|C0036525;C1522484|Metastatic to;metastatic qualifier|metastatic
Disorder|Neoplastic Process|Hospital Course|11519,11537|false|false|false|C0027627;C2939419;C2939420|Metastatic Neoplasm;Metastatic malignant neoplasm;Neoplasm Metastasis|metastatic disease
Finding|Finding|Hospital Course|11519,11537|false|false|false|C1513183|Metastatic Lesion|metastatic disease
Disorder|Disease or Syndrome|Hospital Course|11530,11537|false|false|false|C0012634|Disease|disease
Anatomy|Body Location or Region|Hospital Course|11545,11549|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11545,11549|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|11545,11549|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|11545,11549|false|false|false|C0740941|Lung Problem|lung
Anatomy|Tissue|Hospital Course|11555,11565|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|Hospital Course|11555,11565|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Finding|Body Substance|Hospital Course|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11571,11578|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|Hospital Course|11581,11584|false|false|false|C1420310|SON gene|son
Finding|Intellectual Product|Hospital Course|11606,11612|false|false|false|C2348314|Doctor - Title|doctor
Event|Occupational Activity|Hospital Course|11617,11621|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|11617,11624|false|false|false|C0750430|Work-up|work up
Anatomy|Body Location or Region|Hospital Course|11629,11633|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11629,11633|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|11629,11633|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|11629,11633|false|false|false|C0740941|Lung Problem|lung
Finding|Finding|Hospital Course|11629,11638|false|false|false|C0149726|Lung mass|lung mass
Finding|Finding|Hospital Course|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|11634,11638|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Idea or Concept|Hospital Course|11650,11657|false|false|false|C0549178|Continuous|ongoing
Finding|Social Behavior|Hospital Course|11658,11668|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11658,11668|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|Hospital Course|11675,11685|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|11675,11685|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Pathologic Function|Hospital Course|11686,11689|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11686,11689|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Disorder|Disease or Syndrome|Hospital Course|11711,11715|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Finding|Gene or Genome|Hospital Course|11711,11715|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Finding|Finding|Hospital Course|11735,11742|false|false|false|C0221198|Lesion|lesions
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11747,11753|false|false|false|C0006141|Breast|Breast
Disorder|Neoplastic Process|Hospital Course|11747,11753|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|Breast
Finding|Finding|Hospital Course|11747,11753|false|false|false|C0567499|Breast problem|Breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11747,11753|false|false|false|C0191838|Procedures on breast|Breast
Finding|Finding|Hospital Course|11747,11758|false|false|false|C0024103|Mass in breast|Breast mass
Finding|Finding|Hospital Course|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|11754,11758|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Finding|Hospital Course|11763,11772|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|Hospital Course|11763,11772|false|false|false|C0024671|Mammography|mammogram
Finding|Intellectual Product|Hospital Course|11781,11788|false|false|false|C1511314|Breast Imaging Reporting and Data System|BI-RADS
Finding|Intellectual Product|Hospital Course|11781,11790|false|false|false|C5960924|Breast Imaging-Reporting and Data System Assessment Category 5|BI-RADS 5
Drug|Biomedical or Dental Material|Hospital Course|11792,11797|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|Solid
Drug|Substance|Hospital Course|11792,11797|false|false|false|C0302909;C1378566|Solid Dose Form;solid substance|Solid
Finding|Finding|Hospital Course|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|11798,11802|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11815,11820|false|false|false|C1743089|CLOCK protein, human|clock
Drug|Enzyme|Hospital Course|11815,11820|false|false|false|C1743089|CLOCK protein, human|clock
Finding|Gene or Genome|Hospital Course|11815,11820|false|false|false|C1413503|CLOCK gene|clock
Finding|Functional Concept|Hospital Course|11821,11825|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11821,11832|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11826,11832|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|11826,11832|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|11826,11832|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11826,11832|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Hospital Course|11860,11885|false|false|false|C4050405|Suspicious for Malignancy|suspicious for malignancy
Disorder|Neoplastic Process|Hospital Course|11875,11885|false|true|false|C0006826;C1306459|Malignant Neoplasms;Primary malignant neoplasm|malignancy
Finding|Body Substance|Hospital Course|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11891,11898|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Gene or Genome|Hospital Course|11901,11904|false|false|false|C1420310|SON gene|son
Finding|Intellectual Product|Hospital Course|11922,11928|false|false|false|C2348314|Doctor - Title|doctor
Finding|Finding|Hospital Course|11948,11951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|11948,11951|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11952,11958|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|11952,11958|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|11952,11958|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11952,11958|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Hospital Course|11952,11963|false|false|false|C0024103|Mass in breast|breast mass
Finding|Finding|Hospital Course|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|11959,11963|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Idea or Concept|Hospital Course|11982,11989|false|false|false|C0549178|Continuous|ongoing
Finding|Social Behavior|Hospital Course|11990,12000|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11990,12000|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Intellectual Product|Hospital Course|12021,12027|false|false|true|C2348314|Doctor - Title|doctor
Finding|Classification|Hospital Course|12032,12042|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12032,12042|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|12058,12062|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Finding|Functional Concept|Hospital Course|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|Hospital Course|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|Hospital Course|12058,12062|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Drug|Organic Chemical|Hospital Course|12092,12104|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12092,12104|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Functional Concept|Hospital Course|12113,12120|true|false|false|C0392747|Changing|changes
Finding|Idea or Concept|Hospital Course|12122,12130|false|false|false|C0750591|consider|Consider
Finding|Idea or Concept|Hospital Course|12132,12142|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|12132,12142|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Drug|Inorganic Chemical|Hospital Course|12153,12161|false|false|false|C0723457|Stop brand of fluoride|stopping
Drug|Pharmacologic Substance|Hospital Course|12153,12161|false|false|false|C0723457|Stop brand of fluoride|stopping
Drug|Organic Chemical|Hospital Course|12162,12174|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|12162,12174|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Classification|Hospital Course|12178,12188|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|12178,12188|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Pharmacologic Substance|Hospital Course|12189,12194|false|false|false|C1874451|Basis|basis
Finding|Functional Concept|Hospital Course|12189,12194|false|false|false|C1527178|Basis - conceptual entity|basis
Disorder|Disease or Syndrome|Hospital Course|12200,12214|false|false|false|C0020676|Hypothyroidism|Hypothyroidism
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12226,12239|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Hormone|Hospital Course|12226,12239|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Organic Chemical|Hospital Course|12226,12239|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Drug|Pharmacologic Substance|Hospital Course|12226,12239|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|levothyroxine
Finding|Functional Concept|Hospital Course|12248,12255|true|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|Hospital Course|12264,12267|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Finding|Gene or Genome|Hospital Course|12264,12267|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Finding|Gene or Genome|Hospital Course|12279,12282|false|false|false|C1420310|SON gene|son
Attribute|Clinical Attribute|Hospital Course|12288,12297|false|false|false|C0804815||physician
Event|Occupational Activity|Hospital Course|12304,12308|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|12304,12308|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|Hospital Course|12304,12315|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|Hospital Course|12309,12315|false|false|false|C5889824||status
Finding|Idea or Concept|Hospital Course|12309,12315|false|false|false|C1546481|What subject filter - Status|status
Event|Occupational Activity|Hospital Course|12322,12326|false|false|false|C0009219|Coding|code
Finding|Intellectual Product|Hospital Course|12322,12326|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|code
Finding|Body Substance|Hospital Course|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|12343,12350|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|12360,12372|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Disorder|Disease or Syndrome|Hospital Course|12416,12426|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Hospital Course|12416,12434|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|Hospital Course|12427,12434|false|false|false|C0012634|Disease|disease
Finding|Functional Concept|Hospital Course|12435,12441|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|Hospital Course|12435,12441|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|Hospital Course|12435,12444|false|false|false|C0589120|Follow-up status|follow up
Procedure|Health Care Activity|Hospital Course|12435,12444|false|false|false|C1522577|follow-up|follow up
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12511,12514|false|false|false|C1137947|SET protein, human|set
Drug|Biologically Active Substance|Hospital Course|12511,12514|false|false|false|C1137947|SET protein, human|set
Finding|Conceptual Entity|Hospital Course|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Functional Concept|Hospital Course|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Gene or Genome|Hospital Course|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Idea or Concept|Hospital Course|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Finding|Mental Process|Hospital Course|12511,12514|false|false|false|C0036849;C1366517;C1442518;C1552652;C1705195|Parameterized Data Type - Set;SET gene;Set (Psychology);Set scale;set (group)|set
Event|Activity|Hospital Course|12511,12517|false|false|false|C1521827|Preparation|set up
Event|Activity|Hospital Course|12521,12532|false|false|false|C0003629|Appointments|appointment
Event|Activity|Hospital Course|12541,12552|false|false|false|C0003629|Appointments|appointment
Attribute|Clinical Attribute|Hospital Course|12576,12586|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|Hospital Course|12576,12586|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|Hospital Course|12579,12586|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|12579,12586|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|12579,12586|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12587,12593|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|12587,12593|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|12587,12593|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|12587,12593|false|false|false|C0812455|Pelvis problem|pelvis
Attribute|Clinical Attribute|Hospital Course|12649,12659|false|false|false|C1644645||CT abdomen
Procedure|Diagnostic Procedure|Hospital Course|12649,12659|false|false|false|C0412620|CT of abdomen|CT abdomen
Anatomy|Body Location or Region|Hospital Course|12652,12659|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|Hospital Course|12652,12659|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|Hospital Course|12652,12659|false|false|false|C0941288|Abdomen problem|abdomen
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12662,12668|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Hospital Course|12662,12668|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Hospital Course|12662,12668|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Hospital Course|12662,12668|false|false|false|C0812455|Pelvis problem|pelvis
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|12675,12683|false|false|false|C0009924|Contrast Media|contrast
Finding|Intellectual Product|Hospital Course|12691,12695|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Gene or Genome|Hospital Course|12729,12732|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Finding|Intellectual Product|Hospital Course|12729,12732|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|lab
Anatomy|Cell Component|Hospital Course|12757,12760|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Procedure|Laboratory Procedure|Hospital Course|12757,12760|false|false|false|C0009555|Complete Blood Count|CBC
Finding|Idea or Concept|Hospital Course|12767,12779|false|false|false|C1549478|Amount type - Differential|differential
Drug|Biologically Active Substance|Hospital Course|12781,12784|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|Hospital Course|12781,12784|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Procedure|Laboratory Procedure|Hospital Course|12781,12784|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Anatomy|Body Space or Junction|Hospital Course|12790,12793|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|Hospital Course|12790,12793|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|Hospital Course|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|Hospital Course|12790,12793|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Finding|Gene or Genome|Hospital Course|12790,12793|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Disorder|Neoplastic Process|Hospital Course|12795,12798|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12795,12798|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|Hospital Course|12795,12798|false|false|false|C0001899|Alanine Transaminase|ALT
Finding|Gene or Genome|Hospital Course|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|Hospital Course|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|Hospital Course|12795,12798|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12795,12798|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12804,12807|false|false|false|C1663627|ALK protein, human|ALK
Drug|Enzyme|Hospital Course|12804,12807|false|false|false|C1663627|ALK protein, human|ALK
Finding|Gene or Genome|Hospital Course|12804,12807|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Finding|Receptor|Hospital Course|12804,12807|false|false|false|C1332080;C1663627;C1704943|ALK gene;ALK protein, human;ALK wt Allele|ALK
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12804,12812|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Drug|Enzyme|Hospital Course|12804,12812|false|false|false|C0002059|Alkaline Phosphatase|ALK PHOS
Procedure|Laboratory Procedure|Hospital Course|12804,12812|false|false|false|C0201850|Alkaline phosphatase measurement|ALK PHOS
Finding|Gene or Genome|Hospital Course|12818,12821|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Finding|Intellectual Product|Hospital Course|12818,12821|false|false|false|C1825793;C5420098;C5420670|AML Lab Table;EWS Lab Table;LAT2 gene|LAB
Event|Activity|Hospital Course|12822,12830|false|false|false|C1272683||REQUESTS
Finding|Idea or Concept|Hospital Course|12842,12851|false|false|false|C1552657|Annotated - ParameterizedDataType|ANNOTATED
Finding|Idea or Concept|Hospital Course|12879,12882|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Intellectual Product|Hospital Course|12879,12882|false|false|false|C1547563;C1549619|Authorization Mode - Fax;Fax Number|FAX
Finding|Finding|Hospital Course|12896,12904|false|false|false|C0332149|Possible|possible
Drug|Antibiotic|Hospital Course|12918,12927|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|Hospital Course|12918,12927|false|false|false|C1120106|ertapenem|ertapenem
Finding|Finding|Hospital Course|12937,12941|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Hospital Course|12937,12941|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Hospital Course|12937,12941|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Daily or Recreational Activity|Hospital Course|12977,12993|false|false|false|C0871707|daily activities|daily activities
Event|Activity|Hospital Course|12983,12993|false|false|false|C0441655|Activities|activities
Finding|Finding|Hospital Course|12983,12993|false|false|false|C2239122|activities (history)|activities
Drug|Antibiotic|Hospital Course|13031,13040|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|Hospital Course|13031,13040|false|false|false|C1120106|ertapenem|ertapenem
Finding|Idea or Concept|Hospital Course|13064,13069|false|false|false|C1546485|Diagnosis Type - Final|final
Finding|Conceptual Entity|Hospital Course|13070,13079|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Hospital Course|13070,13079|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Hospital Course|13070,13079|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13070,13079|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Disorder|Disease or Syndrome|Hospital Course|13106,13116|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Hospital Course|13106,13124|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|Hospital Course|13117,13124|false|false|false|C0012634|Disease|disease
Finding|Idea or Concept|Hospital Course|13146,13153|false|false|false|C0549178|Continuous|ongoing
Finding|Social Behavior|Hospital Course|13154,13164|false|false|false|C2584313|Discussion (communication)|discussion
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13154,13164|false|false|false|C0557061|Discussion (procedure)|discussion
Finding|Classification|Hospital Course|13170,13180|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|13170,13180|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|13181,13184|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|13181,13184|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Finding|Gene or Genome|Hospital Course|13181,13184|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|13181,13184|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Pathologic Function|Hospital Course|13189,13192|false|false|false|C0019080|Hemorrhage|hem
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13189,13192|false|false|false|C0280599|altretamine/etoposide/methotrexate protocol|hem
Finding|Finding|Hospital Course|13222,13225|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|13222,13225|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13226,13232|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|13226,13232|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|13226,13232|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13226,13232|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Hospital Course|13226,13239|false|false|false|C0567489|Lesion of breast|breast lesion
Finding|Finding|Hospital Course|13233,13239|false|false|false|C0221198;C1546698|Lesion|lesion
Finding|Intellectual Product|Hospital Course|13233,13239|false|false|false|C0221198;C1546698|Lesion|lesion
Anatomy|Body Location or Region|Hospital Course|13244,13248|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|13244,13248|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Hospital Course|13244,13248|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Hospital Course|13244,13248|false|false|false|C0740941|Lung Problem|lung
Anatomy|Tissue|Hospital Course|13249,13259|false|false|false|C0031153;C0230198;C4482223|Abdomen>Peritoneum;Peritoneum;Serous layer of peritoneum|peritoneum
Disorder|Neoplastic Process|Hospital Course|13249,13259|false|false|false|C0496874;C0496954|Benign neoplasm of peritoneum;Neoplasm of uncertain or unknown behavior of peritoneum|peritoneum
Finding|Finding|Hospital Course|13261,13268|false|false|false|C0221198|Lesion|lesions
Finding|Functional Concept|Hospital Course|13286,13290|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Hospital Course|13286,13294|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Drug|Organic Chemical|Hospital Course|13295,13307|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13295,13307|false|false|false|C0286651|atorvastatin|atorvastatin
Finding|Classification|Hospital Course|13322,13332|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|13322,13332|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|13385,13394|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|Hospital Course|13395,13409|false|false|false|C0020295|Hydronephrosis|hydronephrosis
Attribute|Clinical Attribute|Hospital Course|13413,13424|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|13413,13424|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|13413,13424|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|13413,13437|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|13428,13437|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|13456,13466|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|13456,13466|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|13456,13471|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|13467,13471|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|13488,13496|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|13488,13496|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|13488,13496|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|13501,13514|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|13501,13514|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|13501,13514|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|13533,13545|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|13533,13545|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|13563,13573|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|13563,13573|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|Hospital Course|13563,13580|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|13563,13580|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13574,13580|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|13574,13580|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13574,13580|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Idea or Concept|Hospital Course|13620,13624|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|Hospital Course|13625,13632|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|13625,13632|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|13625,13632|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|13633,13647|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|13633,13647|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|13648,13652|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|13657,13670|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|13657,13677|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13671,13677|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|13671,13677|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13671,13677|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|13699,13708|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|Hospital Course|13699,13708|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|Hospital Course|13730,13733|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|13734,13741|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|13734,13741|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|Hospital Course|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|13746,13755|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|13746,13755|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|13746,13767|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|13756,13767|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|13756,13767|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|13756,13767|false|false|false|C4284232|Medications|Medications
Drug|Antibiotic|Hospital Course|13773,13782|false|false|false|C1120106|ertapenem|Ertapenem
Drug|Organic Chemical|Hospital Course|13773,13782|false|false|false|C1120106|ertapenem|Ertapenem
Drug|Organic Chemical|Hospital Course|13773,13789|false|false|false|C1170745|ertapenem sodium|Ertapenem Sodium
Drug|Pharmacologic Substance|Hospital Course|13773,13789|false|false|false|C1170745|ertapenem sodium|Ertapenem Sodium
Drug|Biologically Active Substance|Hospital Course|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13783,13789|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|13783,13789|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13783,13789|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Pharmacologic Substance|Hospital Course|13800,13808|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Drug|Antibiotic|Hospital Course|13830,13839|false|false|false|C1120106|ertapenem|ertapenem
Drug|Organic Chemical|Hospital Course|13830,13839|false|false|false|C1120106|ertapenem|ertapenem
Finding|Functional Concept|Hospital Course|13879,13888|false|false|false|C0521102|Interferes with|interfere
Finding|Daily or Recreational Activity|Hospital Course|13898,13914|false|false|false|C0871707|daily activities|daily activities
Event|Activity|Hospital Course|13904,13914|false|false|false|C0441655|Activities|activities
Finding|Finding|Hospital Course|13904,13914|false|false|false|C2239122|activities (history)|activities
Drug|Food|Hospital Course|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Immunologic Factor|Hospital Course|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Pharmacologic Substance|Hospital Course|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Drug|Substance|Hospital Course|13921,13925|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|Milk
Finding|Body Substance|Hospital Course|13921,13925|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Finding|Intellectual Product|Hospital Course|13921,13925|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|Milk
Drug|Clinical Drug|Hospital Course|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|Hospital Course|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Pharmacologic Substance|Hospital Course|13921,13937|false|false|false|C0591789;C0782828|Milk of Magnesia (Brand Name);magnesium hydroxide Oral Suspension|Milk of Magnesia
Drug|Inorganic Chemical|Hospital Course|13929,13937|false|false|false|C0024477|magnesium oxide|Magnesia
Drug|Pharmacologic Substance|Hospital Course|13929,13937|false|false|false|C0024477|magnesium oxide|Magnesia
Finding|Gene or Genome|Hospital Course|13951,13954|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|Hospital Course|13955,13967|false|false|false|C0009806|Constipation|constipation
Drug|Organic Chemical|Hospital Course|13974,13984|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Pharmacologic Substance|Hospital Course|13974,13984|false|false|false|C0206460|enoxaparin|Enoxaparin
Drug|Organic Chemical|Hospital Course|13974,13991|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Pharmacologic Substance|Hospital Course|13974,13991|false|false|false|C0724579|enoxaparin sodium|Enoxaparin Sodium
Drug|Biologically Active Substance|Hospital Course|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|13985,13991|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|13985,13991|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|13985,13991|false|false|false|C0337443|Sodium measurement|Sodium
Finding|Idea or Concept|Hospital Course|14039,14043|false|false|false|C1552851|next - HtmlLinkType|Next
Finding|Idea or Concept|Hospital Course|14044,14051|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Finding|Intellectual Product|Hospital Course|14044,14051|false|false|false|C1546402;C1547137;C1547582;C1548424;C1549563;C1561591|Admission Type - Routine;Extended Priority Codes - Routine;Level of Care - Routine;Processing priority - Routine;Referral priority - Routine;Report priority - Routine|Routine
Procedure|Laboratory Procedure|Hospital Course|14044,14051|false|false|false|C1979801|Routine coag|Routine
Event|Occupational Activity|Hospital Course|14052,14066|false|false|false|C0001554|Administration occupational activities|Administration
Procedure|Therapeutic or Preventive Procedure|Hospital Course|14052,14066|false|false|false|C1533734|Administration (procedure)|Administration
Finding|Finding|Hospital Course|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Idea or Concept|Hospital Course|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Finding|Intellectual Product|Hospital Course|14068,14072|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|Time
Drug|Organic Chemical|Hospital Course|14079,14092|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|14079,14092|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|14079,14092|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Drug|Organic Chemical|Hospital Course|14113,14125|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|14113,14125|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Hormone|Hospital Course|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Organic Chemical|Hospital Course|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Pharmacologic Substance|Hospital Course|14145,14158|false|false|false|C0040165;C1881373|Synthetic Levothyroxine;levothyroxine|Levothyroxine
Drug|Amino Acid, Peptide, or Protein|Hospital Course|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Hormone|Hospital Course|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Pharmacologic Substance|Hospital Course|14145,14165|false|false|false|C0079691|levothyroxine sodium|Levothyroxine Sodium
Drug|Biologically Active Substance|Hospital Course|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|14159,14165|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|14159,14165|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|14159,14165|false|false|false|C0337443|Sodium measurement|Sodium
Drug|Organic Chemical|Hospital Course|14189,14198|false|false|false|C0024002|lorazepam|LORazepam
Drug|Pharmacologic Substance|Hospital Course|14189,14198|false|false|false|C0024002|lorazepam|LORazepam
Finding|Gene or Genome|Hospital Course|14220,14223|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|14224,14231|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Finding|Sign or Symptom|Hospital Course|14224,14231|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Body Substance|Hospital Course|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14237,14246|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14237,14246|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|14237,14258|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|14237,14258|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|14247,14258|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|14247,14258|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|14260,14268|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|14260,14268|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|14260,14273|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|14269,14273|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|14269,14273|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|14269,14273|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|14276,14284|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|14292,14301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|14292,14301|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|14292,14311|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|14302,14311|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|14302,14311|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|14302,14311|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14302,14311|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Hospital Course|14313,14330|false|false|false|C0801658||Primary diagnosis
Attribute|Clinical Attribute|Hospital Course|14321,14330|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|14321,14330|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|14321,14330|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14321,14330|false|false|false|C0011900|Diagnosis|diagnosis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14332,14338|false|false|false|C0030797|Pelvis|Pelvic
Disorder|Disease or Syndrome|Hospital Course|14332,14355|false|false|false|C1697454|Pelvic fluid collection|Pelvic fluid collection
Drug|Substance|Hospital Course|14339,14344|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Hospital Course|14339,14344|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Hospital Course|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Hospital Course|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Hospital Course|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Hospital Course|14345,14355|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|Hospital Course|14356,14365|false|false|false|C0009450|Communicable Diseases|infection
Finding|Pathologic Function|Hospital Course|14356,14365|false|false|false|C3714514|Infection|infection
Finding|Intellectual Product|Hospital Course|14372,14377|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|14379,14384|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|14379,14384|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|14379,14389|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Finding|Pathologic Function|Hospital Course|14379,14389|false|false|false|C0019080;C3163616|Blood Loss;Hemorrhage|blood loss
Disorder|Disease or Syndrome|Hospital Course|14379,14396|false|false|false|C0154286;C0154298;C0948824|Acute posthaemorrhagic anaemia;Anemia due to blood loss;Iron deficiency anemia secondary to chronic blood loss|blood loss anemia
Finding|Finding|Hospital Course|14385,14389|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Hospital Course|14390,14396|false|false|false|C0002871|Anemia|anemia
Disorder|Neoplastic Process|Hospital Course|14398,14407|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|14398,14407|false|false|false|C1522484|metastatic qualifier|Secondary
Attribute|Clinical Attribute|Hospital Course|14398,14417|false|false|false|C4255018||Secondary diagnosis
Finding|Finding|Hospital Course|14398,14417|false|false|false|C0332138|Secondary diagnosis|Secondary diagnosis
Attribute|Clinical Attribute|Hospital Course|14408,14417|false|false|false|C0945731||diagnosis
Finding|Classification|Hospital Course|14408,14417|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Finding|Functional Concept|Hospital Course|14408,14417|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|diagnosis
Procedure|Diagnostic Procedure|Hospital Course|14408,14417|false|false|false|C0011900|Diagnosis|diagnosis
Finding|Intellectual Product|Hospital Course|14419,14424|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|Hospital Course|14419,14438|false|false|false|C0022660|Kidney Failure, Acute|acute renal failure
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14425,14430|false|false|false|C0022646|Kidney|renal
Disorder|Disease or Syndrome|Hospital Course|14425,14430|false|false|false|C0042075|Urologic Diseases|renal
Disorder|Disease or Syndrome|Hospital Course|14425,14438|false|false|false|C0035078|Kidney Failure|renal failure
Disorder|Disease or Syndrome|Hospital Course|14425,14445|false|false|false|C0022660|Kidney Failure, Acute|renal failure, acute
Finding|Functional Concept|Hospital Course|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Idea or Concept|Hospital Course|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Individual Behavior|Hospital Course|14431,14438|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|failure
Finding|Intellectual Product|Hospital Course|14440,14445|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|Hospital Course|14449,14456|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|14449,14456|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|Hospital Course|14458,14464|false|false|false|C0002871|Anemia|anemia
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14473,14482|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|14473,14482|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|14473,14482|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Finding|Pathologic Function|Hospital Course|14473,14491|false|false|false|C0034065|Pulmonary Embolism|pulmonary embolism
Finding|Finding|Hospital Course|14483,14491|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Pathologic Function|Hospital Course|14483,14491|false|false|false|C0013922;C1704212|Embolism;Embolus|embolism
Finding|Finding|Hospital Course|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|14502,14506|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Classification|Hospital Course|14507,14512|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Finding|Finding|Hospital Course|14507,14512|false|false|false|C0441800;C0919553;C3244287|Grade;Histopathologic Grade;School Grade|grade
Disorder|Neoplastic Process|Hospital Course|14514,14534|false|false|false|C0007138;C2145472|Carcinoma, Transitional Cell;Urothelial Carcinoma|urothelial carcinoma
Disorder|Neoplastic Process|Hospital Course|14525,14534|false|false|false|C0007097|Carcinoma|carcinoma
Finding|Functional Concept|Hospital Course|14536,14540|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14536,14547|false|false|false|C0222601|Left breast|left breast
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|14541,14547|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Hospital Course|14541,14547|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Hospital Course|14541,14547|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Hospital Course|14541,14547|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Hospital Course|14541,14552|false|false|false|C0024103|Mass in breast|breast mass
Finding|Finding|Hospital Course|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Gene or Genome|Hospital Course|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|14548,14552|false|false|false|C0577559;C0577573;C1414542;C1546709;C2700045;C4283905|FBN1 gene;FBN1 wt Allele;Mass of body region;Mass of body structure;Morphology, Attenuation, Size, and Structure Criteria|mass
Finding|Intellectual Product|Hospital Course|14554,14560|false|false|false|C1511314|Breast Imaging Reporting and Data System|BIRADS
Disorder|Disease or Syndrome|Hospital Course|14566,14580|false|false|false|C0020676|Hypothyroidism|hypothyroidism
Finding|Mental Process|Discharge Condition|14607,14613|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|14607,14620|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|14607,14620|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|14614,14620|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14614,14620|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|14622,14627|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|14632,14640|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|14642,14664|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|14642,14664|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|14651,14664|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|14651,14664|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|14666,14671|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|14666,14671|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|14666,14671|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|14666,14671|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14676,14687|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|14689,14697|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|14689,14697|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|14689,14697|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|14698,14704|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14698,14704|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|14706,14716|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|14706,14716|false|false|false|C1561560|ambulatory encounter|Ambulatory
Finding|Social Behavior|Discharge Condition|14728,14738|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|14742,14745|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|14742,14745|false|false|false|C1454018|AICDA protein, human|aid
Finding|Gene or Genome|Discharge Condition|14742,14745|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|14742,14745|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Finding|Gene or Genome|Discharge Instructions|14792,14796|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Idea or Concept|Discharge Instructions|14827,14835|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Finding|Discharge Instructions|14848,14861|false|false|false|C0849970|Feeling tired|feeling tired
Finding|Finding|Discharge Instructions|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Intellectual Product|Discharge Instructions|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Finding|Sign or Symptom|Discharge Instructions|14856,14861|false|false|false|C0015672;C0849970;C3539029|Fatigue;Feel Tired question;Feeling tired|tired
Drug|Substance|Discharge Instructions|14871,14876|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Discharge Instructions|14871,14876|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Conceptual Entity|Discharge Instructions|14877,14883|false|false|false|C1709366|system output|output
Procedure|Health Care Activity|Discharge Instructions|14877,14883|false|false|false|C3251815|Measurement of fluid output|output
Finding|Finding|Discharge Instructions|14888,14894|false|false|false|C4554530|Bloody|bloody
Finding|Idea or Concept|Discharge Instructions|14919,14927|false|false|false|C1547192|Organization unit type - Hospital|hospital
Procedure|Diagnostic Procedure|Discharge Instructions|14933,14940|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|Discharge Instructions|14936,14940|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Finding|Finding|Discharge Instructions|14948,14958|false|false|false|C0450093|Very large|very large
Finding|Gene or Genome|Discharge Instructions|14953,14958|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|Discharge Instructions|14959,14964|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|14959,14964|false|false|false|C1546638|Fluid Specimen Code|fluid
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|14985,14991|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Anatomy|Body Space or Junction|Discharge Instructions|14985,14991|false|false|false|C0030797;C0559769;C4266535|Pelvic cavity structure;Pelvis;Pelvis+|pelvis
Disorder|Neoplastic Process|Discharge Instructions|14985,14991|false|false|false|C0153663|Malignant neoplasm of pelvis|pelvis
Finding|Finding|Discharge Instructions|14985,14991|false|false|false|C0812455|Pelvis problem|pelvis
Drug|Substance|Discharge Instructions|15027,15032|false|false|false|C1550628|Drain - SpecimenType|drain
Finding|Intellectual Product|Discharge Instructions|15027,15032|false|false|false|C1546604|Drain Specimen Code|drain
Finding|Intellectual Product|Discharge Instructions|15048,15052|false|false|false|C1720092|Once - dosing instruction fragment|once
Finding|Gene or Genome|Discharge Instructions|15075,15080|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Substance|Discharge Instructions|15081,15086|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|Discharge Instructions|15081,15086|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Conceptual Entity|Discharge Instructions|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Functional Concept|Discharge Instructions|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Idea or Concept|Discharge Instructions|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Finding|Intellectual Product|Discharge Instructions|15087,15097|false|false|false|C0600644;C1516698;C1704814;C1704815|Collection (action);Collection Object - UML Entity;Collections (publication);Item Collection|collection
Disorder|Disease or Syndrome|Discharge Instructions|15126,15131|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|15126,15131|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15126,15143|false|false|false|C0005841|Blood Transfusion|blood transfusion
Finding|Functional Concept|Discharge Instructions|15132,15143|false|false|false|C0199960||transfusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15132,15143|false|false|false|C0005841;C1879316|Blood Transfusion;Transfusion (procedure)|transfusion
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15158,15162|false|false|false|C2049629|Peripherally Inserted Central Catheter Line Insertion|PICC
Drug|Antibiotic|Discharge Instructions|15200,15211|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Finding|Idea or Concept|Discharge Instructions|15246,15254|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Discharge Instructions|15296,15304|false|false|false|C1547192|Organization unit type - Hospital|hospital
Anatomy|Body Location or Region|Discharge Instructions|15362,15366|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15362,15366|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|15362,15366|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|15362,15366|false|false|false|C0740941|Lung Problem|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15371,15377|false|false|false|C0006141|Breast|breast
Disorder|Neoplastic Process|Discharge Instructions|15371,15377|false|false|false|C0496956|Neoplasm of uncertain or unknown behavior of breast|breast
Finding|Finding|Discharge Instructions|15371,15377|false|false|false|C0567499|Breast problem|breast
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15371,15377|false|false|false|C0191838|Procedures on breast|breast
Finding|Finding|Discharge Instructions|15371,15385|false|false|false|C0567489|Lesion of breast|breast lesions
Finding|Finding|Discharge Instructions|15378,15385|false|false|false|C0221198|Lesion|lesions
Finding|Idea or Concept|Discharge Instructions|15403,15418|false|false|false|C0034866|Recommendation|recommendations
Finding|Idea or Concept|Discharge Instructions|15423,15431|false|false|false|C0549178|Continuous|Continue
Drug|Organic Chemical|Discharge Instructions|15439,15446|false|false|false|C0728963|Lovenox|Lovenox
Drug|Pharmacologic Substance|Discharge Instructions|15439,15446|false|false|false|C0728963|Lovenox|Lovenox
Finding|Idea or Concept|Discharge Instructions|15453,15456|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|15453,15456|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Disorder|Disease or Syndrome|Discharge Instructions|15470,15475|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|15470,15475|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|Discharge Instructions|15470,15480|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clot
Drug|Organic Chemical|Discharge Instructions|15476,15480|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|15476,15480|false|false|false|C0009074|clotrimazole|clot
Finding|Pathologic Function|Discharge Instructions|15476,15480|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Location or Region|Discharge Instructions|15490,15494|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15490,15494|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Discharge Instructions|15490,15494|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Discharge Instructions|15490,15494|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Discharge Instructions|15506,15516|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Discharge Instructions|15506,15524|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|Discharge Instructions|15517,15524|false|false|false|C0012634|Disease|disease
Finding|Intellectual Product|Discharge Instructions|15525,15531|false|false|false|C2348314|Doctor - Title|doctor
Finding|Idea or Concept|Discharge Instructions|15588,15594|false|false|false|C1554106|MDF AttributeType - Number|number
Event|Activity|Discharge Instructions|15608,15619|false|false|false|C0003629|Appointments|appointment
Finding|Intellectual Product|Discharge Instructions|15642,15646|false|false|false|C4724437|SURE Test|sure
Finding|Functional Concept|Discharge Instructions|15658,15664|false|false|false|C0205341;C1705914|Repeat;Repeat Object|repeat
Procedure|Diagnostic Procedure|Discharge Instructions|15665,15672|false|false|false|C0040405|X-Ray Computed Tomography|CT scan
Procedure|Diagnostic Procedure|Discharge Instructions|15668,15672|false|false|false|C0034606;C0441633|Radionuclide Imaging;Scanning|scan
Event|Activity|Discharge Instructions|15691,15702|false|false|false|C0003629|Appointments|appointment
Disorder|Disease or Syndrome|Discharge Instructions|15712,15722|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Discharge Instructions|15712,15730|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|Discharge Instructions|15723,15730|false|false|false|C0012634|Disease|disease
Finding|Intellectual Product|Discharge Instructions|15731,15737|false|false|false|C2348314|Doctor - Title|doctor
Drug|Antibiotic|Discharge Instructions|15763,15774|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Disorder|Disease or Syndrome|Discharge Instructions|15799,15809|false|false|false|C0009450|Communicable Diseases|infectious
Disorder|Disease or Syndrome|Discharge Instructions|15799,15817|false|false|false|C0009450|Communicable Diseases|infectious disease
Disorder|Disease or Syndrome|Discharge Instructions|15810,15817|false|false|false|C0012634|Disease|disease
Finding|Intellectual Product|Discharge Instructions|15818,15824|false|false|false|C2348314|Doctor - Title|doctor
Finding|Intellectual Product|Discharge Instructions|15887,15895|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|15887,15895|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|15903,15907|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|15903,15907|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|15903,15907|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|15903,15910|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|Discharge Instructions|15934,15942|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|15943,15955|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|15943,15955|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

