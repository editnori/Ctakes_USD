 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|43,52|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|43,52|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|43,57|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|77,86|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|77,86|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|77,86|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|77,91|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|109,114|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|133,136|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|133,136|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|144,151|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|144,151|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|SIMPLE_SEGMENT|153,160|false|false|false|||SURGERY
Finding|Finding|SIMPLE_SEGMENT|153,160|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|SIMPLE_SEGMENT|153,160|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|SIMPLE_SEGMENT|153,160|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|153,160|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Drug|Organic Chemical|Allergies|175,182|false|false|false|C0591292|Corgard|Corgard
Drug|Pharmacologic Substance|Allergies|175,182|false|false|false|C0591292|Corgard|Corgard
Drug|Amino Acid, Peptide, or Protein|Allergies|185,192|false|false|false|C0728763|Vasotec|Vasotec
Drug|Pharmacologic Substance|Allergies|185,192|false|false|false|C0728763|Vasotec|Vasotec
Event|Event|Allergies|195,204|false|false|false|||Attending
Finding|Functional Concept|Allergies|195,204|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|230,242|false|false|false|||incarcerated
Finding|Finding|Chief Complaint|230,242|false|false|false|C0392751|In prison (finding)|incarcerated
Disorder|Acquired Abnormality|Chief Complaint|230,258|false|false|false|C0401074|Irreducible inguinal hernia|incarcerated inguinal hernia
Anatomy|Body Location or Region|Chief Complaint|243,251|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|Chief Complaint|243,258|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Disorder|Anatomical Abnormality|Chief Complaint|252,258|false|false|false|C0019270|Hernia|hernia
Event|Event|Chief Complaint|252,258|false|false|false|||hernia
Finding|Classification|Chief Complaint|261,266|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|267,275|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|279,297|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|288,297|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|288,297|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|288,297|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|288,297|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|288,297|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Functional Concept|Chief Complaint|299,303|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Disorder|Acquired Abnormality|Chief Complaint|299,319|false|false|false|C0262537|Left inguinal hernia|Left inguinal hernia
Anatomy|Body Location or Region|Chief Complaint|304,312|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|Chief Complaint|304,319|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|304,326|false|false|false|C0021446|Repair of inguinal hernia|inguinal hernia repair
Disorder|Anatomical Abnormality|Chief Complaint|313,319|false|false|false|C0019270|Hernia|hernia
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|313,326|false|false|false|C0019328|Herniorrhaphy|hernia repair
Event|Event|Chief Complaint|320,326|false|false|false|||repair
Finding|Functional Concept|Chief Complaint|320,326|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Chief Complaint|320,326|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Chief Complaint|320,326|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|320,326|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Disorder|Disease or Syndrome|History of Present Illness|366,370|false|false|false|C0004238|Atrial Fibrillation|afib
Event|Event|History of Present Illness|366,370|false|false|false|||afib
Lab|Laboratory or Test Result|History of Present Illness|366,370|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|afib
Event|Event|History of Present Illness|374,382|false|false|false|||apixiban
Disorder|Disease or Syndrome|History of Present Illness|384,387|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|384,387|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|384,387|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|384,387|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|384,387|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|384,387|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|384,387|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|384,387|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Event|Event|History of Present Illness|392,396|false|false|false|||CABG
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|392,396|false|false|false|C0010055|Coronary Artery Bypass Surgery|CABG
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|402,409|false|false|false|C0007272|Carotid Arteries|carotid
Disorder|Disease or Syndrome|History of Present Illness|402,417|false|false|false|C0741975|carotid disease|carotid disease
Disorder|Disease or Syndrome|History of Present Illness|410,417|false|false|false|C0012634|Disease|disease
Event|Event|History of Present Illness|410,417|false|false|false|||disease
Disorder|Disease or Syndrome|History of Present Illness|420,424|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|420,424|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|420,424|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|420,424|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|425,434|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|History of Present Illness|425,434|false|false|false|||emphysema
Finding|Pathologic Function|History of Present Illness|425,434|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Disorder|Disease or Syndrome|History of Present Illness|447,456|false|false|false|C0032285|Pneumonia|pneumonia
Event|Event|History of Present Illness|447,456|false|false|false|||pneumonia
Event|Event|History of Present Illness|457,465|false|false|false|||presents
Finding|Functional Concept|History of Present Illness|470,478|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Finding|Intellectual Product|History of Present Illness|470,478|false|false|false|C1546398;C1546846;C1561552|Act Priority - elective;Admission Type - Elective;Visit Priority Code - Elective|elective
Event|Event|History of Present Illness|479,483|false|false|false|||left
Finding|Functional Concept|History of Present Illness|479,483|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|History of Present Illness|485,493|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|History of Present Illness|485,500|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|485,507|false|false|false|C0021446|Repair of inguinal hernia|inguinal hernia repair
Disorder|Anatomical Abnormality|History of Present Illness|494,500|false|false|false|C0019270|Hernia|hernia
Event|Event|History of Present Illness|494,500|false|false|false|||hernia
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|494,507|false|false|false|C0019328|Herniorrhaphy|hernia repair
Event|Event|History of Present Illness|501,507|false|false|false|||repair
Finding|Functional Concept|History of Present Illness|501,507|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|History of Present Illness|501,507|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|History of Present Illness|501,507|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|501,507|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Event|Event|History of Present Illness|509,514|false|false|false|||large
Finding|Gene or Genome|History of Present Illness|509,514|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Finding|History of Present Illness|521,533|false|false|false|C0392751|In prison (finding)|incarcerated
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|534,541|false|false|false|C0227391|Sigmoid colon|sigmoid
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|534,547|false|false|false|C0227391|Sigmoid colon|sigmoid colon
Disorder|Neoplastic Process|History of Present Illness|534,547|false|false|false|C0153436;C0496864|Benign neoplasm of sigmoid colon;Malignant neoplasm of sigmoid colon|sigmoid colon
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|542,547|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|History of Present Illness|542,547|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|History of Present Illness|542,547|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|History of Present Illness|542,547|false|false|false|C0750873|COLON PROBLEM|colon
Finding|Finding|Past Medical History|606,614|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Finding|Intellectual Product|Past Medical History|606,614|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|MODERATE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|615,622|false|false|false|C0007272|Carotid Arteries|CAROTID
Disorder|Disease or Syndrome|Past Medical History|615,630|false|false|false|C0741975|carotid disease|CAROTID DISEASE
Disorder|Disease or Syndrome|Past Medical History|623,630|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|623,630|false|false|false|||DISEASE
Disorder|Disease or Syndrome|Past Medical History|632,656|false|false|false|C0018802|Congestive heart failure|CONGESTIVE HEART FAILURE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|643,648|false|false|false|C0018787;C4037974|Chest>Heart;Heart|HEART
Disorder|Neoplastic Process|Past Medical History|643,648|false|false|false|C0153500;C0153957|Malignant neoplasm of heart;benign neoplasm of heart|HEART
Finding|Sign or Symptom|Past Medical History|643,648|false|false|false|C0795691|HEART PROBLEM|HEART
Disorder|Disease or Syndrome|Past Medical History|643,656|false|false|false|C0018801;C0018802|Congestive heart failure;Heart failure|HEART FAILURE
Event|Event|Past Medical History|649,656|false|false|false|||FAILURE
Finding|Functional Concept|Past Medical History|649,656|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Idea or Concept|Past Medical History|649,656|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Finding|Individual Behavior|Past Medical History|649,656|false|false|false|C0231174;C0680095;C5200924|Failure;Failure (biologic function);Personal failure|FAILURE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|658,666|false|false|false|C0018787|Heart|CORONARY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|658,673|false|false|false|C0205042|Coronary artery|CORONARY ARTERY
Disorder|Disease or Syndrome|Past Medical History|658,681|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|CORONARY ARTERY DISEASE
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|667,673|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Anatomy|Body System|Past Medical History|667,673|false|false|false|C0003842;C0226004|Arterial system;Arteries|ARTERY
Disorder|Disease or Syndrome|Past Medical History|667,681|false|false|false|C0852949|Arteriopathic disease|ARTERY DISEASE
Disorder|Disease or Syndrome|Past Medical History|674,681|false|false|false|C0012634|Disease|DISEASE
Event|Event|Past Medical History|674,681|false|false|false|||DISEASE
Anatomy|Body Location or Region|Past Medical History|683,699|false|false|false|C0744316|gastroesophageal|GASTROESOPHAGEAL
Disorder|Disease or Syndrome|Past Medical History|683,706|false|false|false|C0017168|Gastroesophageal reflux disease|GASTROESOPHAGEAL REFLUX
Finding|Finding|Past Medical History|683,706|false|false|false|C3813607;C4317146|Acid reflux;Infantile Gastroesophageal Reflux|GASTROESOPHAGEAL REFLUX
Event|Event|Past Medical History|700,706|false|false|false|||REFLUX
Finding|Pathologic Function|Past Medical History|700,706|false|false|false|C0232483|Reflux|REFLUX
Disorder|Disease or Syndrome|Past Medical History|708,720|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|708,720|false|false|false|||HYPERTENSION
Finding|Finding|Past Medical History|722,728|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Finding|Intellectual Product|Past Medical History|722,728|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|SEVERE
Disorder|Disease or Syndrome|Past Medical History|729,738|false|false|false|C0034067|Pulmonary Emphysema|EMPHYSEMA
Event|Event|Past Medical History|729,738|false|false|false|||EMPHYSEMA
Finding|Pathologic Function|Past Medical History|729,738|false|false|false|C0013990|Pathological accumulation of air in tissues|EMPHYSEMA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|740,749|false|false|false|C0024109|Lung|PULMONARY
Attribute|Clinical Attribute|Past Medical History|740,749|false|false|false|C2707265||PULMONARY
Finding|Finding|Past Medical History|740,749|false|false|false|C4522268|Pulmonary (intended site)|PULMONARY
Finding|Pathologic Function|Past Medical History|740,762|false|false|false|C0020542|Pulmonary Hypertension|PULMONARY HYPERTENSION
Disorder|Disease or Syndrome|Past Medical History|750,762|false|false|false|C0020538|Hypertensive disease|HYPERTENSION
Event|Event|Past Medical History|750,762|false|false|false|||HYPERTENSION
Finding|Functional Concept|Past Medical History|764,769|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|764,783|false|false|false|C0225916|Structure of right branch of atrioventricular bundle|RIGHT BUNDLE BRANCH
Disorder|Disease or Syndrome|Past Medical History|764,789|false|false|false|C0085615|Right bundle branch block|RIGHT BUNDLE BRANCH BLOCK
Finding|Finding|Past Medical History|764,789|false|false|false|C0344421||RIGHT BUNDLE BRANCH BLOCK
Disorder|Disease or Syndrome|Past Medical History|770,789|false|false|false|C0006384;C1879286|Bundle-Branch Block;Hereditary bundle branch system defect|BUNDLE BRANCH BLOCK
Drug|Chemical Viewed Structurally|Past Medical History|777,783|false|false|false|C1881507|Macromolecular Branch|BRANCH
Drug|Biomedical or Dental Material|Past Medical History|784,789|false|false|false|C1706085|Block Dosage Form|BLOCK
Event|Event|Past Medical History|784,789|false|false|false|||BLOCK
Finding|Body Substance|Past Medical History|784,789|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Finding|Past Medical History|784,789|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Functional Concept|Past Medical History|784,789|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|BLOCK
Finding|Pathologic Function|Past Medical History|791,819|false|false|false|C1704272|Benign Prostatic Hyperplasia|BENIGN PROSTATIC HYPERTROPHY
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|798,807|false|false|false|C0033572|Prostate|PROSTATIC
Disorder|Disease or Syndrome|Past Medical History|798,819|false|false|false|C1739363|Prostatic Hypertrophy|PROSTATIC HYPERTROPHY
Finding|Pathologic Function|Past Medical History|798,819|false|false|false|C1704272;C2937421|Benign Prostatic Hyperplasia;Prostatic Hyperplasia|PROSTATIC HYPERTROPHY
Event|Event|Past Medical History|808,819|false|false|false|||HYPERTROPHY
Finding|Pathologic Function|Past Medical History|808,819|false|false|false|C0020564|Hypertrophy|HYPERTROPHY
Disorder|Disease or Syndrome|Past Medical History|821,835|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|HYPERLIPIDEMIA
Event|Event|Past Medical History|821,835|false|false|false|||HYPERLIPIDEMIA
Finding|Finding|Past Medical History|821,835|false|false|false|C0428465|Serum lipids high (finding)|HYPERLIPIDEMIA
Event|Event|Past Medical History|837,847|false|false|false|||PAROXYSMAL
Disorder|Disease or Syndrome|Past Medical History|837,867|false|false|false|C0235480|Paroxysmal atrial fibrillation|PAROXYSMAL ATRIAL FIBRILLATION
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|848,854|false|false|false|C0018792|Heart Atrium|ATRIAL
Attribute|Clinical Attribute|Past Medical History|848,867|false|false|false|C2926591||ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|848,867|false|false|false|C0004238|Atrial Fibrillation|ATRIAL FIBRILLATION
Lab|Laboratory or Test Result|Past Medical History|848,867|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|ATRIAL FIBRILLATION
Disorder|Disease or Syndrome|Past Medical History|855,867|false|false|false|C0232197|Fibrillation|FIBRILLATION
Event|Event|Past Medical History|855,867|false|false|false|||FIBRILLATION
Event|Event|Past Surgical History|914,927|false|false|false|||CARDIOVERSION
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|914,927|false|false|false|C0013778|Electric Countershock|CARDIOVERSION
Finding|Functional Concept|Past Surgical History|933,938|false|false|false|C1552823|Table Cell Horizontal Align - right|RIGHT
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|933,949|false|false|false|C1261075|Structure of right lower lobe of lung|RIGHT LOWER LOBE
Anatomy|Body Location or Region|Past Surgical History|939,944|false|false|false|C1548802|Body Site Modifier - Lower|LOWER
Event|Activity|Past Surgical History|939,944|false|false|false|C2003888|Lower (action)|LOWER
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|939,949|false|false|false|C0225758|Structure of lower lobe of lung|LOWER LOBE
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|945,949|false|false|false|C0796494|lobe|LOBE
Finding|Gene or Genome|Past Surgical History|945,949|false|false|false|C1428707;C3539671|AKT1S1 gene;AKT1S1 wt Allele|LOBE
Event|Event|Past Surgical History|950,959|false|false|false|||LOBECTOMY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|950,959|false|true|false|C0023928|Lobectomy|LOBECTOMY
Anatomy|Body Part, Organ, or Organ Component|Past Surgical History|965,973|false|false|false|C0018787|Heart|CORONARY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|965,980|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|965,988|false|false|false|C0010055|Coronary Artery Bypass Surgery|CORONARY BYPASS SURGERY
Event|Event|Past Surgical History|974,980|false|false|false|||BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|974,980|false|false|false|C0813207|Creation of shunt|BYPASS
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|974,988|false|false|false|C1536078|Bypass surgery|BYPASS SURGERY
Event|Event|Past Surgical History|981,988|false|false|false|||SURGERY
Finding|Finding|Past Surgical History|981,988|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Functional Concept|Past Surgical History|981,988|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Finding|Idea or Concept|Past Surgical History|981,988|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|SURGERY
Procedure|Therapeutic or Preventive Procedure|Past Surgical History|981,988|false|false|false|C0543467|Operative Surgical Procedures|SURGERY
Finding|Classification|General Exam|1067,1070|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Finding|Gene or Genome|General Exam|1067,1070|false|false|false|C2239486;C4084748;C4521767|GEN1 gene;GEN1 wt Allele;United States Military Commissioned Officer O10 (qualifier value)|Gen
Event|Event|General Exam|1072,1077|false|false|false|||Awake
Attribute|Clinical Attribute|General Exam|1082,1087|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|1082,1087|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|1082,1087|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|1082,1087|false|false|false|||alert
Finding|Finding|General Exam|1082,1087|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|1082,1087|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|1082,1087|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|1114,1120|false|false|false|||rhythm
Finding|Finding|General Exam|1114,1120|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|1114,1120|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Activity|General Exam|1129,1133|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|1129,1133|false|false|false|||rate
Finding|Idea or Concept|General Exam|1129,1133|false|false|false|C1549480|Amount type - Rate|rate
Attribute|Clinical Attribute|General Exam|1134,1138|false|false|false|C0231832|Respiratory rate|Resp
Disorder|Disease or Syndrome|General Exam|1134,1138|false|false|false|C0851355|Respiratory, thoracic and mediastinal disorders|Resp
Event|Event|General Exam|1134,1138|false|false|false|||Resp
Drug|Organic Chemical|General Exam|1140,1144|false|false|false|C0951233|cetrimonium bromide|CTAB
Event|Event|General Exam|1140,1144|false|false|false|||CTAB
Disorder|Disease or Syndrome|General Exam|1149,1153|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|1149,1153|false|false|false|||Soft
Anatomy|Body Location or Region|General Exam|1181,1189|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|General Exam|1181,1189|false|false|false|C0332803|Surgical wound|incision
Event|Event|General Exam|1181,1189|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|General Exam|1181,1189|false|false|false|C0184898|Surgical incisions|incision
Anatomy|Body Location or Region|General Exam|1205,1213|false|false|false|C2338258|Cranial incision point|Incision
Disorder|Injury or Poisoning|General Exam|1205,1213|false|false|false|C0332803|Surgical wound|Incision
Procedure|Therapeutic or Preventive Procedure|General Exam|1205,1213|false|false|false|C0184898|Surgical incisions|Incision
Event|Activity|General Exam|1214,1219|false|false|false|C1947930|Cleaning (activity)|clean
Event|Event|General Exam|1230,1236|false|false|false|||intact
Finding|Finding|General Exam|1230,1236|false|false|false|C1554187|Gender Status - Intact|intact
Disorder|Disease or Syndrome|General Exam|1245,1253|false|false|false|C0041834|Erythema|erythema
Event|Event|General Exam|1245,1253|false|false|false|||erythema
Disorder|Congenital Abnormality|General Exam|1254,1257|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|1254,1257|false|false|false|||Ext
Finding|Gene or Genome|General Exam|1254,1257|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|1259,1263|false|false|false|||Warm
Finding|Finding|General Exam|1259,1263|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|1259,1263|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|1268,1272|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|1273,1281|false|false|false|||perfused
Event|Event|Hospital Course|1342,1350|false|false|false|||admitted
Event|Event|Hospital Course|1387,1393|false|false|false|||repair
Finding|Functional Concept|Hospital Course|1387,1393|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Hospital Course|1387,1393|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Hospital Course|1387,1393|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1387,1393|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Finding|Functional Concept|Hospital Course|1399,1403|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Finding|Hospital Course|1405,1417|false|false|false|C0392751|In prison (finding)|incarcerated
Disorder|Acquired Abnormality|Hospital Course|1405,1433|false|false|false|C0401074|Irreducible inguinal hernia|incarcerated inguinal hernia
Anatomy|Body Location or Region|Hospital Course|1418,1426|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|Hospital Course|1418,1433|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Disorder|Anatomical Abnormality|Hospital Course|1427,1433|false|false|false|C0019270|Hernia|hernia
Event|Event|Hospital Course|1427,1433|false|false|false|||hernia
Event|Event|Hospital Course|1439,1446|false|false|false|||details
Attribute|Clinical Attribute|Hospital Course|1454,1463|false|false|false|C0945766||procedure
Event|Event|Hospital Course|1454,1463|false|false|false|||procedure
Event|Occupational Activity|Hospital Course|1454,1463|false|false|false|C1546467|Act Class - procedure|procedure
Finding|Functional Concept|Hospital Course|1454,1463|false|false|false|C2700391|Procedure (set of actions)|procedure
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1454,1463|false|false|false|C0184661|Interventional procedure|procedure
Event|Event|Hospital Course|1473,1478|false|false|false|||refer
Finding|Intellectual Product|Hospital Course|1486,1502|false|false|false|C1269801|Operative report|operative report
Attribute|Clinical Attribute|Hospital Course|1496,1502|false|false|false|C4255046||report
Event|Event|Hospital Course|1496,1502|false|false|false|||report
Finding|Intellectual Product|Hospital Course|1496,1502|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Hospital Course|1496,1502|false|false|false|C0700287|Reporting|report
Event|Event|Hospital Course|1522,1528|false|false|false|||course
Event|Event|Hospital Course|1534,1547|false|false|false|||uncomplicated
Finding|Intellectual Product|Hospital Course|1557,1562|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|brief
Event|Event|Hospital Course|1563,1567|false|false|false|||stay
Event|Event|Hospital Course|1589,1600|false|false|false|||transferred
Event|Event|Hospital Course|1616,1623|false|false|false|||nursing
Finding|Organism Function|Hospital Course|1616,1623|false|false|false|C0006147|Breast Feeding|nursing
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1616,1623|false|false|false|C0028678|RNAx nursing therapy actions|nursing
Anatomy|Anatomical Structure|Hospital Course|1624,1629|false|false|false|C3714591|Floor (anatomic)|floor
Attribute|Clinical Attribute|Hospital Course|1635,1639|false|false|false|C2598155||pain
Event|Event|Hospital Course|1635,1639|false|false|false|||pain
Finding|Functional Concept|Hospital Course|1635,1639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1635,1639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|1645,1655|false|false|false|||controlled
Drug|Pharmacologic Substance|Hospital Course|1661,1674|false|false|false|C1971835|IV medication|IV medication
Drug|Pharmacologic Substance|Hospital Course|1664,1674|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|1664,1674|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|1664,1674|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|1694,1701|false|false|false|||started
Finding|Daily or Recreational Activity|Hospital Course|1708,1720|false|false|false|C0184625||regular diet
Drug|Food|Hospital Course|1716,1720|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1716,1720|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1716,1720|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1716,1720|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|Hospital Course|1730,1734|false|false|false|C2598155||pain
Event|Event|Hospital Course|1730,1734|false|false|false|||pain
Finding|Functional Concept|Hospital Course|1730,1734|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1730,1734|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|1739,1749|false|false|false|||controlled
Attribute|Clinical Attribute|Hospital Course|1758,1762|false|false|false|C2598155||pain
Event|Event|Hospital Course|1758,1762|false|false|false|||pain
Finding|Functional Concept|Hospital Course|1758,1762|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1758,1762|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Hospital Course|1764,1774|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|1764,1774|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|1764,1774|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|1779,1785|false|false|false|||voided
Event|Activity|Hospital Course|1794,1799|true|false|false|C5966184|Issue (action)|issue
Event|Event|Hospital Course|1794,1799|false|false|false|||issue
Finding|Finding|Hospital Course|1794,1799|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|Hospital Course|1794,1799|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|Hospital Course|1808,1818|false|false|false|||ambulating
Drug|Organic Chemical|Hospital Course|1841,1846|false|false|false|C2356088|Halls|halls
Drug|Pharmacologic Substance|Hospital Course|1841,1846|false|false|false|C2356088|Halls|halls
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|1863,1868|false|false|false|C0021853|Intestines|bowel
Procedure|Health Care Activity|Hospital Course|1863,1876|false|false|false|C5979615|Bowel Regimen|bowel regimen
Event|Event|Hospital Course|1869,1876|false|false|false|||regimen
Finding|Intellectual Product|Hospital Course|1869,1876|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1869,1876|false|false|false|C0040808|Treatment Protocols|regimen
Event|Event|Hospital Course|1883,1889|false|false|false|||passed
Event|Event|Hospital Course|1890,1896|false|false|false|||flatus
Finding|Sign or Symptom|Hospital Course|1890,1896|false|false|false|C0016204|Flatulence|flatus
Event|Event|Hospital Course|1912,1921|false|false|false|||continued
Event|Event|Hospital Course|1925,1933|false|false|false|||tolerate
Drug|Food|Hospital Course|1938,1942|false|false|false|C0012155;C3668949|Diet;Diet (animal life circumstance)|diet
Event|Event|Hospital Course|1938,1942|false|false|false|||diet
Finding|Functional Concept|Hospital Course|1938,1942|false|false|false|C1549512|diet - supply|diet
Procedure|Health Care Activity|Hospital Course|1938,1942|false|false|false|C0012159|Diet therapy|diet
Attribute|Clinical Attribute|Hospital Course|1949,1953|false|false|false|C2598155||pain
Event|Event|Hospital Course|1949,1953|false|false|false|||pain
Finding|Functional Concept|Hospital Course|1949,1953|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|1949,1953|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|1958,1962|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|1963,1973|false|false|false|||controlled
Anatomy|Body Space or Junction|Hospital Course|1977,1981|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|1977,1981|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|1977,1981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|1977,1981|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Drug|Pharmacologic Substance|Hospital Course|1977,1992|false|false|false|C5848556|Oral medication (substance)|oral medication
Procedure|Therapeutic or Preventive Procedure|Hospital Course|1977,1992|false|false|false|C0175795|Oral Medication|oral medication
Drug|Pharmacologic Substance|Hospital Course|1982,1992|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|1982,1992|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|1982,1992|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|2001,2010|false|false|false|||continued
Event|Event|Hospital Course|2015,2023|false|false|false|||ambulate
Finding|Finding|Hospital Course|2015,2023|false|false|false|C4036205|Ambulate|ambulate
Event|Event|Hospital Course|2046,2056|false|false|false|||discharged
Event|Event|Hospital Course|2057,2061|false|false|false|||home
Finding|Idea or Concept|Hospital Course|2057,2061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|2057,2061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|2057,2061|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|2065,2071|false|false|false|||stable
Finding|Intellectual Product|Hospital Course|2065,2071|false|false|false|C1547311|Patient Condition Code - Stable|stable
Attribute|Clinical Attribute|Hospital Course|2073,2082|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Hospital Course|2073,2082|false|false|false|C0012634|Disease|condition
Event|Event|Hospital Course|2073,2082|false|false|false|||condition
Finding|Conceptual Entity|Hospital Course|2073,2082|false|false|false|C1705253|Logical Condition|condition
Event|Event|Hospital Course|2086,2089|false|false|false|||POD
Event|Event|Hospital Course|2107,2113|false|false|false|||follow
Event|Event|Hospital Course|2134,2143|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|2134,2143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|2134,2143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|2134,2143|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|2134,2143|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|2134,2155|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|2144,2155|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|2144,2155|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|2144,2155|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|2144,2155|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|2160,2170|false|false|false|C0002598|amiodarone|Amiodarone
Drug|Pharmacologic Substance|Hospital Course|2160,2170|false|false|false|C0002598|amiodarone|Amiodarone
Event|Event|Hospital Course|2160,2170|false|false|false|||Amiodarone
Procedure|Laboratory Procedure|Hospital Course|2160,2170|false|false|false|C5399868|Drug assay amiodarone|Amiodarone
Drug|Organic Chemical|Hospital Course|2191,2199|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|2191,2199|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|2208,2211|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2208,2211|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|2208,2211|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|2208,2211|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|2208,2211|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|2216,2223|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|2216,2223|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|2243,2251|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|2243,2251|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|2243,2251|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|2243,2258|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|2243,2258|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|2252,2258|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|2252,2258|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|2252,2258|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|2252,2258|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|2252,2258|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|2252,2258|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|2269,2272|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|2269,2272|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|2269,2272|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|2269,2272|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|2269,2272|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|2277,2285|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Hospital Course|2277,2285|false|false|false|C0126174|losartan|Losartan
Event|Event|Hospital Course|2277,2285|false|false|false|||Losartan
Drug|Organic Chemical|Hospital Course|2277,2295|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Hospital Course|2277,2295|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Hospital Course|2286,2295|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Hospital Course|2286,2295|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Hospital Course|2286,2295|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Hospital Course|2286,2295|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Hospital Course|2286,2295|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Hospital Course|2286,2295|false|false|false|||Potassium
Finding|Physiologic Function|Hospital Course|2286,2295|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Hospital Course|2286,2295|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Hospital Course|2315,2325|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Pharmacologic Substance|Hospital Course|2315,2325|false|false|false|C0028978|omeprazole|Omeprazole
Drug|Organic Chemical|Hospital Course|2345,2356|false|false|false|C0040869|triamterene|Triamterene
Drug|Pharmacologic Substance|Hospital Course|2345,2356|false|false|false|C0040869|triamterene|Triamterene
Drug|Organic Chemical|Hospital Course|2357,2361|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Drug|Pharmacologic Substance|Hospital Course|2357,2361|false|false|false|C0020261|hydrochlorothiazide|HCTZ
Event|Event|Hospital Course|2357,2361|false|false|false|||HCTZ
Disorder|Congenital Abnormality|Hospital Course|2374,2377|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|2374,2377|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|2374,2377|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|2374,2377|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2374,2377|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|2391,2404|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|2391,2404|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|2391,2404|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|2391,2404|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|2420,2423|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|2424,2428|false|false|false|C2598155||pain
Event|Event|Hospital Course|2424,2428|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2424,2428|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2424,2428|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|2432,2437|false|false|false|||fever
Finding|Finding|Hospital Course|2432,2437|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|2432,2437|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Hospital Course|2446,2452|false|false|false|||exceed
Finding|Idea or Concept|Hospital Course|2465,2468|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|2465,2468|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Drug|Organic Chemical|Hospital Course|2475,2488|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|Hospital Course|2475,2488|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|Hospital Course|2475,2488|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|Hospital Course|2475,2488|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Drug|Biomedical or Dental Material|Hospital Course|2500,2506|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|2500,2506|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|2510,2518|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|2513,2518|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|2513,2518|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|2544,2550|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|2551,2558|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|2551,2558|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|2565,2574|false|false|false|C0030049|oxycodone|OxycoDONE
Drug|Pharmacologic Substance|Hospital Course|2565,2574|false|false|false|C0030049|oxycodone|OxycoDONE
Event|Event|Hospital Course|2565,2574|false|false|false|||OxycoDONE
Procedure|Laboratory Procedure|Hospital Course|2565,2574|false|false|false|C0524222|Oxycodone measurement|OxycoDONE
Finding|Idea or Concept|Hospital Course|2576,2585|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Finding|Intellectual Product|Hospital Course|2576,2585|false|false|false|C1548167;C1697779|Query Priority - Immediate;immediate - ResponseCode|Immediate
Drug|Biomedical or Dental Material|Hospital Course|2576,2593|false|false|false|C1708470|Immediate Release Dosage Form|Immediate Release
Event|Event|Hospital Course|2586,2593|false|false|false|||Release
Finding|Functional Concept|Hospital Course|2586,2593|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|2586,2593|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2586,2593|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Finding|Gene or Genome|Hospital Course|2608,2611|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|2612,2616|false|false|false|C2598155||pain
Event|Event|Hospital Course|2612,2616|false|false|false|||pain
Finding|Functional Concept|Hospital Course|2612,2616|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|2612,2616|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Hospital Course|2618,2620|false|false|false|||RX
Drug|Organic Chemical|Hospital Course|2622,2631|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|2622,2631|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|2622,2631|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|2622,2631|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Biomedical or Dental Material|Hospital Course|2641,2647|false|false|false|C0039225|Tablet Dosage Form|tablet
Event|Event|Hospital Course|2641,2647|false|false|false|||tablet
Finding|Functional Concept|Hospital Course|2651,2659|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Hospital Course|2654,2659|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|2654,2659|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Activity|Hospital Course|2674,2678|false|false|false|C1880359|Dispense (activity)|Disp
Finding|Gene or Genome|Hospital Course|2674,2678|false|false|false|C2828567|PRSS30P gene|Disp
Drug|Biomedical or Dental Material|Hospital Course|2685,2691|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|2692,2699|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|2692,2699|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|2707,2712|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|2707,2712|false|false|false|C3489575|sennosides, USP|Senna
Drug|Organic Chemical|Hospital Course|2759,2768|false|false|false|C0030049|oxycodone|oxycodone
Drug|Pharmacologic Substance|Hospital Course|2759,2768|false|false|false|C0030049|oxycodone|oxycodone
Event|Event|Hospital Course|2759,2768|false|false|false|||oxycodone
Procedure|Laboratory Procedure|Hospital Course|2759,2768|false|false|false|C0524222|Oxycodone measurement|oxycodone
Drug|Organic Chemical|Hospital Course|2775,2785|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|Hospital Course|2775,2785|false|false|false|C3489575|sennosides, USP|sennosides
Event|Event|Hospital Course|2775,2785|false|false|false|||sennosides
Procedure|Therapeutic or Preventive Procedure|Hospital Course|2787,2791|false|false|false|C0058928|ECHO protocol|Evac
Drug|Organic Chemical|Hospital Course|2787,2797|false|false|false|C0720314;C1995730|Evac-U-Gen;Evac-U-Gen Reformulated Jan 2008|Evac-U-Gen
Drug|Pharmacologic Substance|Hospital Course|2787,2797|false|false|false|C0720314;C1995730|Evac-U-Gen;Evac-U-Gen Reformulated Jan 2008|Evac-U-Gen
Drug|Organic Chemical|Hospital Course|2799,2809|false|false|false|C3489575|sennosides, USP|sennosides
Drug|Pharmacologic Substance|Hospital Course|2799,2809|false|false|false|C3489575|sennosides, USP|sennosides
Event|Event|Hospital Course|2799,2809|false|false|false|||sennosides
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|2821,2828|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|2821,2828|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|2821,2828|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Location or Region|Hospital Course|2833,2838|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Hospital Course|2833,2838|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Drug|Biomedical or Dental Material|Hospital Course|2855,2861|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Hospital Course|2862,2869|false|false|false|||Refills
Finding|Idea or Concept|Hospital Course|2862,2869|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Hospital Course|2877,2882|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|2877,2882|false|false|false|C2369992|Align|Align
Drug|Pharmacologic Substance|Hospital Course|2884,2908|false|false|false|C4019097|herbal medicines bifidobacterium infantis|bifidobacterium infantis
Event|Event|Hospital Course|2900,2908|false|false|false|||infantis
Anatomy|Body Space or Junction|Hospital Course|2915,2919|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2915,2919|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2915,2919|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2915,2919|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|2920,2925|false|false|false|||DAILY
Drug|Biologically Active Substance|Hospital Course|2931,2939|false|false|false|C0009235|Coenzymes|coenzyme
Drug|Organic Chemical|Hospital Course|2931,2939|false|false|false|C0009235|Coenzymes|coenzyme
Event|Event|Hospital Course|2931,2939|false|false|false|||coenzyme
Drug|Biologically Active Substance|Hospital Course|2931,2943|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Organic Chemical|Hospital Course|2931,2943|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Drug|Pharmacologic Substance|Hospital Course|2931,2943|false|false|false|C0041536|ubidecarenone|coenzyme Q10
Event|Event|Hospital Course|2940,2943|false|false|false|||Q10
Finding|Gene or Genome|Hospital Course|2940,2943|false|false|false|C1414333;C2827473|AGO2 gene;AGO2 wt Allele|Q10
Anatomy|Body Space or Junction|Hospital Course|2951,2955|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|2951,2955|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|2951,2955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|2951,2955|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|2956,2961|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|2967,2979|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Drug|Pharmacologic Substance|Hospital Course|2967,2979|false|false|false|C0965129|rosuvastatin|Rosuvastatin
Event|Event|Hospital Course|2967,2979|false|false|false|||Rosuvastatin
Drug|Organic Chemical|Hospital Course|2967,2987|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Pharmacologic Substance|Hospital Course|2967,2987|false|false|false|C1101751|rosuvastatin calcium|Rosuvastatin Calcium
Drug|Biologically Active Substance|Hospital Course|2980,2987|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Hospital Course|2980,2987|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Hospital Course|2980,2987|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Hospital Course|2980,2987|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Hospital Course|2980,2987|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|Hospital Course|2980,2987|false|false|false|||Calcium
Finding|Physiologic Function|Hospital Course|2980,2987|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Hospital Course|2980,2987|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Biologically Active Substance|Hospital Course|2980,2990|false|false|false|C0006675|calcium|Calcium 40
Drug|Element, Ion, or Isotope|Hospital Course|2980,2990|false|false|false|C0006675|calcium|Calcium 40
Drug|Pharmacologic Substance|Hospital Course|2980,2990|false|false|false|C0006675|calcium|Calcium 40
Event|Event|Hospital Course|2997,3000|false|false|false|||QPM
Drug|Organic Chemical|Hospital Course|3006,3013|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|3006,3013|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|3006,3013|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|3006,3015|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|3006,3015|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|3006,3015|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|3006,3015|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|3006,3015|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|3014,3015|false|false|false|||D
Event|Event|Hospital Course|3021,3025|false|false|false|||UNIT
Event|Event|Hospital Course|3039,3048|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3039,3048|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3039,3048|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3039,3048|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3039,3048|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|3039,3060|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|3039,3060|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|3049,3060|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|3049,3060|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|3049,3060|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Hospital Course|3062,3066|false|false|false|||Home
Finding|Idea or Concept|Hospital Course|3062,3066|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|3062,3066|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|3062,3066|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Hospital Course|3072,3079|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Hospital Course|3072,3079|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Hospital Course|3082,3090|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|3082,3090|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Hospital Course|3098,3107|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|3098,3107|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|3098,3107|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|3098,3107|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|3098,3107|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|3098,3117|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|3108,3117|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|3108,3117|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|3108,3117|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|3108,3117|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|3108,3117|false|false|false|C0011900|Diagnosis|Diagnosis
Anatomy|Body Location or Region|Hospital Course|3119,3127|false|false|false|C0018246|Inguinal region|Inguinal
Disorder|Anatomical Abnormality|Hospital Course|3119,3134|false|false|false|C0019294|Hernia, Inguinal|Inguinal hernia
Disorder|Anatomical Abnormality|Hospital Course|3128,3134|false|false|false|C0019270|Hernia|hernia
Event|Event|Hospital Course|3128,3134|false|false|false|||hernia
Finding|Mental Process|Discharge Condition|3158,3164|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|3158,3171|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|3158,3171|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|3165,3171|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|3165,3171|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|3173,3178|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|3173,3178|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|3183,3191|false|false|false|||coherent
Finding|Finding|Discharge Condition|3183,3191|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|3193,3198|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|3193,3215|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|3193,3215|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|3202,3215|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|3202,3215|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|3202,3215|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|3217,3222|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|3217,3222|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|3217,3222|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|3217,3222|false|false|false|||Alert
Finding|Finding|Discharge Condition|3217,3222|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|3217,3222|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|3217,3222|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|3227,3238|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|3227,3238|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|3240,3248|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|3240,3248|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|3240,3248|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|3249,3255|false|false|false|C5889824||Status
Event|Event|Discharge Condition|3249,3255|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|3249,3255|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|3257,3267|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|3257,3267|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|3257,3267|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|3257,3267|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|3257,3267|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|3270,3281|false|false|false|||Independent
Finding|Finding|Discharge Condition|3270,3281|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|3270,3281|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|3309,3313|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|3332,3340|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|3332,3340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|3332,3340|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|3348,3352|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|3348,3352|false|false|false|||care
Finding|Finding|Discharge Instructions|3348,3352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|3348,3352|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|3348,3355|false|false|false|C1555558|care of - AddressPartType|care of
Event|Event|Discharge Instructions|3387,3395|false|false|false|||admitted
Finding|Idea or Concept|Discharge Instructions|3403,3411|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|3430,3436|false|false|false|||repair
Finding|Functional Concept|Discharge Instructions|3430,3436|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Finding|Organism Function|Discharge Instructions|3430,3436|false|false|false|C0043240;C4319951|Repair;Wound Healing|repair
Procedure|Health Care Activity|Discharge Instructions|3430,3436|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3430,3436|false|false|false|C0374711;C1705181|Repair - Remedial Action;Surgical repair|repair
Anatomy|Body Location or Region|Discharge Instructions|3445,3453|false|false|false|C0018246|Inguinal region|inguinal
Disorder|Anatomical Abnormality|Discharge Instructions|3445,3460|false|false|false|C0019294|Hernia, Inguinal|inguinal hernia
Disorder|Anatomical Abnormality|Discharge Instructions|3454,3460|false|false|false|C0019270|Hernia|hernia
Event|Event|Discharge Instructions|3454,3460|false|false|false|||hernia
Event|Event|Discharge Instructions|3472,3481|false|false|false|||recovered
Event|Event|Discharge Instructions|3487,3494|false|false|false|||surgery
Finding|Finding|Discharge Instructions|3487,3494|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|3487,3494|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|3487,3494|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|3487,3494|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|3507,3512|false|false|false|||ready
Event|Event|Discharge Instructions|3519,3529|false|false|false|||discharged
Event|Event|Discharge Instructions|3530,3534|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|3530,3534|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|3530,3534|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|3530,3534|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|3555,3570|false|false|false|||recommendations
Finding|Idea or Concept|Discharge Instructions|3555,3570|false|false|false|C0034866|Recommendation|recommendations
Event|Event|Discharge Instructions|3580,3586|false|false|false|||ensure
Finding|Finding|Discharge Instructions|3601,3611|false|false|false|C5453124|Uneventful|uneventful
Event|Activity|Discharge Instructions|3612,3620|false|false|false|C0237820||recovery
Event|Event|Discharge Instructions|3612,3620|false|false|false|||recovery
Finding|Organism Function|Discharge Instructions|3612,3620|false|false|false|C2004454|Recovery - healing process|recovery
Event|Activity|Discharge Instructions|3625,3633|false|false|false|C0441655|Activities|ACTIVITY
Event|Event|Discharge Instructions|3625,3633|false|false|false|||ACTIVITY
Finding|Daily or Recreational Activity|Discharge Instructions|3625,3633|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Finding|Finding|Discharge Instructions|3625,3633|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|ACTIVITY
Event|Event|Discharge Instructions|3644,3649|false|false|false|||drive
Event|Event|Discharge Instructions|3673,3679|false|false|false|||taking
Attribute|Clinical Attribute|Discharge Instructions|3680,3684|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|3680,3684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|3680,3684|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|3680,3693|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|3680,3693|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|3680,3693|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|3685,3693|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|3685,3693|false|false|false|||medicine
Event|Event|Discharge Instructions|3714,3721|false|false|false|||respond
Event|Event|Discharge Instructions|3728,3737|false|false|false|||emergency
Finding|Finding|Discharge Instructions|3728,3737|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|3728,3737|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|3728,3737|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|3728,3737|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|3728,3737|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|3728,3737|false|false|false|C1553500|emergency encounter|emergency
Event|Event|Discharge Instructions|3755,3761|false|false|false|||stairs
Finding|Finding|Discharge Instructions|3755,3761|false|false|false|C4300351|Prior functioning.stairs|stairs
Event|Event|Discharge Instructions|3790,3795|false|false|false|||avoid
Event|Event|Discharge Instructions|3796,3805|false|false|false|||traveling
Event|Event|Discharge Instructions|3811,3820|false|false|false|||distances
Event|Event|Discharge Instructions|3832,3835|false|false|false|||see
Attribute|Clinical Attribute|Discharge Instructions|3841,3848|false|false|false|C5444295||surgeon
Finding|Idea or Concept|Discharge Instructions|3857,3861|false|false|false|C1552851|next - HtmlLinkType|next
Event|Event|Discharge Instructions|3862,3867|false|false|false|||visit
Finding|Social Behavior|Discharge Instructions|3862,3867|false|false|false|C0545082|Visit|visit
Procedure|Laboratory Procedure|Discharge Instructions|3895,3898|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Attribute|Clinical Attribute|Discharge Instructions|3932,3938|false|false|false|C0944911||weight
Event|Event|Discharge Instructions|3932,3938|false|false|false|||weight
Finding|Finding|Discharge Instructions|3932,3938|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Discharge Instructions|3932,3938|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Discharge Instructions|3932,3938|false|false|false|C1305866|Weighing patient|weight
Event|Event|Discharge Instructions|3944,3953|false|false|false|||briefcase
Event|Event|Discharge Instructions|3959,3962|false|false|false|||bag
Finding|Intellectual Product|Discharge Instructions|3959,3962|false|false|false|C1552710|Bag Data Type|bag
Event|Event|Discharge Instructions|3966,3975|false|false|false|||groceries
Finding|Intellectual Product|Discharge Instructions|3983,3993|false|false|false|C1553879|applies to - HL7 Value Set and Coded Concept Property Codes|applies to
Event|Event|Discharge Instructions|4026,4029|false|false|false|||sit
Disorder|Disease or Syndrome|Discharge Instructions|4038,4041|false|false|false|C0396060|Congenital laryngeal adductor palsy|lap
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|4038,4041|false|false|false|C1870042|ACP2 protein, human|lap
Drug|Enzyme|Discharge Instructions|4038,4041|false|false|false|C1870042|ACP2 protein, human|lap
Event|Event|Discharge Instructions|4038,4041|false|false|false|||lap
Finding|Finding|Discharge Instructions|4038,4041|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Finding|Gene or Genome|Discharge Instructions|4038,4041|false|false|false|C0456170;C1412132;C1413323;C1423544;C1424863;C1425522;C2827449;C3540509;C5575443;C5890955|ACP2 gene;ACP2 wt Allele;CEBPB gene;CEBPB wt Allele;CENPJ gene;LAP3 gene;LAP3 wt Allele;Left atrial pressure;PICALM gene;PICALM wt Allele|lap
Procedure|Diagnostic Procedure|Discharge Instructions|4038,4041|false|false|false|C0031150|Laparoscopy|lap
Event|Event|Discharge Instructions|4053,4058|false|false|false|||start
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|4064,4069|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|Discharge Instructions|4064,4069|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|Discharge Instructions|4064,4069|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|Discharge Instructions|4064,4069|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|Discharge Instructions|4064,4069|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|4064,4069|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4064,4069|false|false|false|C0031765|Phototherapy|light
Finding|Daily or Recreational Activity|Discharge Instructions|4064,4078|false|false|false|C1517883|Light Exercise|light exercise
Event|Event|Discharge Instructions|4070,4078|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|4070,4078|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4070,4078|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Discharge Instructions|4093,4104|false|false|false|||comfortable
Finding|Finding|Discharge Instructions|4093,4104|false|false|false|C5546696|Feeling comfortable|comfortable
Event|Event|Discharge Instructions|4117,4121|false|false|false|||need
Event|Event|Discharge Instructions|4125,4129|false|false|false|||stay
Event|Event|Discharge Instructions|4137,4145|false|false|false|||bathtubs
Finding|Daily or Recreational Activity|Discharge Instructions|4149,4157|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|Discharge Instructions|4149,4157|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Event|Event|Discharge Instructions|4158,4163|false|false|false|||pools
Finding|Finding|Discharge Instructions|4171,4175|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|4171,4175|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|4171,4175|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Anatomy|Body Location or Region|Discharge Instructions|4187,4195|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|4187,4195|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|4187,4195|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4187,4195|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|4199,4206|false|false|false|||healing
Event|Event|Discharge Instructions|4208,4211|false|false|false|||Ask
Event|Event|Discharge Instructions|4217,4223|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|4217,4223|false|false|true|C2348314|Doctor - Title|doctor
Finding|Gene or Genome|Discharge Instructions|4245,4248|false|false|false|C1421225|TUB gene|tub
Event|Event|Discharge Instructions|4249,4254|false|false|false|||baths
Procedure|Health Care Activity|Discharge Instructions|4249,4254|false|false|false|C0150141|Bathing|baths
Event|Event|Discharge Instructions|4258,4266|false|false|false|||swimming
Finding|Daily or Recreational Activity|Discharge Instructions|4258,4266|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|Discharge Instructions|4258,4266|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Event|Event|Discharge Instructions|4276,4284|false|false|false|||exercise
Finding|Daily or Recreational Activity|Discharge Instructions|4276,4284|false|false|false|C0015259|Exercise|exercise
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4276,4284|false|false|false|C1522704|Exercise Pain Management|exercise
Event|Event|Discharge Instructions|4292,4299|false|false|false|||started
Event|Event|Discharge Instructions|4319,4322|false|false|false|||use
Event|Event|Discharge Instructions|4323,4329|false|false|false|||common
Finding|Functional Concept|Discharge Instructions|4323,4329|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Discharge Instructions|4323,4329|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Event|Event|Discharge Instructions|4331,4336|false|false|false|||sense
Finding|Organ or Tissue Function|Discharge Instructions|4331,4336|false|false|false|C0036658|Sensory perception|sense
Event|Event|Discharge Instructions|4341,4343|false|false|false|||go
Event|Event|Discharge Instructions|4371,4377|false|false|false|||resume
Finding|Behavior|Discharge Instructions|4378,4384|false|false|false|C0036864|Sex Behavior|sexual
Finding|Behavior|Discharge Instructions|4378,4393|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Finding|Individual Behavior|Discharge Instructions|4378,4393|false|false|false|C0036864;C5575036|Sex Behavior;Sexual Activity|sexual activity
Event|Activity|Discharge Instructions|4385,4393|false|false|false|C0441655|Activities|activity
Event|Event|Discharge Instructions|4385,4393|false|false|false|||activity
Finding|Daily or Recreational Activity|Discharge Instructions|4385,4393|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Finding|Finding|Discharge Instructions|4385,4393|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|activity
Event|Event|Discharge Instructions|4406,4412|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|4406,4412|false|false|false|C2348314|Doctor - Title|doctor
Event|Event|Discharge Instructions|4452,4456|false|false|false|||FEEL
Finding|Mental Process|Discharge Instructions|4452,4456|false|false|false|C1527305|Feelings|FEEL
Event|Event|Discharge Instructions|4469,4473|false|false|false|||feel
Finding|Intellectual Product|Discharge Instructions|4469,4478|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Finding|Sign or Symptom|Discharge Instructions|4469,4478|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|feel weak
Event|Event|Discharge Instructions|4474,4478|false|false|false|||weak
Finding|Intellectual Product|Discharge Instructions|4474,4478|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Finding|Sign or Symptom|Discharge Instructions|4474,4478|false|false|false|C3538976;C3714552|Feel Weak (question);Weakness|weak
Event|Event|Discharge Instructions|4483,4489|false|false|false|||washed
Event|Event|Discharge Instructions|4518,4522|false|false|false|||want
Drug|Indicator, Reagent, or Diagnostic Aid|Discharge Instructions|4527,4530|false|false|false|C4283878|Neutrophil Activation Probe Imaging Agent|nap
Event|Event|Discharge Instructions|4527,4530|false|false|false|||nap
Finding|Gene or Genome|Discharge Instructions|4527,4530|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Physiologic Function|Discharge Instructions|4527,4530|false|false|false|C0870935;C1423800|CTNNBL1 gene;Napping|nap
Finding|Intellectual Product|Discharge Instructions|4531,4536|false|false|false|C4050225|Often - answer to question|often
Finding|Gene or Genome|Discharge Instructions|4538,4544|false|false|false|C1424587|LITAF gene|Simple
Drug|Hazardous or Poisonous Substance|Discharge Instructions|4555,4562|false|false|false|C0178629|exhaust|exhaust
Finding|Sign or Symptom|Discharge Instructions|4585,4589|false|false|false|C0234233;C1442877|Sore skin;Sore to touch|sore
Disorder|Disease or Syndrome|Discharge Instructions|4585,4596|false|false|false|C0031350|Pharyngitis|sore throat
Drug|Organic Chemical|Discharge Instructions|4585,4596|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Drug|Pharmacologic Substance|Discharge Instructions|4585,4596|false|false|false|C0723402;C3244654|Sore Throat brand of Phenol;Sore Throat brand of benzocaine & menthol|sore throat
Finding|Sign or Symptom|Discharge Instructions|4585,4596|false|false|false|C0242429|Sore Throat|sore throat
Anatomy|Body Location or Region|Discharge Instructions|4590,4596|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4590,4596|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Discharge Instructions|4590,4596|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Discharge Instructions|4590,4596|false|false|false|||throat
Finding|Body Substance|Discharge Instructions|4590,4596|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Discharge Instructions|4590,4596|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Discharge Instructions|4610,4614|false|false|false|||tube
Finding|Functional Concept|Discharge Instructions|4610,4614|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Finding|Gene or Genome|Discharge Instructions|4610,4614|false|false|false|C1427122;C1719071|TUBE1 gene;Unspecified tube|tube
Anatomy|Body Location or Region|Discharge Instructions|4633,4639|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|4633,4639|false|false|false|C0031354;C0230069;C3665375|Anterior portion of neck;Pharyngeal structure;Throat|throat
Drug|Pharmacologic Substance|Discharge Instructions|4633,4639|false|false|false|C1950455|Throat Homeopathic Medication|throat
Event|Event|Discharge Instructions|4633,4639|false|false|false|||throat
Finding|Body Substance|Discharge Instructions|4633,4639|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Finding|Intellectual Product|Discharge Instructions|4633,4639|false|false|false|C1547926;C1550663|Specimen Type - Throat|throat
Event|Event|Discharge Instructions|4647,4654|false|false|false|||surgery
Finding|Finding|Discharge Instructions|4647,4654|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|4647,4654|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|4647,4654|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4647,4654|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|Discharge Instructions|4673,4680|false|false|false|||trouble
Event|Event|Discharge Instructions|4681,4694|false|false|false|||concentrating
Event|Event|Discharge Instructions|4698,4708|false|false|false|||difficulty
Finding|Finding|Discharge Instructions|4698,4708|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|Discharge Instructions|4709,4717|false|false|false|||sleeping
Event|Event|Discharge Instructions|4730,4734|false|false|false|||feel
Finding|Finding|Discharge Instructions|4735,4743|false|false|false|C2984079|Somewhat|somewhat
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|4744,4753|false|false|false|C0344315|Depressed mood|depressed
Event|Event|Discharge Instructions|4744,4753|false|false|false|||depressed
Finding|Intellectual Product|Discharge Instructions|4774,4778|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Attribute|Clinical Attribute|Discharge Instructions|4774,4787|false|false|false|C5671122||poor appetite
Finding|Intellectual Product|Discharge Instructions|4774,4787|false|false|false|C0232462;C4282406|Decrease in appetite;Poor appetite question|poor appetite
Finding|Sign or Symptom|Discharge Instructions|4774,4787|false|false|false|C0232462;C4282406|Decrease in appetite;Poor appetite question|poor appetite
Event|Event|Discharge Instructions|4779,4787|false|false|false|||appetite
Finding|Organism Function|Discharge Instructions|4779,4787|false|false|false|C0003618|Desire for food|appetite
Drug|Food|Discharge Instructions|4801,4805|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|Food
Drug|Immunologic Factor|Discharge Instructions|4801,4805|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|Food
Drug|Pharmacologic Substance|Discharge Instructions|4801,4805|false|false|false|C0016452;C3540798|Food;Food allergenic extracts|Food
Event|Event|Discharge Instructions|4801,4805|false|false|false|||Food
Event|Event|Discharge Instructions|4810,4814|false|false|false|||seem
Event|Event|Discharge Instructions|4816,4827|false|false|false|||unappealing
Event|Event|Discharge Instructions|4844,4852|false|false|false|||feelings
Finding|Intellectual Product|Discharge Instructions|4844,4852|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Finding|Mental Process|Discharge Instructions|4844,4852|false|false|false|C1527305;C4722637|Feelings;Subject's Feelings|feelings
Event|Event|Discharge Instructions|4857,4866|false|false|false|||reactions
Event|Event|Discharge Instructions|4871,4877|false|false|false|||normal
Finding|Finding|Discharge Instructions|4909,4913|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|4909,4913|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|4909,4913|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|4931,4935|false|false|false|||tell
Attribute|Clinical Attribute|Discharge Instructions|4941,4948|false|false|true|C5444295||surgeon
Anatomy|Body Location or Region|Discharge Instructions|4957,4965|false|false|false|C2338258|Cranial incision point|INCISION
Disorder|Injury or Poisoning|Discharge Instructions|4957,4965|false|false|false|C0332803|Surgical wound|INCISION
Event|Event|Discharge Instructions|4957,4965|false|false|false|||INCISION
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4957,4965|false|false|false|C0184898|Surgical incisions|INCISION
Anatomy|Body Location or Region|Discharge Instructions|4974,4982|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|4974,4982|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|4974,4982|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|4974,4982|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|4999,5002|false|false|false|||red
Finding|Finding|Discharge Instructions|4999,5002|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|Discharge Instructions|4999,5002|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Event|Event|Discharge Instructions|5030,5036|false|false|false|||normal
Event|Event|Discharge Instructions|5058,5064|false|false|false|||strips
Event|Event|Discharge Instructions|5073,5079|false|false|false|||remove
Finding|Idea or Concept|Discharge Instructions|5119,5124|false|false|false|C1547566|Paper Authorization|paper
Event|Event|Discharge Instructions|5125,5131|false|false|false|||strips
Anatomy|Body Location or Region|Discharge Instructions|5149,5157|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5149,5157|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5149,5157|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5149,5157|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5173,5177|false|false|false|||fall
Event|Event|Discharge Instructions|5225,5229|false|false|false|||wash
Drug|Substance|Discharge Instructions|5241,5249|false|false|false|C0520510|Materials|material
Event|Event|Discharge Instructions|5241,5249|false|false|false|||material
Anatomy|Body Location or Region|Discharge Instructions|5262,5270|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5262,5270|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5262,5270|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5262,5270|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5280,5286|false|false|false|||normal
Event|Event|Discharge Instructions|5290,5294|false|false|false|||feel
Event|Event|Discharge Instructions|5302,5307|false|false|false|||ridge
Finding|Functional Concept|Discharge Instructions|5302,5307|false|false|false|C0332243|Ridging|ridge
Anatomy|Body Location or Region|Discharge Instructions|5318,5326|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5318,5326|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5318,5326|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5318,5326|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5339,5341|false|false|false|||go
Finding|Intellectual Product|Discharge Instructions|5356,5362|false|false|false|C1552596;C3244286|Direct - PostalAddressUse;direct address|direct
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5363,5366|false|false|false|C0038817|Sunlight|sun
Phenomenon|Phenomenon or Process|Discharge Instructions|5363,5375|false|false|false|C1456711|Sun Exposure|sun exposure
Disorder|Injury or Poisoning|Discharge Instructions|5367,5375|false|false|false|C0274281|Injury due to exposure to external cause|exposure
Event|Event|Discharge Instructions|5367,5375|false|false|false|||exposure
Finding|Finding|Discharge Instructions|5367,5375|false|false|false|C2220266|exposure history|exposure
Phenomenon|Phenomenon or Process|Discharge Instructions|5367,5375|false|false|false|C0728853|Accident due to exposure to weather conditions|exposure
Anatomy|Body Location or Region|Discharge Instructions|5383,5391|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5383,5391|false|false|false|C0332803|Surgical wound|incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5383,5391|false|false|false|C0184898|Surgical incisions|incision
Event|Governmental or Regulatory Activity|Discharge Instructions|5392,5396|false|false|false|C1510751|Academic Research Enhancement Awards|area
Event|Event|Discharge Instructions|5407,5410|false|false|false|||use
Drug|Biomedical or Dental Material|Discharge Instructions|5415,5424|false|false|false|C0028912|Ointments|ointments
Event|Event|Discharge Instructions|5415,5424|false|false|false|||ointments
Anatomy|Body Location or Region|Discharge Instructions|5432,5440|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5432,5440|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5432,5440|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5432,5440|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5457,5461|false|false|false|||told
Event|Event|Discharge Instructions|5484,5487|false|false|false|||see
Event|Event|Discharge Instructions|5496,5502|false|false|false|||amount
Finding|Intellectual Product|Discharge Instructions|5496,5502|false|false|false|C1561574|Amount class - Amount|amount
Event|Event|Discharge Instructions|5506,5511|false|false|false|||clear
Finding|Idea or Concept|Discharge Instructions|5506,5511|false|false|false|C1550016|Remote control command - Clear|clear
Drug|Amino Acid, Peptide, or Protein|Discharge Instructions|5515,5520|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|Discharge Instructions|5515,5520|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|Discharge Instructions|5515,5520|false|false|false|||light
Finding|Finding|Discharge Instructions|5515,5520|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|Discharge Instructions|5515,5520|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|Discharge Instructions|5515,5520|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5515,5520|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5515,5520|false|false|false|C0031765|Phototherapy|light
Phenomenon|Natural Phenomenon or Process|Discharge Instructions|5515,5524|false|false|false|C0563227|Red light (physical force)|light red
Finding|Finding|Discharge Instructions|5521,5524|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|Discharge Instructions|5521,5524|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Drug|Substance|Discharge Instructions|5525,5530|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|Discharge Instructions|5525,5530|false|false|false|||fluid
Finding|Intellectual Product|Discharge Instructions|5525,5530|false|false|false|C1546638|Fluid Specimen Code|fluid
Event|Event|Discharge Instructions|5532,5540|false|false|false|||staining
Drug|Biomedical or Dental Material|Discharge Instructions|5546,5554|false|false|false|C1705365|Dressing Dosage Form|dressing
Event|Event|Discharge Instructions|5546,5554|false|false|false|||dressing
Finding|Daily or Recreational Activity|Discharge Instructions|5546,5554|false|false|false|C0518459;C1305428|Ability to dress|dressing
Finding|Finding|Discharge Instructions|5546,5554|false|false|false|C0518459;C1305428|Ability to dress|dressing
Procedure|Health Care Activity|Discharge Instructions|5546,5554|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5546,5554|false|false|false|C0152053;C0278286|Dressing of skin or wound;Dressing patient (procedure)|dressing
Event|Event|Discharge Instructions|5558,5565|false|false|false|||clothes
Event|Event|Discharge Instructions|5574,5582|false|false|false|||staining
Finding|Finding|Discharge Instructions|5574,5582|false|false|false|C1704680|Staining (finding)|staining
Procedure|Laboratory Procedure|Discharge Instructions|5574,5582|false|false|false|C0487602|Staining method|staining
Event|Event|Discharge Instructions|5586,5592|false|false|false|||severe
Finding|Finding|Discharge Instructions|5586,5592|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|5586,5592|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Discharge Instructions|5602,5606|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|5612,5619|false|false|false|C5444295||surgeon
Event|Event|Discharge Instructions|5631,5637|false|false|false|||shower
Event|Event|Discharge Instructions|5642,5647|false|false|false|||noted
Finding|Idea or Concept|Discharge Instructions|5648,5653|false|false|false|C1552828|Table Frame - above|above
Event|Event|Discharge Instructions|5655,5658|false|false|false|||ask
Event|Event|Discharge Instructions|5664,5670|false|false|false|||doctor
Finding|Intellectual Product|Discharge Instructions|5664,5670|false|false|true|C2348314|Doctor - Title|doctor
Finding|Gene or Genome|Discharge Instructions|5692,5695|false|false|false|C1421225|TUB gene|tub
Event|Event|Discharge Instructions|5696,5701|false|false|false|||baths
Procedure|Health Care Activity|Discharge Instructions|5696,5701|false|false|false|C0150141|Bathing|baths
Event|Event|Discharge Instructions|5705,5713|false|false|false|||swimming
Finding|Daily or Recreational Activity|Discharge Instructions|5705,5713|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Finding|Discharge Instructions|5705,5713|false|false|false|C0039003;C2362608|Swimming;swimming (history)|swimming
Finding|Idea or Concept|Discharge Instructions|5726,5730|false|false|false|C1552851|next - HtmlLinkType|next
Anatomy|Body Location or Region|Discharge Instructions|5748,5756|false|false|false|C2338258|Cranial incision point|incision
Disorder|Injury or Poisoning|Discharge Instructions|5748,5756|false|false|false|C0332803|Surgical wound|incision
Event|Event|Discharge Instructions|5748,5756|false|false|false|||incision
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|5748,5756|false|false|false|C0184898|Surgical incisions|incision
Event|Event|Discharge Instructions|5762,5766|false|false|false|||fade
Event|Event|Discharge Instructions|5771,5777|false|false|false|||become
Event|Event|Discharge Instructions|5784,5793|false|false|false|||prominent
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|5802,5808|false|false|false|C0021853|Intestines|BOWELS
Event|Event|Discharge Instructions|5812,5824|false|false|false|||Constipation
Finding|Sign or Symptom|Discharge Instructions|5812,5824|false|false|false|C0009806|Constipation|Constipation
Finding|Functional Concept|Discharge Instructions|5830,5836|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Intellectual Product|Discharge Instructions|5830,5836|false|false|false|C1522138;C3245511|Common Specifications in HL7 V3 Publishing;shared attribute|common
Finding|Pathologic Function|Discharge Instructions|5837,5848|false|false|false|C0879626|Adverse effects|side effect
Event|Event|Discharge Instructions|5842,5848|false|false|false|||effect
Drug|Pharmacologic Substance|Discharge Instructions|5852,5860|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|5852,5860|false|false|false|||medicine
Drug|Organic Chemical|Discharge Instructions|5870,5878|false|false|false|C0086787|Percocet|Percocet
Drug|Pharmacologic Substance|Discharge Instructions|5870,5878|false|false|false|C0086787|Percocet|Percocet
Event|Event|Discharge Instructions|5870,5878|false|false|false|||Percocet
Drug|Organic Chemical|Discharge Instructions|5882,5889|false|false|false|C0009214|codeine|codeine
Drug|Pharmacologic Substance|Discharge Instructions|5882,5889|false|false|false|C0009214|codeine|codeine
Event|Event|Discharge Instructions|5882,5889|false|false|false|||codeine
Event|Event|Discharge Instructions|5894,5900|false|false|false|||needed
Event|Event|Discharge Instructions|5910,5914|false|false|false|||take
Finding|Body Substance|Discharge Instructions|5917,5922|false|false|false|C0015733|Feces|stool
Drug|Organic Chemical|Discharge Instructions|5917,5931|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Drug|Pharmacologic Substance|Discharge Instructions|5917,5931|false|false|false|C0301470;C1154263|Stool Softener;Stool Softener brand of docusate sodium|stool softener
Event|Event|Discharge Instructions|5923,5931|false|false|false|||softener
Drug|Organic Chemical|Discharge Instructions|5942,5948|false|false|false|C0282139|Colace|Colace
Drug|Pharmacologic Substance|Discharge Instructions|5942,5948|false|false|false|C0282139|Colace|Colace
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|5954,5961|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Discharge Instructions|5954,5961|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Discharge Instructions|5954,5961|false|false|false|C0006935|capsule (pharmacologic)|capsule
Drug|Organic Chemical|Discharge Instructions|5966,5972|false|false|false|C0720654|Gentle|gentle
Drug|Pharmacologic Substance|Discharge Instructions|5966,5972|false|false|false|C0720654|Gentle|gentle
Drug|Organic Chemical|Discharge Instructions|5966,5981|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|Discharge Instructions|5966,5981|false|false|false|C0720655|Gentle Laxative|gentle laxative
Drug|Pharmacologic Substance|Discharge Instructions|5973,5981|false|false|false|C0282090|Laxatives|laxative
Event|Event|Discharge Instructions|5973,5981|false|false|false|||laxative
Drug|Food|Discharge Instructions|5991,5995|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Immunologic Factor|Discharge Instructions|5991,5995|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Pharmacologic Substance|Discharge Instructions|5991,5995|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Drug|Substance|Discharge Instructions|5991,5995|false|false|false|C0349374;C0444318;C1446647;C2702362;C2825079;C5551141;C5552693|Cow's milk;Milk Beverage;Milk Specimen;Milk antigen;Plant-Based Milk;cow milk allergenic extract|milk
Event|Event|Discharge Instructions|5991,5995|false|false|false|||milk
Finding|Body Substance|Discharge Instructions|5991,5995|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Finding|Intellectual Product|Discharge Instructions|5991,5995|false|false|false|C0026131;C1546713|Milk (body substance);Milk Specimen Code|milk
Drug|Inorganic Chemical|Discharge Instructions|6000,6008|false|false|false|C0024477|magnesium oxide|magnesia
Drug|Pharmacologic Substance|Discharge Instructions|6000,6008|false|false|false|C0024477|magnesium oxide|magnesia
Event|Event|Discharge Instructions|6000,6008|false|false|false|||magnesia
Disorder|Disease or Syndrome|Discharge Instructions|6012,6015|false|false|false|C0265246|Townes syndrome|tbs
Event|Event|Discharge Instructions|6012,6015|false|false|false|||tbs
Finding|Finding|Discharge Instructions|6012,6015|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Finding|Gene or Genome|Discharge Instructions|6012,6015|false|false|false|C1419808;C5780809;C5958753|SALL1 gene;SALL1 wt Allele;Toxicity Burden Score|tbs
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6012,6015|false|false|false|C5889868|theta-burst stimulation|tbs
Finding|Idea or Concept|Discharge Instructions|6025,6028|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|6025,6028|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|6042,6046|false|false|false|||both
Drug|Pharmacologic Substance|Discharge Instructions|6057,6066|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|6057,6066|false|false|false|||medicines
Attribute|Clinical Attribute|Discharge Instructions|6077,6089|true|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Discharge Instructions|6077,6089|false|false|false|||prescription
Finding|Intellectual Product|Discharge Instructions|6077,6089|true|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Discharge Instructions|6077,6089|true|false|false|C0033080|Prescription (procedure)|prescription
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6122,6127|false|false|false|C0021853|Intestines|bowel
Finding|Organism Function|Discharge Instructions|6122,6136|true|false|false|C0011135|Defecation|bowel movement
Event|Event|Discharge Instructions|6128,6136|false|false|false|||movement
Finding|Organism Function|Discharge Instructions|6128,6136|true|false|false|C0026649|Movement|movement
Finding|Intellectual Product|Discharge Instructions|6141,6150|false|false|false|C2984058|Have Pain|have pain
Attribute|Clinical Attribute|Discharge Instructions|6146,6150|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6146,6150|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6146,6150|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6146,6150|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|6152,6158|false|false|false|||moving
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|6164,6170|false|false|false|C0021853|Intestines|bowels
Event|Event|Discharge Instructions|6172,6176|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|6182,6189|false|false|false|C5444295||surgeon
Event|Activity|Discharge Instructions|6204,6214|false|false|false|C3241922|Operation Activity|operations
Event|Event|Discharge Instructions|6204,6214|false|false|false|||operations
Finding|Functional Concept|Discharge Instructions|6204,6214|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Finding|Intellectual Product|Discharge Instructions|6204,6214|false|false|false|C0038895;C3244305;C3244306|ActInformationPrivacyReason - operations;HL7PublishingSubSection - operations;Surgical aspects|operations
Event|Event|Discharge Instructions|6216,6224|false|false|false|||diarrhea
Finding|Finding|Discharge Instructions|6216,6224|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|6216,6224|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|Discharge Instructions|6229,6234|false|false|false|||occur
Event|Event|Discharge Instructions|6248,6256|false|false|false|||diarrhea
Finding|Finding|Discharge Instructions|6248,6256|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|Discharge Instructions|6248,6256|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Drug|Organic Chemical|Discharge Instructions|6269,6282|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|Discharge Instructions|6269,6282|false|false|false|C0718564|Anti-Diarrhea|anti-diarrhea
Drug|Pharmacologic Substance|Discharge Instructions|6283,6292|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Discharge Instructions|6283,6292|false|false|false|||medicines
Drug|Substance|Discharge Instructions|6311,6317|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|6311,6317|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|6311,6317|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6311,6317|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Discharge Instructions|6322,6325|false|false|false|||see
Event|Event|Discharge Instructions|6332,6336|false|false|false|||goes
Event|Event|Discharge Instructions|6358,6360|false|false|false|||go
Event|Event|Discharge Instructions|6374,6380|false|false|false|||severe
Finding|Finding|Discharge Instructions|6374,6380|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|6374,6380|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|6389,6397|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|Discharge Instructions|6389,6397|false|false|false|C0231218;C0557911;C2987492|Feel Ill Question;Feeling bad emotionally;Malaise|feel ill
Finding|Sign or Symptom|Discharge Instructions|6394,6397|false|false|false|C0231218|Malaise|ill
Event|Event|Discharge Instructions|6406,6410|false|false|false|||call
Attribute|Clinical Attribute|Discharge Instructions|6416,6423|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|Discharge Instructions|6427,6431|false|false|false|C2598155||PAIN
Event|Event|Discharge Instructions|6427,6431|false|false|false|||PAIN
Finding|Functional Concept|Discharge Instructions|6427,6431|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Finding|Sign or Symptom|Discharge Instructions|6427,6431|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|PAIN
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6427,6442|false|false|false|C0002766|Pain management (procedure)|PAIN MANAGEMENT
Event|Event|Discharge Instructions|6432,6442|false|false|false|||MANAGEMENT
Event|Occupational Activity|Discharge Instructions|6432,6442|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|MANAGEMENT
Procedure|Health Care Activity|Discharge Instructions|6432,6442|false|false|false|C0376636|Disease Management|MANAGEMENT
Event|Event|Discharge Instructions|6452,6458|false|false|false|||normal
Event|Event|Discharge Instructions|6462,6466|false|false|false|||feel
Event|Event|Discharge Instructions|6472,6482|false|false|false|||discomfort
Finding|Sign or Symptom|Discharge Instructions|6472,6482|false|false|false|C2364135|Discomfort|discomfort
Attribute|Clinical Attribute|Discharge Instructions|6483,6487|false|true|false|C2598155||pain
Event|Event|Discharge Instructions|6483,6487|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6483,6487|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6483,6487|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|Discharge Instructions|6498,6507|false|false|false|C0000726|Abdomen|abdominal
Event|Event|Discharge Instructions|6509,6516|false|false|false|||surgery
Finding|Finding|Discharge Instructions|6509,6516|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|Discharge Instructions|6509,6516|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|Discharge Instructions|6509,6516|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|6509,6516|false|false|false|C0543467|Operative Surgical Procedures|surgery
Attribute|Clinical Attribute|Discharge Instructions|6523,6527|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6523,6527|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6523,6527|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6523,6527|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Intellectual Product|Discharge Instructions|6531,6536|false|false|false|C4050225|Often - answer to question|often
Event|Event|Discharge Instructions|6537,6546|false|false|false|||described
Event|Event|Discharge Instructions|6551,6559|false|false|false|||soreness
Finding|Sign or Symptom|Discharge Instructions|6551,6559|false|false|false|C0234233|Sore to touch|soreness
Attribute|Clinical Attribute|Discharge Instructions|6570,6574|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6570,6574|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6570,6574|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6570,6574|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|6586,6592|false|false|false|||better
Finding|Idea or Concept|Discharge Instructions|6586,6592|false|false|false|C1550462|Observation Interpretation - better|better
Finding|Idea or Concept|Discharge Instructions|6593,6596|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|6593,6596|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Idea or Concept|Discharge Instructions|6600,6603|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Discharge Instructions|6600,6603|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Discharge Instructions|6612,6616|false|false|false|||find
Attribute|Clinical Attribute|Discharge Instructions|6621,6625|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6621,6625|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6621,6625|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6621,6625|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|6638,6643|false|false|false|||worse
Finding|Finding|Discharge Instructions|6638,6643|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|6638,6643|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|6655,6661|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|6670,6677|false|false|false|||contact
Attribute|Clinical Attribute|Discharge Instructions|6683,6690|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|Discharge Instructions|6712,6724|false|false|false|C5886759|Prescription (attribute)|prescription
Event|Event|Discharge Instructions|6712,6724|false|false|false|||prescription
Finding|Intellectual Product|Discharge Instructions|6712,6724|false|false|false|C1521941|prescription document|prescription
Procedure|Health Care Activity|Discharge Instructions|6712,6724|false|false|false|C0033080|Prescription (procedure)|prescription
Attribute|Clinical Attribute|Discharge Instructions|6735,6742|false|false|false|C5444295||surgeon
Attribute|Clinical Attribute|Discharge Instructions|6747,6751|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6747,6751|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6747,6751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6747,6751|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Pharmacologic Substance|Discharge Instructions|6753,6761|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6753,6761|false|false|false|||medicine
Event|Event|Discharge Instructions|6765,6769|false|false|false|||take
Finding|Functional Concept|Discharge Instructions|6770,6778|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Discharge Instructions|6773,6778|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|6773,6778|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Discharge Instructions|6786,6795|false|false|false|||important
Event|Event|Discharge Instructions|6799,6803|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|6809,6817|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6809,6817|false|false|false|||medicine
Event|Event|Discharge Instructions|6822,6830|false|false|false|||directed
Event|Event|Discharge Instructions|6842,6846|false|false|false|||take
Event|Event|Discharge Instructions|6871,6881|false|false|false|||prescribed
Event|Event|Discharge Instructions|6890,6894|false|false|false|||take
Drug|Pharmacologic Substance|Discharge Instructions|6901,6909|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6901,6909|false|false|false|||medicine
Finding|Intellectual Product|Discharge Instructions|6913,6921|false|false|false|C3241998|one time|one time
Finding|Finding|Discharge Instructions|6917,6921|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|6917,6921|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|6917,6921|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Discharge Instructions|6927,6937|false|false|false|||prescribed
Attribute|Clinical Attribute|Discharge Instructions|6946,6950|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|6946,6950|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|6946,6950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|6946,6950|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|6946,6959|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|6946,6959|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|6946,6959|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|6951,6959|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|6951,6959|false|false|false|||medicine
Event|Event|Discharge Instructions|6965,6969|false|false|false|||work
Finding|Idea or Concept|Discharge Instructions|6970,6976|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|6984,6988|false|false|false|||take
Attribute|Clinical Attribute|Discharge Instructions|7005,7009|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7005,7009|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7005,7009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7005,7009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7010,7014|false|false|false|||gets
Event|Event|Discharge Instructions|7019,7025|false|false|false|||severe
Finding|Finding|Discharge Instructions|7019,7025|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|7019,7025|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Attribute|Clinical Attribute|Discharge Instructions|7057,7061|true|false|false|C2598155||pain
Event|Event|Discharge Instructions|7057,7061|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7057,7061|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7057,7061|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7069,7073|false|false|false|||okay
Event|Event|Discharge Instructions|7077,7081|false|false|false|||skip
Event|Event|Discharge Instructions|7084,7088|false|false|false|||dose
Attribute|Clinical Attribute|Discharge Instructions|7093,7097|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7093,7097|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7093,7097|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7093,7097|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Hazardous or Poisonous Substance|Discharge Instructions|7093,7106|false|false|false|C0002771|Analgesics|pain medicine
Drug|Organic Chemical|Discharge Instructions|7093,7106|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|7093,7106|false|false|false|C0002771|Analgesics|pain medicine
Drug|Pharmacologic Substance|Discharge Instructions|7098,7106|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Discharge Instructions|7098,7106|false|false|false|||medicine
Event|Event|Discharge Instructions|7115,7125|false|false|false|||experience
Event|Event|Discharge Instructions|7155,7162|false|false|false|||contact
Attribute|Clinical Attribute|Discharge Instructions|7169,7176|false|false|false|C5444295||surgeon
Finding|Finding|Discharge Instructions|7180,7185|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Gene or Genome|Discharge Instructions|7180,7185|false|false|false|C1444775;C1539835;C3890003|SPEN gene;SPEN wt Allele;Sharp sensation quality|sharp
Finding|Sign or Symptom|Discharge Instructions|7180,7190|false|false|false|C0455270|Sharp pain|sharp pain
Attribute|Clinical Attribute|Discharge Instructions|7186,7190|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7186,7190|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7186,7190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7186,7190|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Discharge Instructions|7198,7204|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Discharge Instructions|7198,7204|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Finding|Discharge Instructions|7198,7209|false|false|false|C0278140;C4050465;C4521229|Neck Pain Score 6;Severe Extremity Pain;Severe pain|severe pain
Attribute|Clinical Attribute|Discharge Instructions|7205,7209|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7205,7209|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7205,7209|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7205,7209|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7215,7220|false|false|false|||lasts
Event|Event|Discharge Instructions|7229,7234|false|false|false|||hours
Attribute|Clinical Attribute|Discharge Instructions|7237,7241|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7237,7241|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7237,7241|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7237,7241|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7258,7263|false|false|false|||worse
Finding|Finding|Discharge Instructions|7258,7263|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Idea or Concept|Discharge Instructions|7258,7263|false|false|false|C1457868;C1550463|Observation Interpretation - worse;Worse|worse
Finding|Finding|Discharge Instructions|7269,7273|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|7269,7273|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|7269,7273|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Attribute|Clinical Attribute|Discharge Instructions|7276,7280|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7276,7280|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7276,7280|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7276,7280|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Discharge Instructions|7281,7292|false|false|false|||accompanied
Finding|Finding|Discharge Instructions|7296,7301|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Discharge Instructions|7296,7301|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|Discharge Instructions|7331,7337|false|false|false|||change
Finding|Functional Concept|Discharge Instructions|7331,7337|false|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|7331,7337|false|false|false|C4319952|Change - procedure|change
Finding|Functional Concept|Discharge Instructions|7331,7340|false|false|false|C0392747|Changing|change in
Event|Event|Discharge Instructions|7341,7347|false|false|false|||nature
Finding|Functional Concept|Discharge Instructions|7341,7347|false|false|false|C0349590;C1262865|Nature;Natures|nature
Finding|Idea or Concept|Discharge Instructions|7341,7347|false|false|false|C0349590;C1262865|Nature;Natures|nature
Event|Event|Discharge Instructions|7351,7358|false|false|false|||quality
Attribute|Clinical Attribute|Discharge Instructions|7367,7371|false|false|false|C2598155||pain
Event|Event|Discharge Instructions|7367,7371|false|false|false|||pain
Finding|Functional Concept|Discharge Instructions|7367,7371|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|7367,7371|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|Medications|7389,7393|false|false|false|||Take
Drug|Pharmacologic Substance|Medications|7402,7411|false|false|false|C0013227|Pharmaceutical Preparations|medicines
Event|Event|Medications|7402,7411|false|false|false|||medicines
Event|Activity|Medications|7435,7444|false|false|false|C3241922|Operation Activity|operation
Event|Event|Medications|7435,7444|false|false|false|||operation
Procedure|Machine Activity|Medications|7435,7444|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Procedure|Therapeutic or Preventive Procedure|Medications|7435,7444|false|false|false|C0543467;C1880161|Computer Operation;Operative Surgical Procedures|operation
Event|Event|Medications|7491,7495|false|false|false|||told
Event|Event|Medications|7527,7536|false|false|false|||questions
Drug|Pharmacologic Substance|Medications|7548,7556|false|false|false|C0013227|Pharmaceutical Preparations|medicine
Event|Event|Medications|7548,7556|false|false|false|||medicine
Event|Event|Medications|7560,7564|false|false|false|||take
Procedure|Health Care Activity|Medications|7576,7580|false|false|false|C1515187|Take|take
Event|Event|Medications|7589,7593|false|false|false|||call
Attribute|Clinical Attribute|Medications|7599,7606|false|false|false|C5444295||surgeon
Procedure|Health Care Activity|Medications|7611,7619|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Medications|7620,7632|false|false|false|C3263700||Instructions
Event|Event|Medications|7620,7632|false|false|false|||Instructions
Finding|Intellectual Product|Medications|7620,7632|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

