 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|27,31
No|32,34
:|34,35
_|38,39
_|39,40
_|40,41
<EOL>|41,42
<EOL>|43,44
Admission|44,53
Date|54,58
:|58,59
_|61,62
_|62,63
_|63,64
Discharge|78,87
Date|88,92
:|92,93
_|96,97
_|97,98
_|98,99
<EOL>|99,100
<EOL>|101,102
Date|102,106
of|107,109
Birth|110,115
:|115,116
_|118,119
_|119,120
_|120,121
Sex|134,137
:|137,138
M|141,142
<EOL>|142,143
<EOL>|144,145
Service|145,152
:|152,153
MEDICINE|154,162
<EOL>|162,163
<EOL>|164,165
No|177,179
Known|180,185
Allergies|186,195
/|196,197
Adverse|198,205
Drug|206,210
Reactions|211,220
<EOL>|220,221
<EOL>|222,223
Attending|223,232
:|232,233
_|234,235
_|235,236
_|236,237
<EOL>|237,238
<EOL>|239,240
Epistaxis|257,266
<EOL>|266,267
<EOL>|268,269
Major|269,274
Surgical|275,283
or|284,286
Invasive|287,295
Procedure|296,305
:|305,306
<EOL>|306,307
None|307,311
<EOL>|311,312
<EOL>|312,313
<EOL>|314,315
Mr.|343,346
_|347,348
_|348,349
_|349,350
is|351,353
an|354,356
_|357,358
_|358,359
_|359,360
with|361,365
history|366,373
of|374,376
AAA|377,380
s|381,382
/|382,383
p|383,384
repair|385,391
<EOL>|392,393
complicated|393,404
by|405,407
MI|408,410
,|410,411
hypertension|412,424
,|424,425
and|426,429
hyperlipidemia|430,444
who|445,448
presents|449,457
<EOL>|458,459
upon|459,463
transfer|464,472
from|473,477
outside|478,485
hospital|486,494
with|495,499
nasal|500,505
fractures|506,515
and|516,519
<EOL>|520,521
epistaxis|521,530
secondary|531,540
to|541,543
fall|544,548
.|548,549
The|550,553
patient|554,561
reports|562,569
that|570,574
he|575,577
was|578,581
at|582,584
<EOL>|585,586
the|586,589
_|590,591
_|591,592
_|592,593
earlier|594,601
this|602,606
afternoon|607,616
.|616,617
While|618,623
coughing|624,632
,|632,633
he|634,636
tripped|637,644
<EOL>|645,646
on|646,648
the|649,652
curb|653,657
and|658,661
suffered|662,670
trauma|671,677
to|678,680
his|681,684
face|685,689
.|689,690
He|691,693
had|694,697
no|698,700
loss|701,705
of|706,708
<EOL>|709,710
consciousness|710,723
.|723,724
However|725,732
,|732,733
he|734,736
had|737,740
a|741,742
persistent|743,753
nosebleed|754,763
and|764,767
<EOL>|768,769
appeared|769,777
to|778,780
have|781,785
some|786,790
trauma|791,797
to|798,800
his|801,804
face|805,809
,|809,810
thus|811,815
was|816,819
transferred|820,831
<EOL>|832,833
to|833,835
_|836,837
_|837,838
_|838,839
for|840,843
further|844,851
care|852,856
.|856,857
There|858,863
,|863,864
a|865,866
CT|867,869
scan|870,874
of|875,877
<EOL>|878,879
the|879,882
head|883,887
,|887,888
neck|889,893
,|893,894
and|895,898
face|899,903
were|904,908
remarkable|909,919
for|920,923
a|924,925
nasal|926,931
bone|932,936
and|937,940
<EOL>|941,942
septal|942,948
fracture|949,957
.|957,958
Given|959,964
persistent|965,975
epistaxis|976,985
,|985,986
bilateral|987,996
<EOL>|997,998
RhinoRockets|998,1010
were|1011,1015
placed|1016,1022
.|1022,1023
He|1024,1026
had|1027,1030
a|1031,1032
small|1033,1038
abrasion|1039,1047
to|1048,1050
the|1051,1054
bridge|1055,1061
<EOL>|1062,1063
of|1063,1065
his|1066,1069
nose|1070,1074
which|1075,1080
was|1081,1084
not|1085,1088
closed|1089,1095
.|1095,1096
Bleeding|1097,1105
was|1106,1109
well|1110,1114
controlled|1115,1125
.|1125,1126
<EOL>|1127,1128
While|1128,1133
in|1134,1136
the|1137,1140
OSH|1141,1144
ED|1145,1147
,|1147,1148
he|1149,1151
had|1152,1155
an|1156,1158
episode|1159,1166
of|1167,1169
nausea|1170,1176
and|1177,1180
coughed|1181,1188
up|1189,1191
<EOL>|1192,1193
some|1193,1197
blood|1198,1203
.|1203,1204
At|1205,1207
that|1208,1212
time|1213,1217
,|1217,1218
he|1219,1221
began|1222,1227
to|1228,1230
feel|1231,1235
lightheaded|1236,1247
and|1248,1251
was|1252,1255
<EOL>|1256,1257
noted|1257,1262
to|1263,1265
be|1266,1268
hypotensive|1269,1280
and|1281,1284
bradycardic|1285,1296
.|1296,1297
Per|1298,1301
report|1302,1308
,|1308,1309
he|1310,1312
had|1313,1316
a|1317,1318
<EOL>|1319,1320
brief|1320,1325
loss|1326,1330
of|1331,1333
consciousness|1334,1347
,|1347,1348
though|1349,1355
quickly|1356,1363
returned|1364,1372
to|1373,1375
his|1376,1379
<EOL>|1380,1381
baseline|1381,1389
.|1389,1390
His|1391,1394
family|1395,1401
noted|1402,1407
that|1408,1412
his|1413,1416
eyes|1417,1421
rolled|1422,1428
back|1429,1433
into|1434,1438
his|1439,1442
<EOL>|1443,1444
head|1444,1448
.|1448,1449
The|1450,1453
patient|1454,1461
recalls|1462,1469
the|1470,1473
event|1474,1479
and|1480,1483
denies|1484,1490
post-event|1491,1501
<EOL>|1502,1503
confusion|1503,1512
.|1512,1513
He|1514,1516
had|1517,1520
no|1521,1523
further|1524,1531
episodes|1532,1540
of|1541,1543
syncope|1544,1551
or|1552,1554
hemodynamic|1555,1566
<EOL>|1567,1568
changes|1568,1575
.|1575,1576
Given|1578,1583
the|1584,1587
syncopal|1588,1596
event|1597,1602
and|1603,1606
epistaxis|1607,1616
,|1616,1617
the|1618,1621
patient|1622,1629
<EOL>|1630,1631
was|1631,1634
transferred|1635,1646
for|1647,1650
further|1651,1658
care|1659,1663
.|1663,1664
<EOL>|1664,1665
<EOL>|1665,1666
In|1666,1668
the|1669,1672
ED|1673,1675
,|1675,1676
initial|1677,1684
vital|1685,1690
signs|1691,1696
98.9|1697,1701
92|1702,1704
140|1705,1708
/|1708,1709
77|1709,1711
18|1712,1714
100|1715,1718
%|1718,1719
/|1719,1720
RA|1720,1722
.|1722,1723
Labs|1724,1728
<EOL>|1729,1730
were|1730,1734
notable|1735,1742
for|1743,1746
WBC|1747,1750
11.3|1751,1755
(|1756,1757
91|1757,1759
%|1759,1760
N|1760,1761
)|1761,1762
,|1762,1763
H|1764,1765
/|1765,1766
H|1766,1767
14.1|1768,1772
/|1772,1773
40|1773,1775
.|1775,1776
2|1776,1777
,|1777,1778
plt|1779,1782
147|1783,1786
,|1786,1787
BUN|1788,1791
/|1791,1792
Cr|1792,1794
<EOL>|1795,1796
36|1796,1798
/|1798,1799
1.5|1799,1802
.|1802,1803
HCTs|1804,1808
were|1809,1813
repeated|1814,1822
which|1823,1828
were|1829,1833
stable|1834,1840
.|1840,1841
A|1842,1843
urinalysis|1844,1854
was|1855,1858
<EOL>|1859,1860
negative|1860,1868
.|1868,1869
A|1870,1871
CXR|1872,1875
demonstrated|1876,1888
a|1889,1890
focal|1891,1896
consolidation|1897,1910
at|1911,1913
the|1914,1917
left|1918,1922
<EOL>|1923,1924
lung|1924,1928
base|1929,1933
,|1933,1934
possibly|1935,1943
representing|1944,1956
aspiration|1957,1967
or|1968,1970
developing|1971,1981
<EOL>|1982,1983
pneumonia|1983,1992
.|1992,1993
The|1994,1997
patient|1998,2005
was|2006,2009
given|2010,2015
Tdap|2016,2020
,|2020,2021
amoxicillin|2022,2033
-|2033,2034
clavulanate|2034,2045
<EOL>|2046,2047
for|2047,2050
antibiotic|2051,2061
prophylaxis|2062,2073
,|2073,2074
ondansetron|2075,2086
,|2086,2087
500cc|2088,2093
NS|2094,2096
,|2096,2097
and|2098,2101
<EOL>|2102,2103
metoprolol|2103,2113
tartrate|2114,2122
50mg|2123,2127
.|2127,2128
Clopidogrel|2129,2140
was|2141,2144
held|2145,2149
.|2149,2150
<EOL>|2150,2151
<EOL>|2152,2153
MI|2175,2177
after|2178,2183
AAA|2184,2187
repair|2188,2194
when|2195,2199
he|2200,2202
was|2203,2206
_|2207,2208
_|2208,2209
_|2209,2210
y|2211,2212
/|2212,2213
o|2213,2214
<EOL>|2214,2215
HTN|2215,2218
<EOL>|2218,2219
Hypercholesterolemia|2219,2239
<EOL>|2239,2240
<EOL>|2241,2242
:|2256,2257
<EOL>|2257,2258
_|2258,2259
_|2259,2260
_|2260,2261
<EOL>|2261,2262
:|2276,2277
<EOL>|2277,2278
Patient|2278,2285
is|2286,2288
unaware|2289,2296
of|2297,2299
a|2300,2301
family|2302,2308
history|2309,2316
of|2317,2319
bleeding|2320,2328
diathesis|2329,2338
.|2338,2339
<EOL>|2339,2340
<EOL>|2340,2341
<EOL>|2342,2343
ADMISSION|2358,2367
:|2367,2368
<EOL>|2368,2369
VS|2369,2371
:|2371,2372
98.5|2373,2377
142|2378,2381
/|2381,2382
65|2382,2384
95|2385,2387
18|2388,2390
98RA|2391,2395
<EOL>|2395,2396
GENERAL|2396,2403
:|2403,2404
Alert|2405,2410
,|2410,2411
oriented|2412,2420
,|2420,2421
no|2422,2424
acute|2425,2430
distress|2431,2439
<EOL>|2441,2442
HEENT|2442,2447
:|2447,2448
Sclerae|2449,2456
anicteric|2457,2466
,|2466,2467
MMM|2468,2471
,|2471,2472
oropharynx|2473,2483
clear|2484,2489
,|2489,2490
bruising|2491,2499
under|2500,2505
<EOL>|2506,2507
both|2507,2511
eyes|2512,2516
,|2516,2517
swollen|2518,2525
nose|2526,2530
with|2531,2535
mild|2536,2540
tenderness|2541,2551
,|2551,2552
RhinoRockets|2553,2565
in|2566,2568
<EOL>|2569,2570
place|2570,2575
<EOL>|2577,2578
NECK|2578,2582
:|2582,2583
Supple|2584,2590
,|2590,2591
without|2592,2599
LAD|2600,2603
<EOL>|2605,2606
RESP|2606,2610
:|2610,2611
Generally|2612,2621
CTA|2622,2625
bilaterally|2626,2637
<EOL>|2639,2640
CV|2640,2642
:|2642,2643
RRR|2644,2647
,|2647,2648
(|2649,2650
+|2650,2651
)|2651,2652
S1|2652,2654
/|2654,2655
S2|2655,2657
no|2658,2660
m|2661,2662
/|2662,2663
r|2663,2664
/|2664,2665
g|2665,2666
<EOL>|2668,2669
ABD|2669,2672
:|2672,2673
Soft|2674,2678
,|2678,2679
non-tender|2680,2690
,|2690,2691
non-distended|2692,2705
<EOL>|2705,2706
GU|2706,2708
:|2708,2709
Deferred|2710,2718
<EOL>|2719,2720
EXT|2720,2723
:|2723,2724
Warm|2725,2729
,|2729,2730
well|2731,2735
perfused|2736,2744
,|2744,2745
2|2746,2747
+|2747,2748
pulses|2749,2755
,|2755,2756
no|2757,2759
clubbing|2760,2768
,|2768,2769
cyanosis|2770,2778
or|2779,2781
<EOL>|2782,2783
edema|2783,2788
<EOL>|2790,2791
NEURO|2791,2796
:|2796,2797
CN|2798,2800
II|2801,2803
-|2803,2804
XII|2804,2807
grossly|2808,2815
intact|2816,2822
,|2822,2823
motor|2824,2829
function|2830,2838
grossly|2839,2846
normal|2847,2853
<EOL>|2853,2854
SKIN|2854,2858
:|2858,2859
No|2860,2862
excoriations|2863,2875
or|2876,2878
rash|2879,2883
.|2883,2884
<EOL>|2884,2885
<EOL>|2885,2886
DISCHARGE|2886,2895
:|2895,2896
<EOL>|2896,2897
VS|2897,2899
:|2899,2900
98.4|2901,2905
125|2906,2909
/|2909,2910
55|2910,2912
73|2913,2915
18|2916,2918
94RA|2919,2923
<EOL>|2923,2924
GENERAL|2924,2931
:|2931,2932
Alert|2933,2938
,|2938,2939
oriented|2940,2948
,|2948,2949
no|2950,2952
acute|2953,2958
distress|2959,2967
<EOL>|2969,2970
HEENT|2970,2975
:|2975,2976
Sclerae|2977,2984
anicteric|2985,2994
,|2994,2995
MMM|2996,2999
,|2999,3000
oropharynx|3001,3011
clear|3012,3017
,|3017,3018
bruising|3019,3027
under|3028,3033
<EOL>|3034,3035
both|3035,3039
eyes|3040,3044
,|3044,3045
swollen|3046,3053
nose|3054,3058
with|3059,3063
mild|3064,3068
tenderness|3069,3079
,|3079,3080
RhinoRockets|3081,3093
in|3094,3096
<EOL>|3097,3098
place|3098,3103
<EOL>|3105,3106
NECK|3106,3110
:|3110,3111
Supple|3112,3118
,|3118,3119
without|3120,3127
LAD|3128,3131
<EOL>|3133,3134
RESP|3134,3138
:|3138,3139
Generally|3140,3149
CTA|3150,3153
bilaterally|3154,3165
<EOL>|3167,3168
CV|3168,3170
:|3170,3171
RRR|3172,3175
,|3175,3176
(|3177,3178
+|3178,3179
)|3179,3180
S1|3180,3182
/|3182,3183
S2|3183,3185
no|3186,3188
m|3189,3190
/|3190,3191
r|3191,3192
/|3192,3193
g|3193,3194
<EOL>|3196,3197
ABD|3197,3200
:|3200,3201
Soft|3202,3206
,|3206,3207
non-tender|3208,3218
,|3218,3219
non-distended|3220,3233
<EOL>|3233,3234
GU|3234,3236
:|3236,3237
Deferred|3238,3246
<EOL>|3247,3248
EXT|3248,3251
:|3251,3252
Warm|3253,3257
,|3257,3258
well|3259,3263
perfused|3264,3272
,|3272,3273
2|3274,3275
+|3275,3276
pulses|3277,3283
,|3283,3284
no|3285,3287
clubbing|3288,3296
,|3296,3297
cyanosis|3298,3306
or|3307,3309
<EOL>|3310,3311
edema|3311,3316
<EOL>|3318,3319
NEURO|3319,3324
:|3324,3325
CN|3326,3328
II|3329,3331
-|3331,3332
XII|3332,3335
grossly|3336,3343
intact|3344,3350
,|3350,3351
motor|3352,3357
function|3358,3366
grossly|3367,3374
normal|3375,3381
<EOL>|3381,3382
SKIN|3382,3386
:|3386,3387
No|3388,3390
excoriations|3391,3403
or|3404,3406
rash|3407,3411
.|3411,3412
<EOL>|3412,3413
<EOL>|3414,3415
Pertinent|3415,3424
Results|3425,3432
:|3432,3433
<EOL>|3433,3434
ADMISSION|3434,3443
:|3443,3444
<EOL>|3444,3445
_|3445,3446
_|3446,3447
_|3447,3448
08|3449,3451
:|3451,3452
15PM|3452,3456
BLOOD|3457,3462
WBC|3463,3466
-|3466,3467
11|3467,3469
.|3469,3470
3|3470,3471
*|3471,3472
RBC|3473,3476
-|3476,3477
4|3477,3478
.|3478,3479
30|3479,3481
*|3481,3482
Hgb|3483,3486
-|3486,3487
14.1|3487,3491
Hct|3492,3495
-|3495,3496
40.2|3496,3500
<EOL>|3501,3502
MCV|3502,3505
-|3505,3506
93|3506,3508
MCH|3509,3512
-|3512,3513
32|3513,3515
.|3515,3516
8|3516,3517
*|3517,3518
MCHC|3519,3523
-|3523,3524
35|3524,3526
.|3526,3527
1|3527,3528
*|3528,3529
RDW|3530,3533
-|3533,3534
12.8|3534,3538
Plt|3539,3542
_|3543,3544
_|3544,3545
_|3545,3546
<EOL>|3546,3547
_|3547,3548
_|3548,3549
_|3549,3550
08|3551,3553
:|3553,3554
15PM|3554,3558
BLOOD|3559,3564
Neuts|3565,3570
-|3570,3571
91|3571,3573
.|3573,3574
1|3574,3575
*|3575,3576
Lymphs|3577,3583
-|3583,3584
4|3584,3585
.|3585,3586
7|3586,3587
*|3587,3588
Monos|3589,3594
-|3594,3595
3.8|3595,3598
Eos|3599,3602
-|3602,3603
0.3|3603,3606
<EOL>|3607,3608
Baso|3608,3612
-|3612,3613
0.1|3613,3616
<EOL>|3616,3617
_|3617,3618
_|3618,3619
_|3619,3620
08|3621,3623
:|3623,3624
15PM|3624,3628
BLOOD|3629,3634
_|3635,3636
_|3636,3637
_|3637,3638
PTT|3639,3642
-|3642,3643
26.8|3643,3647
_|3648,3649
_|3649,3650
_|3650,3651
<EOL>|3651,3652
_|3652,3653
_|3653,3654
_|3654,3655
08|3656,3658
:|3658,3659
15PM|3659,3663
BLOOD|3664,3669
Glucose|3670,3677
-|3677,3678
159|3678,3681
*|3681,3682
UreaN|3683,3688
-|3688,3689
36|3689,3691
*|3691,3692
Creat|3693,3698
-|3698,3699
1|3699,3700
.|3700,3701
5|3701,3702
*|3702,3703
Na|3704,3706
-|3706,3707
141|3707,3710
<EOL>|3711,3712
K|3712,3713
-|3713,3714
4.1|3714,3717
Cl|3718,3720
-|3720,3721
106|3721,3724
HCO3|3725,3729
-|3729,3730
21|3730,3732
*|3732,3733
AnGap|3734,3739
-|3739,3740
18|3740,3742
<EOL>|3742,3743
_|3743,3744
_|3744,3745
_|3745,3746
06|3747,3749
:|3749,3750
03AM|3750,3754
BLOOD|3755,3760
CK|3761,3763
(|3763,3764
CPK|3764,3767
)|3767,3768
-|3768,3769
594|3769,3772
*|3772,3773
<EOL>|3773,3774
<EOL>|3774,3775
CARDIAC|3775,3782
MARKER|3783,3789
TREND|3790,3795
:|3795,3796
<EOL>|3796,3797
_|3797,3798
_|3798,3799
_|3799,3800
07|3801,3803
:|3803,3804
45AM|3804,3808
BLOOD|3809,3814
cTropnT|3815,3822
-|3822,3823
0|3823,3824
.|3824,3825
04|3825,3827
*|3827,3828
<EOL>|3828,3829
_|3829,3830
_|3830,3831
_|3831,3832
06|3833,3835
:|3835,3836
03AM|3836,3840
BLOOD|3841,3846
CK|3847,3849
-|3849,3850
MB|3850,3852
-|3852,3853
36|3853,3855
*|3855,3856
MB|3857,3859
Indx|3860,3864
-|3864,3865
6|3865,3866
.|3866,3867
1|3867,3868
*|3868,3869
cTropnT|3870,3877
-|3877,3878
0|3878,3879
.|3879,3880
57|3880,3882
*|3882,3883
<EOL>|3883,3884
_|3884,3885
_|3885,3886
_|3886,3887
03|3888,3890
:|3890,3891
03PM|3891,3895
BLOOD|3896,3901
CK|3902,3904
-|3904,3905
MB|3905,3907
-|3907,3908
23|3908,3910
*|3910,3911
MB|3912,3914
Indx|3915,3919
-|3919,3920
4.2|3920,3923
cTropnT|3924,3931
-|3931,3932
0|3932,3933
.|3933,3934
89|3934,3936
*|3936,3937
<EOL>|3937,3938
_|3938,3939
_|3939,3940
_|3940,3941
05|3942,3944
:|3944,3945
59AM|3945,3949
BLOOD|3950,3955
CK|3956,3958
-|3958,3959
MB|3959,3961
-|3961,3962
8|3962,3963
cTropnT|3964,3971
-|3971,3972
1|3972,3973
.|3973,3974
28|3974,3976
*|3976,3977
<EOL>|3977,3978
_|3978,3979
_|3979,3980
_|3980,3981
01|3982,3984
:|3984,3985
16PM|3985,3989
BLOOD|3990,3995
CK|3996,3998
-|3998,3999
MB|3999,4001
-|4001,4002
5|4002,4003
cTropnT|4004,4011
-|4011,4012
1|4012,4013
.|4013,4014
29|4014,4016
*|4016,4017
<EOL>|4017,4018
_|4018,4019
_|4019,4020
_|4020,4021
06|4022,4024
:|4024,4025
10AM|4025,4029
BLOOD|4030,4035
CK|4036,4038
-|4038,4039
MB|4039,4041
-|4041,4042
4|4042,4043
cTropnT|4044,4051
-|4051,4052
1|4052,4053
.|4053,4054
48|4054,4056
*|4056,4057
<EOL>|4057,4058
_|4058,4059
_|4059,4060
_|4060,4061
07|4062,4064
:|4064,4065
28AM|4065,4069
BLOOD|4070,4075
CK|4076,4078
-|4078,4079
MB|4079,4081
-|4081,4082
2|4082,4083
cTropnT|4084,4091
-|4091,4092
1|4092,4093
.|4093,4094
50|4094,4096
*|4096,4097
<EOL>|4097,4098
<EOL>|4098,4099
DISCHARGE|4099,4108
LABS|4109,4113
:|4113,4114
<EOL>|4114,4115
_|4115,4116
_|4116,4117
_|4117,4118
07|4119,4121
:|4121,4122
28AM|4122,4126
BLOOD|4127,4132
WBC|4133,4136
-|4136,4137
4.2|4137,4140
RBC|4141,4144
-|4144,4145
3|4145,4146
.|4146,4147
85|4147,4149
*|4149,4150
Hgb|4151,4154
-|4154,4155
12|4155,4157
.|4157,4158
5|4158,4159
*|4159,4160
Hct|4161,4164
-|4164,4165
36|4165,4167
.|4167,4168
0|4168,4169
*|4169,4170
<EOL>|4171,4172
MCV|4172,4175
-|4175,4176
94|4176,4178
MCH|4179,4182
-|4182,4183
32|4183,4185
.|4185,4186
5|4186,4187
*|4187,4188
MCHC|4189,4193
-|4193,4194
34.7|4194,4198
RDW|4199,4202
-|4202,4203
12.9|4203,4207
Plt|4208,4211
_|4212,4213
_|4213,4214
_|4214,4215
<EOL>|4215,4216
_|4216,4217
_|4217,4218
_|4218,4219
07|4220,4222
:|4222,4223
28AM|4223,4227
BLOOD|4228,4233
Glucose|4234,4241
-|4241,4242
104|4242,4245
*|4245,4246
UreaN|4247,4252
-|4252,4253
30|4253,4255
*|4255,4256
Creat|4257,4262
-|4262,4263
1|4263,4264
.|4264,4265
6|4265,4266
*|4266,4267
Na|4268,4270
-|4270,4271
142|4271,4274
<EOL>|4275,4276
K|4276,4277
-|4277,4278
4.3|4278,4281
Cl|4282,4284
-|4284,4285
106|4285,4288
HCO3|4289,4293
-|4293,4294
26|4294,4296
AnGap|4297,4302
-|4302,4303
14|4303,4305
<EOL>|4305,4306
<EOL>|4306,4307
IMAGING|4307,4314
:|4314,4315
<EOL>|4315,4316
_|4316,4317
_|4317,4318
_|4318,4319
CXR|4320,4323
<EOL>|4323,4324
PA|4324,4326
and|4327,4330
lateral|4331,4338
views|4339,4344
of|4345,4347
the|4348,4351
chest|4352,4357
provided|4358,4366
.|4366,4367
The|4368,4371
lungs|4372,4377
are|4378,4381
<EOL>|4382,4383
adequately|4383,4393
<EOL>|4394,4395
aerated|4395,4402
.|4402,4403
There|4404,4409
is|4410,4412
a|4413,4414
focal|4415,4420
consolidation|4421,4434
at|4435,4437
the|4438,4441
left|4442,4446
lung|4447,4451
base|4452,4456
<EOL>|4457,4458
adjacent|4458,4466
to|4467,4469
the|4470,4473
lateral|4474,4481
hemidiaphragm|4482,4495
.|4495,4496
There|4497,4502
is|4503,4505
mild|4506,4510
vascular|4511,4519
<EOL>|4520,4521
engorgement|4521,4532
.|4532,4533
There|4534,4539
is|4540,4542
bilateral|4543,4552
apical|4553,4559
pleural|4560,4567
thickening|4568,4578
.|4578,4579
The|4580,4583
<EOL>|4584,4585
cardiomediastinal|4585,4602
silhouette|4603,4613
is|4614,4616
remarkable|4617,4627
for|4628,4631
aortic|4632,4638
arch|4639,4643
<EOL>|4644,4645
calcifications|4645,4659
.|4659,4660
The|4661,4664
heart|4665,4670
is|4671,4673
top|4674,4677
normal|4678,4684
in|4685,4687
size|4688,4692
.|4692,4693
<EOL>|4694,4695
<EOL>|4695,4696
_|4696,4697
_|4697,4698
_|4698,4699
ECHO|4700,4704
<EOL>|4704,4705
The|4705,4708
left|4709,4713
atrium|4714,4720
is|4721,4723
mildly|4724,4730
dilated|4731,4738
.|4738,4739
Left|4740,4744
ventricular|4745,4756
wall|4757,4761
<EOL>|4762,4763
thicknesses|4763,4774
and|4775,4778
cavity|4779,4785
size|4786,4790
are|4791,4794
normal|4795,4801
.|4801,4802
There|4803,4808
is|4809,4811
mild|4812,4816
regional|4817,4825
<EOL>|4826,4827
left|4827,4831
ventricular|4832,4843
systolic|4844,4852
dysfunction|4853,4864
with|4865,4869
focal|4870,4875
apical|4876,4882
<EOL>|4883,4884
hypokinesis|4884,4895
.|4895,4896
The|4897,4900
remaining|4901,4910
segments|4911,4919
contract|4920,4928
normally|4929,4937
(|4938,4939
LVEF|4939,4943
=|4944,4945
55|4946,4948
<EOL>|4949,4950
%|4950,4951
)|4951,4952
.|4952,4953
No|4954,4956
masses|4957,4963
or|4964,4966
thrombi|4967,4974
are|4975,4978
seen|4979,4983
in|4984,4986
the|4987,4990
left|4991,4995
ventricle|4996,5005
.|5005,5006
Right|5007,5012
<EOL>|5013,5014
ventricular|5014,5025
chamber|5026,5033
size|5034,5038
and|5039,5042
free|5043,5047
wall|5048,5052
motion|5053,5059
are|5060,5063
normal|5064,5070
.|5070,5071
There|5072,5077
<EOL>|5078,5079
are|5079,5082
three|5083,5088
aortic|5089,5095
valve|5096,5101
leaflets|5102,5110
.|5110,5111
There|5112,5117
is|5118,5120
mild|5121,5125
aortic|5126,5132
valve|5133,5138
<EOL>|5139,5140
stenosis|5140,5148
(|5149,5150
valve|5150,5155
area|5156,5160
1.7|5161,5164
cm2|5164,5167
)|5167,5168
.|5168,5169
Mild|5170,5174
(|5175,5176
1|5176,5177
+|5177,5178
)|5178,5179
aortic|5180,5186
regurgitation|5187,5200
is|5201,5203
<EOL>|5204,5205
seen|5205,5209
.|5209,5210
The|5211,5214
mitral|5215,5221
valve|5222,5227
leaflets|5228,5236
are|5237,5240
mildly|5241,5247
thickened|5248,5257
.|5257,5258
Trivial|5259,5266
<EOL>|5267,5268
mitral|5268,5274
regurgitation|5275,5288
is|5289,5291
seen|5292,5296
.|5296,5297
The|5298,5301
pulmonary|5302,5311
artery|5312,5318
systolic|5319,5327
<EOL>|5328,5329
pressure|5329,5337
could|5338,5343
not|5344,5347
be|5348,5350
determined|5351,5361
.|5361,5362
There|5363,5368
is|5369,5371
a|5372,5373
trivial|5374,5381
/|5381,5382
physiologic|5382,5393
<EOL>|5394,5395
pericardial|5395,5406
effusion|5407,5415
.|5415,5416
<EOL>|5417,5418
<EOL>|5418,5419
IMPRESSION|5419,5429
:|5429,5430
Normal|5431,5437
left|5438,5442
ventricular|5443,5454
cavity|5455,5461
size|5462,5466
with|5467,5471
mild|5472,5476
<EOL>|5477,5478
regional|5478,5486
systolic|5487,5495
dysfunction|5496,5507
most|5508,5512
c|5513,5514
/|5514,5515
w|5515,5516
CAD|5517,5520
(|5521,5522
distal|5522,5528
LAD|5529,5532
<EOL>|5533,5534
distribution|5534,5546
)|5546,5547
.|5547,5548
Mild|5549,5553
aortic|5554,5560
valve|5561,5566
stenosis|5567,5575
.|5575,5576
Mild|5577,5581
aortic|5582,5588
<EOL>|5589,5590
regurgitation|5590,5603
.|5603,5604
<EOL>|5605,5606
<EOL>|5607,5608
Mr.|5631,5634
_|5635,5636
_|5636,5637
_|5637,5638
is|5639,5641
an|5642,5644
_|5645,5646
_|5646,5647
_|5647,5648
with|5649,5653
history|5654,5661
of|5662,5664
AAA|5665,5668
s|5669,5670
/|5670,5671
p|5671,5672
repair|5673,5679
<EOL>|5680,5681
complicated|5681,5692
by|5693,5695
MI|5696,5698
,|5698,5699
hypertension|5700,5712
,|5712,5713
and|5714,5717
hyperlipidemia|5718,5732
who|5733,5736
<EOL>|5737,5738
presented|5738,5747
with|5748,5752
nasal|5753,5758
fractures|5759,5768
and|5769,5772
epistaxis|5773,5782
after|5783,5788
mechanical|5789,5799
<EOL>|5800,5801
fall|5801,5805
with|5806,5810
hospital|5811,5819
course|5820,5826
complicated|5827,5838
by|5839,5841
NSTEMI|5842,5848
.|5848,5849
<EOL>|5849,5850
<EOL>|5850,5851
#|5851,5852
Epistaxis|5852,5861
,|5861,5862
nasal|5863,5868
fractures|5869,5878
<EOL>|5878,5879
Patient|5879,5886
presenting|5887,5897
after|5898,5903
mechanical|5904,5914
fall|5915,5919
with|5920,5924
Rhinorockets|5925,5937
<EOL>|5938,5939
placed|5939,5945
at|5946,5948
outside|5949,5956
hospital|5957,5965
for|5966,5969
ongoing|5970,5977
epistaxis|5978,5987
.|5987,5988
CT|5989,5991
scan|5992,5996
from|5997,6001
<EOL>|6002,6003
that|6003,6007
hospital|6008,6016
demonstrated|6017,6029
nasal|6030,6035
bone|6036,6040
and|6041,6044
septal|6045,6051
fractures|6052,6061
.|6061,6062
The|6063,6066
<EOL>|6067,6068
Rhinorockets|6068,6080
were|6081,6085
maintained|6086,6096
while|6097,6102
inpatient|6103,6112
and|6113,6116
discontinued|6117,6129
<EOL>|6130,6131
prior|6131,6136
to|6137,6139
discharge|6140,6149
.|6149,6150
He|6151,6153
was|6154,6157
encouraged|6158,6168
to|6169,6171
use|6172,6175
oxymetolazone|6176,6189
nasal|6190,6195
<EOL>|6196,6197
spray|6197,6202
and|6203,6206
hold|6207,6211
pressure|6212,6220
should|6221,6227
bleeding|6228,6236
reoccur|6237,6244
.|6244,6245
<EOL>|6246,6247
<EOL>|6247,6248
#|6248,6249
NSTEMI|6249,6255
<EOL>|6255,6256
Patient|6256,6263
found|6264,6269
to|6270,6272
have|6273,6277
mild|6278,6282
elevation|6283,6292
of|6293,6295
troponin|6296,6304
in|6305,6307
the|6308,6311
ED|6312,6314
.|6314,6315
This|6316,6320
<EOL>|6321,6322
was|6322,6325
trended|6326,6333
and|6334,6337
eventually|6338,6348
rose|6349,6353
to|6354,6356
1.5|6357,6360
,|6360,6361
though|6362,6368
MB|6369,6371
component|6372,6381
<EOL>|6382,6383
downtrended|6383,6394
during|6395,6401
course|6402,6408
of|6409,6411
admission|6412,6421
.|6421,6422
The|6423,6426
patient|6427,6434
was|6435,6438
without|6439,6446
<EOL>|6447,6448
chest|6448,6453
pain|6454,6458
or|6459,6461
other|6462,6467
cardiac|6468,6475
symptoms|6476,6484
.|6484,6485
Cardiology|6486,6496
was|6497,6500
consulted|6501,6510
<EOL>|6511,6512
who|6512,6515
thought|6516,6523
that|6524,6528
this|6529,6533
was|6534,6537
most|6538,6542
likely|6543,6549
secondary|6550,6559
to|6560,6562
demand|6563,6569
<EOL>|6570,6571
ischemia|6571,6579
(|6580,6581
type|6581,6585
II|6586,6588
MI|6589,6591
)|6591,6592
secondary|6593,6602
to|6603,6605
his|6606,6609
fall|6610,6614
.|6614,6615
An|6616,6618
echocardiogram|6619,6633
<EOL>|6634,6635
demonstrated|6635,6647
aortic|6648,6654
stenosis|6655,6663
and|6664,6667
likely|6668,6674
distal|6675,6681
LAD|6682,6685
disease|6686,6693
based|6694,6699
<EOL>|6700,6701
on|6701,6703
wall|6704,6708
motion|6709,6715
abnormalities|6716,6729
.|6729,6730
The|6731,6734
patient|6735,6742
's|6742,6744
metoprolol|6745,6755
was|6756,6759
<EOL>|6760,6761
uptitrated|6761,6771
,|6771,6772
his|6773,6776
pravastatin|6777,6788
was|6789,6792
converted|6793,6802
to|6803,6805
atorvastatin|6806,6818
,|6818,6819
his|6820,6823
<EOL>|6824,6825
clopidogrel|6825,6836
was|6837,6840
maintained|6841,6851
,|6851,6852
and|6853,6856
he|6857,6859
was|6860,6863
started|6864,6871
on|6872,6874
aspirin|6875,6882
.|6882,6883
<EOL>|6883,6884
<EOL>|6884,6885
#|6885,6886
Hypoxemia|6886,6895
/|6895,6896
L|6896,6897
basilar|6898,6905
consolidation|6906,6919
<EOL>|6919,6920
Patient|6920,6927
reported|6928,6936
to|6937,6939
be|6940,6942
mildly|6943,6949
hypoxic|6950,6957
in|6958,6960
the|6961,6964
ED|6965,6967
,|6967,6968
though|6969,6975
he|6976,6978
<EOL>|6979,6980
maintained|6980,6990
normal|6991,6997
oxygen|6998,7004
saturations|7005,7016
on|7017,7019
room|7020,7024
air|7025,7028
.|7028,7029
He|7030,7032
denied|7033,7039
<EOL>|7040,7041
shortness|7041,7050
of|7051,7053
breath|7054,7060
or|7061,7063
cough|7064,7069
,|7069,7070
fevers|7071,7077
,|7077,7078
or|7079,7081
other|7082,7087
infectious|7088,7098
<EOL>|7099,7100
symptoms|7100,7108
and|7109,7112
had|7113,7116
no|7117,7119
leukocytosis|7120,7132
.|7132,7133
A|7134,7135
CXR|7136,7139
revealed|7140,7148
consolidation|7149,7162
<EOL>|7163,7164
in|7164,7166
left|7167,7171
lung|7172,7176
,|7176,7177
thought|7178,7185
to|7186,7188
be|7189,7191
possibly|7192,7200
related|7201,7208
to|7209,7211
aspirated|7212,7221
blood|7222,7227
.|7227,7228
<EOL>|7229,7230
-|7230,7231
monitor|7231,7238
O2|7239,7241
saturation|7242,7252
,|7252,7253
temperature|7254,7265
,|7265,7266
trend|7267,7272
WBC|7273,7276
.|7276,7277
He|7278,7280
was|7281,7284
convered|7285,7293
<EOL>|7294,7295
with|7295,7299
antibiotics|7300,7311
while|7312,7317
inpatient|7318,7327
as|7328,7330
he|7331,7333
required|7334,7342
prophylaxis|7343,7354
for|7355,7358
<EOL>|7359,7360
the|7360,7363
Rhinorockets|7364,7376
,|7376,7377
but|7378,7381
this|7382,7386
was|7387,7390
discontinued|7391,7403
upon|7404,7408
discharge|7409,7418
.|7418,7419
<EOL>|7419,7420
<EOL>|7420,7421
#|7421,7422
Acute|7422,7427
kidney|7428,7434
injury|7435,7441
<EOL>|7441,7442
Patient|7442,7449
presented|7450,7459
with|7460,7464
creatinine|7465,7475
of|7476,7478
1.5|7479,7482
with|7483,7487
last|7488,7492
creatinine|7493,7503
at|7504,7506
<EOL>|7507,7508
PCP|7508,7511
1.8|7512,7515
.|7515,7516
Patient|7517,7524
was|7525,7528
unaware|7529,7536
of|7537,7539
a|7540,7541
history|7542,7549
of|7550,7552
kidney|7553,7559
disease|7560,7567
.|7567,7568
The|7569,7572
<EOL>|7573,7574
patient|7574,7581
was|7582,7585
discharged|7586,7596
with|7597,7601
a|7602,7603
stable|7604,7610
creatinine|7611,7621
.|7621,7622
<EOL>|7622,7623
<EOL>|7623,7624
#|7624,7625
Peripheral|7625,7635
vascular|7636,7644
disease|7645,7652
<EOL>|7652,7653
Patient|7653,7660
had|7661,7664
a|7665,7666
history|7667,7674
of|7675,7677
AAA|7678,7681
repair|7682,7688
in|7689,7691
_|7692,7693
_|7693,7694
_|7694,7695
without|7696,7703
history|7704,7711
of|7712,7714
<EOL>|7715,7716
MI|7716,7718
per|7719,7722
PCP|7723,7726
.|7726,7727
Patient|7728,7735
denied|7736,7742
history|7743,7750
of|7751,7753
CABG|7754,7758
or|7759,7761
cardiac|7762,7769
/|7769,7770
peripheral|7770,7780
<EOL>|7781,7782
stents|7782,7788
.|7788,7789
A|7790,7791
cardiac|7792,7799
regimen|7800,7807
was|7808,7811
continued|7812,7821
,|7821,7822
as|7823,7825
above|7826,7831
.|7831,7832
<EOL>|7832,7833
<EOL>|7833,7834
TRANSITIONAL|7834,7846
ISSUES|7847,7853
<EOL>|7853,7854
-|7854,7855
Outpatient|7855,7865
stress|7866,7872
echo|7873,7877
for|7878,7881
futher|7882,7888
evaluation|7889,7899
distal|7900,7906
LAD|7907,7910
disease|7911,7918
<EOL>|7919,7920
(|7920,7921
possibly|7921,7929
a|7930,7931
large|7932,7937
myocardial|7938,7948
territory|7949,7958
at|7959,7961
risk|7962,7966
)|7966,7967
.|7967,7968
<EOL>|7969,7970
-|7970,7971
Repeat|7971,7977
echocardiogram|7978,7992
in|7993,7995
_|7996,7997
_|7997,7998
_|7998,7999
years|8000,8005
to|8006,8008
monitor|8009,8016
mild|8017,8021
AS|8022,8024
/|8024,8025
AR|8025,8027
.|8027,8028
<EOL>|8028,8029
-|8029,8030
If|8030,8032
epistaxis|8033,8042
returns|8043,8050
,|8050,8051
can|8052,8055
use|8056,8059
oxymetolazone|8060,8073
nasal|8074,8079
spray|8080,8085
.|8085,8086
<EOL>|8086,8087
-|8087,8088
Repeat|8088,8094
chest|8095,8100
x-ray|8101,8106
in|8107,8109
_|8110,8111
_|8111,8112
_|8112,8113
weeks|8114,8119
to|8120,8122
ensure|8123,8129
resolution|8130,8140
of|8141,8143
the|8144,8147
LLL|8148,8151
<EOL>|8152,8153
infiltrative|8153,8165
process|8166,8173
.|8173,8174
<EOL>|8174,8175
-|8175,8176
Consider|8176,8184
follow|8185,8191
-|8191,8192
up|8192,8194
with|8195,8199
ENT|8200,8203
or|8204,8206
Plastic|8207,8214
Surgery|8215,8222
for|8223,8226
later|8227,8232
<EOL>|8233,8234
evaluation|8234,8244
of|8245,8247
nasal|8248,8253
fractures|8254,8263
.|8263,8264
<EOL>|8264,8265
-|8265,8266
Repeat|8266,8272
CBC|8273,8276
in|8277,8279
one|8280,8283
week|8284,8288
to|8289,8291
ensure|8292,8298
stability|8299,8308
of|8309,8311
HCT|8312,8315
and|8316,8319
<EOL>|8320,8321
platelets|8321,8330
.|8330,8331
<EOL>|8331,8332
-|8332,8333
Consider|8333,8341
conversion|8342,8352
of|8353,8355
metoprolol|8356,8366
tartrate|8367,8375
to|8376,8378
succinate|8379,8388
for|8389,8392
<EOL>|8393,8394
ease|8394,8398
-|8398,8399
of|8399,8401
-|8401,8402
administration|8402,8416
.|8416,8417
<EOL>|8417,8418
<EOL>|8419,8420
Medications|8420,8431
on|8432,8434
Admission|8435,8444
:|8444,8445
<EOL>|8445,8446
The|8446,8449
Preadmission|8450,8462
Medication|8463,8473
list|8474,8478
is|8479,8481
accurate|8482,8490
and|8491,8494
complete|8495,8503
.|8503,8504
<EOL>|8504,8505
1.|8505,8507
Clopidogrel|8508,8519
75|8520,8522
mg|8523,8525
PO|8526,8528
DAILY|8529,8534
<EOL>|8535,8536
2.|8536,8538
Metoprolol|8539,8549
Tartrate|8550,8558
50|8559,8561
mg|8562,8564
PO|8565,8567
TID|8568,8571
<EOL>|8572,8573
3.|8573,8575
Pravastatin|8576,8587
80|8588,8590
mg|8591,8593
PO|8594,8596
QPM|8597,8600
<EOL>|8601,8602
<EOL>|8602,8603
<EOL>|8604,8605
Discharge|8605,8614
Medications|8615,8626
:|8626,8627
<EOL>|8627,8628
1.|8628,8630
Clopidogrel|8631,8642
75|8643,8645
mg|8646,8648
PO|8649,8651
DAILY|8652,8657
<EOL>|8658,8659
2.|8659,8661
Acetaminophen|8662,8675
650|8676,8679
mg|8680,8682
PO|8683,8685
Q8H|8686,8689
:|8689,8690
PRN|8690,8693
pain|8694,8698
<EOL>|8699,8700
Please|8700,8706
avoid|8707,8712
NSAID|8713,8718
medications|8719,8730
like|8731,8735
ibuprofen|8736,8745
given|8746,8751
your|8752,8756
<EOL>|8757,8758
bleeding|8758,8766
.|8766,8767
<EOL>|8768,8769
3.|8769,8771
Aspirin|8772,8779
81|8780,8782
mg|8783,8785
PO|8786,8788
DAILY|8789,8794
Duration|8795,8803
:|8803,8804
30|8805,8807
Days|8808,8812
<EOL>|8813,8814
4.|8814,8816
Metoprolol|8817,8827
Tartrate|8828,8836
75|8837,8839
mg|8840,8842
PO|8843,8845
TID|8846,8849
<EOL>|8850,8851
RX|8851,8853
*|8854,8855
metoprolol|8855,8865
tartrate|8866,8874
25|8875,8877
mg|8878,8880
3|8881,8882
tablet|8883,8889
(|8889,8890
s|8890,8891
)|8891,8892
by|8893,8895
mouth|8896,8901
three|8902,8907
times|8908,8913
<EOL>|8914,8915
daily|8915,8920
Disp|8921,8925
#|8926,8927
*|8927,8928
270|8928,8931
Tablet|8932,8938
Refills|8939,8946
:|8946,8947
*|8947,8948
0|8948,8949
<EOL>|8949,8950
5.|8950,8952
Atorvastatin|8953,8965
40|8966,8968
mg|8969,8971
PO|8972,8974
QPM|8975,8978
<EOL>|8979,8980
RX|8980,8982
*|8983,8984
atorvastatin|8984,8996
40|8997,8999
mg|9000,9002
1|9003,9004
tablet|9005,9011
(|9011,9012
s|9012,9013
)|9013,9014
by|9015,9017
mouth|9018,9023
every|9024,9029
evening|9030,9037
Disp|9038,9042
<EOL>|9043,9044
#|9044,9045
*|9045,9046
30|9046,9048
Tablet|9049,9055
Refills|9056,9063
:|9063,9064
*|9064,9065
0|9065,9066
<EOL>|9066,9067
6.|9067,9069
Oxymetazoline|9070,9083
1|9084,9085
SPRY|9086,9090
NU|9091,9093
BID|9094,9097
:|9097,9098
PRN|9098,9101
nosebleed|9102,9111
<EOL>|9112,9113
This|9113,9117
can|9118,9121
be|9122,9124
purchased|9125,9134
over-the|9135,9143
-|9143,9144
counter|9144,9151
,|9151,9152
the|9153,9156
brand|9157,9162
name|9163,9167
is|9168,9170
_|9171,9172
_|9172,9173
_|9173,9174
.|9174,9175
<EOL>|9176,9177
<EOL>|9177,9178
<EOL>|9178,9179
<EOL>|9180,9181
Discharge|9181,9190
Disposition|9191,9202
:|9202,9203
<EOL>|9203,9204
Home|9204,9208
With|9209,9213
Service|9214,9221
<EOL>|9221,9222
<EOL>|9223,9224
Facility|9224,9232
:|9232,9233
<EOL>|9233,9234
_|9234,9235
_|9235,9236
_|9236,9237
<EOL>|9237,9238
<EOL>|9239,9240
Discharge|9240,9249
Diagnosis|9250,9259
:|9259,9260
<EOL>|9260,9261
Nasal|9261,9266
fracture|9267,9275
<EOL>|9275,9276
Epistaxis|9276,9285
<EOL>|9285,9286
NSTEMI|9286,9292
<EOL>|9292,9293
<EOL>|9293,9294
<EOL>|9295,9296
Mental|9317,9323
Status|9324,9330
:|9330,9331
Clear|9332,9337
and|9338,9341
coherent|9342,9350
.|9350,9351
<EOL>|9351,9352
Level|9352,9357
of|9358,9360
Consciousness|9361,9374
:|9374,9375
Alert|9376,9381
and|9382,9385
interactive|9386,9397
.|9397,9398
<EOL>|9398,9399
Activity|9399,9407
Status|9408,9414
:|9414,9415
Ambulatory|9416,9426
-|9427,9428
Independent|9429,9440
.|9440,9441
<EOL>|9441,9442
<EOL>|9442,9443
<EOL>|9444,9445
Mr.|9469,9472
_|9473,9474
_|9474,9475
_|9475,9476
,|9476,9477
<EOL>|9477,9478
You|9478,9481
were|9482,9486
admitted|9487,9495
after|9496,9501
you|9502,9505
fell|9506,9510
and|9511,9514
broke|9515,9520
your|9521,9525
nose|9526,9530
.|9530,9531
You|9532,9535
had|9536,9539
<EOL>|9540,9541
nose|9541,9545
bleeds|9546,9552
that|9553,9557
were|9558,9562
difficult|9563,9572
to|9573,9575
control|9576,9583
,|9583,9584
thus|9585,9589
plugs|9590,9595
were|9596,9600
<EOL>|9601,9602
placed|9602,9608
in|9609,9611
your|9612,9616
nose|9617,9621
to|9622,9624
stop|9625,9629
the|9630,9633
bleeding|9634,9642
.|9642,9643
During|9644,9650
your|9651,9655
hospital|9656,9664
<EOL>|9665,9666
course|9666,9672
,|9672,9673
you|9674,9677
were|9678,9682
found|9683,9688
to|9689,9691
have|9692,9696
high|9697,9701
troponins|9702,9711
,|9711,9712
a|9713,9714
blood|9715,9720
test|9721,9725
for|9726,9729
<EOL>|9730,9731
the|9731,9734
heart|9735,9740
.|9740,9741
A|9742,9743
ultrasound|9744,9754
of|9755,9757
your|9758,9762
heart|9763,9768
was|9769,9772
performed|9773,9782
.|9782,9783
You|9784,9787
should|9788,9794
<EOL>|9795,9796
follow|9796,9802
-|9802,9803
up|9803,9805
with|9806,9810
your|9811,9815
PCP|9816,9819
to|9820,9822
discuss|9823,9830
stress|9831,9837
test|9838,9842
.|9842,9843
<EOL>|9843,9844
<EOL>|9844,9845
It|9845,9847
was|9848,9851
a|9852,9853
pleasure|9854,9862
participating|9863,9876
in|9877,9879
your|9880,9884
care|9885,9889
,|9889,9890
thank|9891,9896
you|9897,9900
for|9901,9904
<EOL>|9905,9906
choosing|9906,9914
_|9915,9916
_|9916,9917
_|9917,9918
.|9918,9919
<EOL>|9919,9920
<EOL>|9921,9922
Followup|9922,9930
Instructions|9931,9943
:|9943,9944
<EOL>|9944,9945
_|9945,9946
_|9946,9947
_|9947,9948
<EOL>|9948,9949

