 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|39,48|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|73,82|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|160,169|false|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|160,169|false|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|160,169|false|false|false|C0020517|Hypersensitivity|Allergies
Attribute|Clinical Attribute|SIMPLE_SEGMENT|181,190|true|false|false|C1717415||Allergies
Event|Event|SIMPLE_SEGMENT|181,190|true|false|false|||Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|181,190|true|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|SIMPLE_SEGMENT|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|201,205|true|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|SIMPLE_SEGMENT|201,205|true|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|SIMPLE_SEGMENT|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|SIMPLE_SEGMENT|206,215|true|false|false|||Reactions
Event|Event|SIMPLE_SEGMENT|218,227|false|false|false|||Attending
Finding|Functional Concept|SIMPLE_SEGMENT|218,227|false|false|false|C1999232|Attending (action)|Attending
Finding|Finding|SIMPLE_SEGMENT|236,251|false|false|false|C0277786|Chief complaint (finding)|Chief Complaint
Attribute|Clinical Attribute|SIMPLE_SEGMENT|242,251|false|false|false|C3864418||Complaint
Event|Event|SIMPLE_SEGMENT|242,251|false|false|false|||Complaint
Finding|Finding|SIMPLE_SEGMENT|242,251|false|false|false|C5441521|Complaint (finding)|Complaint
Anatomy|Body Location or Region|SIMPLE_SEGMENT|253,256|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|253,256|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|253,256|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|253,256|false|false|false|||DVT
Finding|Classification|SIMPLE_SEGMENT|259,264|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|SIMPLE_SEGMENT|265,273|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|265,273|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|277,295|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|SIMPLE_SEGMENT|286,295|false|false|false|C0945766||Procedure
Event|Event|SIMPLE_SEGMENT|286,295|false|false|false|||Procedure
Event|Occupational Activity|SIMPLE_SEGMENT|286,295|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|SIMPLE_SEGMENT|286,295|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|286,295|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|SIMPLE_SEGMENT|297,300|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|297,300|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|304,311|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|304,311|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|304,311|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|304,311|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|304,314|false|false|false|C0262926|Medical History|History of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|304,330|false|false|false|C0488508||History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|304,330|false|false|false|C0262512|History of present illness (finding)|History of Present Illness
Finding|Finding|SIMPLE_SEGMENT|315,322|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Idea or Concept|SIMPLE_SEGMENT|315,322|false|false|false|C0150312;C0449450|Present;Presentation|Present
Finding|Finding|SIMPLE_SEGMENT|315,330|false|false|false|C4264312|Present illness|Present Illness
Finding|Sign or Symptom|SIMPLE_SEGMENT|323,330|false|false|false|C0221423|Illness (finding)|Illness
Event|Event|SIMPLE_SEGMENT|367,378|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|367,378|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|383,386|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|383,386|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|383,386|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|383,386|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|383,386|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|388,391|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|388,391|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|393,396|false|false|false|||HLD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|405,408|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|409,414|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|409,417|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|419,422|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|SIMPLE_SEGMENT|419,422|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|419,422|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|SIMPLE_SEGMENT|436,440|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|453,460|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|462,468|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|462,468|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|471,479|false|false|false|||presents
Anatomy|Body Location or Region|SIMPLE_SEGMENT|485,490|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|485,490|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|485,499|false|false|false|C0230443|Structure of left lower leg|lower Left leg
Finding|Functional Concept|SIMPLE_SEGMENT|491,495|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|491,499|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|Left leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|491,508|false|false|false|C2219779|numbness of left leg|Left leg numbness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|496,499|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|496,508|false|true|false|C0857160|Numbness in leg|leg numbness
Event|Event|SIMPLE_SEGMENT|500,508|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|500,508|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|500,508|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|513,517|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|513,517|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|513,517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|513,517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|535,542|false|false|false|||evening
Event|Event|SIMPLE_SEGMENT|548,556|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|548,556|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|548,556|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|557,564|false|false|false|||started
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|579,582|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|SIMPLE_SEGMENT|579,582|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|589,594|false|false|false|||onset
Event|Event|SIMPLE_SEGMENT|599,606|false|false|false|||gradual
Event|Event|SIMPLE_SEGMENT|619,629|false|false|false|||associated
Attribute|Clinical Attribute|SIMPLE_SEGMENT|635,639|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|635,639|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|635,639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|635,639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|640,648|false|false|false|C0026821|Muscle Cramp|cramping
Anatomy|Body Location or Region|SIMPLE_SEGMENT|667,671|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|667,671|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Event|Event|SIMPLE_SEGMENT|673,682|false|false|false|||radiating
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|697,701|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|697,701|false|false|false|C0555980|Foot problem|foot
Finding|Finding|SIMPLE_SEGMENT|737,744|false|false|false|C3888388|Usually|usually
Event|Event|SIMPLE_SEGMENT|761,766|true|false|false|||lying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|770,773|true|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|770,773|true|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|770,773|true|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|785,793|true|false|false|||exertion
Finding|Organism Function|SIMPLE_SEGMENT|785,793|true|false|false|C0015264|Exertion|exertion
Event|Event|SIMPLE_SEGMENT|799,805|false|false|false|||denies
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|806,809|true|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Finding|SIMPLE_SEGMENT|806,818|true|false|false|C0427068;C1836296|Monoparesis of lower limb;Muscle Weakness Lower Limb|leg weakness
Event|Event|SIMPLE_SEGMENT|810,818|true|false|false|||weakness
Finding|Sign or Symptom|SIMPLE_SEGMENT|810,818|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|SIMPLE_SEGMENT|827,831|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|827,831|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|827,831|true|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|SIMPLE_SEGMENT|840,844|true|false|false|||able
Finding|Finding|SIMPLE_SEGMENT|840,844|true|false|false|C1299581|Able (qualifier value)|able
Event|Event|SIMPLE_SEGMENT|849,853|true|false|false|||walk
Event|Event|SIMPLE_SEGMENT|862,872|true|false|false|||assistance
Finding|Social Behavior|SIMPLE_SEGMENT|862,872|true|false|false|C0018896|Helping Behavior|assistance
Attribute|Clinical Attribute|SIMPLE_SEGMENT|884,888|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|884,888|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|884,888|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|884,888|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|893,901|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|893,901|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|893,901|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|906,914|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|925,933|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|925,933|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|925,933|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Location or Region|SIMPLE_SEGMENT|949,953|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|949,953|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Event|Event|SIMPLE_SEGMENT|955,961|false|false|false|||Denies
Anatomy|Body Location or Region|SIMPLE_SEGMENT|965,968|true|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|965,968|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|965,968|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|965,968|true|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|971,977|false|false|false|||Denies
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|978,983|true|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|SIMPLE_SEGMENT|978,983|true|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|SIMPLE_SEGMENT|978,983|true|false|false|C0150920|Spine Problem|spine
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|991,997|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Event|Event|SIMPLE_SEGMENT|991,997|true|false|false|||trauma
Procedure|Health Care Activity|SIMPLE_SEGMENT|991,997|true|false|false|C0548346|Trauma assessment and care|trauma
Finding|Sign or Symptom|SIMPLE_SEGMENT|1002,1011|true|false|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1007,1011|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1007,1011|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1007,1011|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1007,1011|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1016,1028|true|false|false|C0021167|Incontinence|incontinence
Event|Event|SIMPLE_SEGMENT|1016,1028|true|false|false|||incontinence
Event|Event|SIMPLE_SEGMENT|1034,1040|true|false|false|||fevers
Finding|Sign or Symptom|SIMPLE_SEGMENT|1034,1040|true|false|false|C0015967|Fever|fevers
Event|Event|SIMPLE_SEGMENT|1041,1047|true|false|false|||chills
Finding|Sign or Symptom|SIMPLE_SEGMENT|1041,1047|true|false|false|C0085593|Chills|chills
Event|Event|SIMPLE_SEGMENT|1052,1060|true|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|1052,1060|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|1052,1060|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Event|Event|SIMPLE_SEGMENT|1090,1096|false|false|false|||denies
Event|Event|SIMPLE_SEGMENT|1098,1106|true|false|false|||headache
Finding|Sign or Symptom|SIMPLE_SEGMENT|1098,1106|true|false|false|C0018681|Headache|headache
Finding|Functional Concept|SIMPLE_SEGMENT|1108,1114|true|false|false|C0234621|Visual|visual
Finding|Finding|SIMPLE_SEGMENT|1108,1122|true|false|false|C0750280|Visual changes|visual changes
Event|Event|SIMPLE_SEGMENT|1115,1122|true|false|false|||changes
Finding|Functional Concept|SIMPLE_SEGMENT|1115,1122|true|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1124,1129|true|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1124,1129|true|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1124,1134|true|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1124,1134|true|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1130,1134|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1130,1134|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1130,1134|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1130,1134|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1130,1141|false|false|false|C0008031|Chest Pain|pain, chest
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1136,1141|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1136,1141|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|SIMPLE_SEGMENT|1136,1150|false|false|false|C0438716|Chest pressure|chest pressure
Event|Event|SIMPLE_SEGMENT|1142,1150|false|false|false|||pressure
Finding|Finding|SIMPLE_SEGMENT|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|SIMPLE_SEGMENT|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|1142,1150|false|false|false|C0033095||pressure
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1152,1157|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|1152,1157|false|false|false|C0741025|Chest problem|chest
Event|Event|SIMPLE_SEGMENT|1159,1171|false|false|false|||palpitations
Finding|Finding|SIMPLE_SEGMENT|1159,1171|false|false|false|C0030252|Palpitations|palpitations
Event|Event|SIMPLE_SEGMENT|1173,1182|false|false|false|||shortness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1173,1192|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|SIMPLE_SEGMENT|1173,1192|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|SIMPLE_SEGMENT|1186,1192|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1193,1202|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|SIMPLE_SEGMENT|1193,1207|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1203,1207|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|1203,1207|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|1203,1207|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|1203,1207|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|1209,1216|false|false|false|||dysuria
Finding|Sign or Symptom|SIMPLE_SEGMENT|1209,1216|false|false|false|C0013428|Dysuria|dysuria
Event|Event|SIMPLE_SEGMENT|1222,1230|false|false|false|||diarrhea
Finding|Finding|SIMPLE_SEGMENT|1222,1230|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|SIMPLE_SEGMENT|1222,1230|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Finding|SIMPLE_SEGMENT|1235,1255|false|false|false|C0262926;C0455458|Medical History;PMH - past medical history|Past Medical History
Event|Event|SIMPLE_SEGMENT|1240,1247|false|false|false|||Medical
Finding|Functional Concept|SIMPLE_SEGMENT|1240,1247|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|SIMPLE_SEGMENT|1240,1247|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|SIMPLE_SEGMENT|1240,1247|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1240,1247|false|false|false|C0199168|Medical service|Medical
Finding|Finding|SIMPLE_SEGMENT|1240,1255|false|false|false|C0262926|Medical History|Medical History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1248,1255|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1259,1271|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|1259,1271|false|false|false|||hypertension
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1276,1284|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Event|Event|SIMPLE_SEGMENT|1276,1284|false|false|false|||diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1292,1295|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1292,1295|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Event|Event|SIMPLE_SEGMENT|1292,1295|false|false|false|||CVA
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1297,1307|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1308,1317|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1318,1324|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|SIMPLE_SEGMENT|1318,1324|false|false|false|||stroke
Finding|Finding|SIMPLE_SEGMENT|1318,1324|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1336,1339|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1336,1339|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1336,1339|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1336,1339|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1336,1339|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1357,1360|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|1357,1360|false|false|false|||BMS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1392,1419|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1403,1411|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1403,1419|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1412,1419|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|1412,1419|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1421,1433|false|true|false|C0021775|Intermittent Claudication|claudication
Event|Event|SIMPLE_SEGMENT|1421,1433|false|false|false|||claudication
Finding|Finding|SIMPLE_SEGMENT|1421,1433|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1448,1456|false|false|false|C0005847|Blood Vessel|vascular
Event|Event|SIMPLE_SEGMENT|1458,1465|false|false|false|||managed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|1483,1488|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|1483,1491|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1492,1495|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|1492,1495|false|false|false|||CKD
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|1497,1505|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|1497,1505|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|1497,1505|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1519,1523|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Event|Event|SIMPLE_SEGMENT|1519,1523|false|false|false|||GERD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1524,1534|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1524,1540|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Event|SIMPLE_SEGMENT|1535,1540|false|false|false|||rings
Finding|Functional Concept|SIMPLE_SEGMENT|1543,1549|false|false|false|C0728831|Social|Social
Finding|Finding|SIMPLE_SEGMENT|1543,1557|false|false|false|C0424945;C3714536|Social History;Social and personal history|Social History
Event|Event|SIMPLE_SEGMENT|1550,1557|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1550,1557|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1550,1557|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1550,1557|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Classification|SIMPLE_SEGMENT|1563,1569|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Conceptual Entity|SIMPLE_SEGMENT|1563,1569|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Idea or Concept|SIMPLE_SEGMENT|1563,1569|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Intellectual Product|SIMPLE_SEGMENT|1563,1569|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|Family
Finding|Finding|SIMPLE_SEGMENT|1563,1577|false|false|false|C0241889|Family Medical History|Family History
Event|Event|SIMPLE_SEGMENT|1570,1577|false|false|false|||History
Finding|Conceptual Entity|SIMPLE_SEGMENT|1570,1577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|SIMPLE_SEGMENT|1570,1577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|SIMPLE_SEGMENT|1570,1577|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Activity|SIMPLE_SEGMENT|1594,1598|false|false|false|C1947906|Sorting|sort
Event|Event|SIMPLE_SEGMENT|1594,1598|false|false|false|||sort
Finding|Cell Function|SIMPLE_SEGMENT|1594,1598|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|SIMPLE_SEGMENT|1594,1598|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1602,1608|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1602,1608|false|false|false|||cancer
Finding|Conceptual Entity|SIMPLE_SEGMENT|1610,1616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|SIMPLE_SEGMENT|1610,1616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Event|Event|SIMPLE_SEGMENT|1617,1621|false|false|false|||died
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1641,1645|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1641,1645|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1641,1645|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|SIMPLE_SEGMENT|1641,1645|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1641,1653|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1646,1653|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|1646,1653|false|false|false|||disease
Finding|Idea or Concept|SIMPLE_SEGMENT|1656,1662|false|false|false|C1546508|Relationship - Mother|Mother
Event|Event|SIMPLE_SEGMENT|1663,1667|false|false|false|||died
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|SIMPLE_SEGMENT|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Event|Event|SIMPLE_SEGMENT|1689,1696|false|false|false|||unknown
Finding|Finding|SIMPLE_SEGMENT|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|SIMPLE_SEGMENT|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|SIMPLE_SEGMENT|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|SIMPLE_SEGMENT|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Event|Event|SIMPLE_SEGMENT|1697,1702|false|false|false|||cause
Finding|Conceptual Entity|SIMPLE_SEGMENT|1697,1702|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|SIMPLE_SEGMENT|1697,1702|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1715,1718|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|1715,1718|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|1715,1718|true|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|1715,1718|true|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|1715,1718|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|SIMPLE_SEGMENT|1722,1742|true|false|false|C0085298|Sudden Cardiac Death|sudden cardiac death
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1729,1736|true|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|SIMPLE_SEGMENT|1729,1736|true|false|false|C1314974|Cardiac attachment|cardiac
Finding|Pathologic Function|SIMPLE_SEGMENT|1729,1742|true|false|false|C0376297|Cardiac Death|cardiac death
Event|Event|SIMPLE_SEGMENT|1737,1742|true|false|false|||death
Finding|Finding|SIMPLE_SEGMENT|1737,1742|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|SIMPLE_SEGMENT|1737,1742|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|SIMPLE_SEGMENT|1737,1742|true|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Event|Event|SIMPLE_SEGMENT|1759,1766|true|false|false|||history
Finding|Conceptual Entity|SIMPLE_SEGMENT|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|SIMPLE_SEGMENT|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|SIMPLE_SEGMENT|1759,1769|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1771,1777|true|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|SIMPLE_SEGMENT|1771,1777|true|false|false|||cancer
Event|Event|SIMPLE_SEGMENT|1781,1789|false|false|false|||Physical
Finding|Finding|SIMPLE_SEGMENT|1781,1789|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Finding|Functional Concept|SIMPLE_SEGMENT|1781,1789|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|Physical
Procedure|Health Care Activity|SIMPLE_SEGMENT|1781,1789|false|false|false|C0031809|Physical Examination|Physical
Finding|Finding|SIMPLE_SEGMENT|1781,1794|false|false|false|C1509143|physical examination (physical finding)|Physical Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1781,1794|false|false|false|C0031809|Physical Examination|Physical Exam
Event|Event|SIMPLE_SEGMENT|1790,1794|false|false|false|||Exam
Finding|Functional Concept|SIMPLE_SEGMENT|1790,1794|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1790,1794|false|false|false|C0582103|Medical Examination|Exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|1796,1805|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|1806,1814|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|1806,1814|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|1806,1819|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1806,1819|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|1815,1819|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|1815,1819|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|1815,1819|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|SIMPLE_SEGMENT|1866,1873|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|1866,1873|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|1866,1873|false|false|false|C3812897|General medical service|General
Finding|Mental Process|SIMPLE_SEGMENT|1875,1883|false|false|false|C2987187|Pleasant|Pleasant
Event|Event|SIMPLE_SEGMENT|1884,1890|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|1884,1890|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|1884,1890|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|1892,1898|false|false|false|||laying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1902,1905|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|1902,1905|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|1902,1905|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|1907,1914|false|false|false|||resting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1931,1934|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1931,1934|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|1931,1934|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|1931,1934|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1938,1943|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1945,1951|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|1945,1951|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|1945,1951|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|1945,1951|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|1952,1961|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|1952,1961|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|1963,1966|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|1963,1966|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|1968,1978|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|1979,1984|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|1979,1984|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|1986,1990|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|1992,1997|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|1992,1997|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2000,2004|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2000,2004|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|2000,2004|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|2006,2012|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|2006,2012|true|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|2014,2017|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2014,2017|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|2022,2030|true|false|false|||elevated
Event|Activity|SIMPLE_SEGMENT|2046,2050|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|2046,2050|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|2046,2050|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|2055,2061|true|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2055,2061|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2055,2061|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|2082,2089|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2082,2089|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2091,2095|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2091,2095|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2098,2105|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2108,2113|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|2133,2141|false|false|false|||crackles
Finding|Finding|SIMPLE_SEGMENT|2133,2141|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Event|Event|SIMPLE_SEGMENT|2142,2150|false|false|false|||improved
Drug|Organic Chemical|SIMPLE_SEGMENT|2156,2161|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2156,2161|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|SIMPLE_SEGMENT|2156,2161|false|false|false|||cough
Finding|Sign or Symptom|SIMPLE_SEGMENT|2156,2161|false|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2165,2172|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2165,2172|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|2165,2172|false|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|2165,2172|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2174,2179|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2174,2179|false|false|false|||obese
Finding|Finding|SIMPLE_SEGMENT|2174,2187|false|false|false|C0426650|Obese abdomen|obese abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2180,2187|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2180,2187|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|2180,2187|false|false|false|C0941288|Abdomen problem|abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2189,2193|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2189,2193|true|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2226,2233|true|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|2237,2245|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|2237,2245|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2249,2252|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|2249,2252|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|2249,2252|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|2254,2258|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|2254,2258|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|2254,2258|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|2260,2264|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|2265,2273|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|2278,2284|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|2278,2284|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|2278,2284|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|2278,2284|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|SIMPLE_SEGMENT|2286,2291|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2286,2296|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2292,2296|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2292,2296|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|SIMPLE_SEGMENT|2292,2305|false|false|false|C0238882|Swollen calf|calf swelling
Event|Event|SIMPLE_SEGMENT|2297,2305|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|2297,2305|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|2297,2305|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|SIMPLE_SEGMENT|2320,2324|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2320,2329|false|false|false|C0489800|Posterior part of left leg|left calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2325,2329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2325,2329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|SIMPLE_SEGMENT|2325,2338|false|false|false|C0238882|Swollen calf|calf swelling
Event|Event|SIMPLE_SEGMENT|2330,2338|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|2330,2338|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|2330,2338|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2343,2347|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2343,2347|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|SIMPLE_SEGMENT|2343,2358|true|false|false|C0238883|CALF TENDERNESS|calf tenderness
Event|Event|SIMPLE_SEGMENT|2348,2358|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|2348,2358|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|2348,2358|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|2362,2371|true|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2362,2371|true|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2380,2388|false|false|false|C0222007|Structure of nail of toe|toenails
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2390,2398|false|false|false|C0043345|Xeroderma|dry skin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2390,2398|false|false|false|C0720057|Dry Skin brand of emollient|dry skin
Finding|Sign or Symptom|SIMPLE_SEGMENT|2390,2398|false|false|false|C0151908|Dry skin|dry skin
Anatomy|Body System|SIMPLE_SEGMENT|2394,2398|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|2394,2398|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2405,2409|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2411,2417|false|false|false|C0018534|Hallux structure|Hallux
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|2418,2424|false|false|false|C0042282|Valgus deformity|valgus
Event|Event|SIMPLE_SEGMENT|2418,2424|false|false|false|||valgus
Event|Event|SIMPLE_SEGMENT|2444,2450|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|2444,2450|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|SIMPLE_SEGMENT|2456,2464|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|2456,2464|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2471,2476|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|2471,2476|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2471,2488|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2477,2488|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|2506,2515|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|2506,2515|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|2506,2515|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|2506,2515|false|false|false|C2229507|sensory exam|sensation
Finding|Body Substance|SIMPLE_SEGMENT|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|2519,2528|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|2529,2537|false|false|false|||PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2529,2537|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|SIMPLE_SEGMENT|2529,2537|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|SIMPLE_SEGMENT|2529,2537|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|SIMPLE_SEGMENT|2529,2542|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2529,2542|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|SIMPLE_SEGMENT|2538,2542|false|false|false|||EXAM
Finding|Functional Concept|SIMPLE_SEGMENT|2538,2542|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|SIMPLE_SEGMENT|2538,2542|false|false|false|C0582103|Medical Examination|EXAM
Attribute|Clinical Attribute|SIMPLE_SEGMENT|2593,2597|false|false|false|C2317096|Saturation of Peripheral Oxygen|SpO2
Event|Event|SIMPLE_SEGMENT|2620,2627|false|false|false|||General
Finding|Classification|SIMPLE_SEGMENT|2620,2627|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|SIMPLE_SEGMENT|2620,2627|false|false|false|C3812897|General medical service|General
Finding|Mental Process|SIMPLE_SEGMENT|2629,2637|false|false|false|C2987187|Pleasant|Pleasant
Event|Event|SIMPLE_SEGMENT|2638,2644|false|false|false|||affect
Finding|Mental Process|SIMPLE_SEGMENT|2638,2644|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|SIMPLE_SEGMENT|2638,2644|false|false|false|C2237113|assessment of affect|affect
Event|Event|SIMPLE_SEGMENT|2646,2652|false|false|false|||laying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2656,2659|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|SIMPLE_SEGMENT|2656,2659|false|false|false|||bed
Finding|Intellectual Product|SIMPLE_SEGMENT|2656,2659|false|false|false|C2346952|Bachelor of Education|bed
Event|Event|SIMPLE_SEGMENT|2661,2668|false|false|false|||resting
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2685,2688|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2685,2688|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|SIMPLE_SEGMENT|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|SIMPLE_SEGMENT|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|SIMPLE_SEGMENT|2685,2688|false|false|false|||NAD
Finding|Finding|SIMPLE_SEGMENT|2685,2688|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2692,2697|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2699,2705|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2699,2705|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|SIMPLE_SEGMENT|2699,2705|false|false|false|||Sclera
Procedure|Health Care Activity|SIMPLE_SEGMENT|2699,2705|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|SIMPLE_SEGMENT|2706,2715|false|false|false|||anicteric
Finding|Finding|SIMPLE_SEGMENT|2706,2715|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2717,2720|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2717,2720|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2722,2732|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|SIMPLE_SEGMENT|2733,2738|false|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2733,2738|false|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|2740,2744|false|false|false|||EOMI
Event|Event|SIMPLE_SEGMENT|2746,2751|false|false|false|||PERRL
Finding|Finding|SIMPLE_SEGMENT|2746,2751|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2754,2758|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|SIMPLE_SEGMENT|2754,2758|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|SIMPLE_SEGMENT|2754,2758|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|SIMPLE_SEGMENT|2760,2766|true|false|false|||Supple
Finding|Functional Concept|SIMPLE_SEGMENT|2760,2766|true|false|false|C0332254|Supple|Supple
Event|Event|SIMPLE_SEGMENT|2768,2771|true|false|false|||JVP
Finding|Finding|SIMPLE_SEGMENT|2768,2771|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|SIMPLE_SEGMENT|2776,2784|true|false|false|||elevated
Event|Activity|SIMPLE_SEGMENT|2800,2804|false|false|false|C0871208|Rating (action)|rate
Event|Event|SIMPLE_SEGMENT|2800,2804|false|false|false|||rate
Finding|Idea or Concept|SIMPLE_SEGMENT|2800,2804|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|SIMPLE_SEGMENT|2809,2815|true|false|false|||rhythm
Finding|Finding|SIMPLE_SEGMENT|2809,2815|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|SIMPLE_SEGMENT|2809,2815|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|SIMPLE_SEGMENT|2836,2843|true|false|false|||murmurs
Finding|Finding|SIMPLE_SEGMENT|2836,2843|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|SIMPLE_SEGMENT|2845,2849|true|false|false|||rubs
Finding|Finding|SIMPLE_SEGMENT|2845,2849|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|SIMPLE_SEGMENT|2852,2859|true|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|2862,2867|false|false|false|C0024109|Lung|Lungs
Event|Event|SIMPLE_SEGMENT|2869,2874|true|false|false|||clear
Finding|Idea or Concept|SIMPLE_SEGMENT|2869,2874|true|false|false|C1550016|Remote control command - Clear|clear
Event|Event|SIMPLE_SEGMENT|2878,2890|true|false|false|||auscultation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|2878,2890|true|false|false|C0004339|Auscultation|auscultation
Event|Event|SIMPLE_SEGMENT|2913,2920|true|false|false|||wheezes
Finding|Sign or Symptom|SIMPLE_SEGMENT|2913,2920|true|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2932,2939|true|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2932,2939|true|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|SIMPLE_SEGMENT|2932,2939|true|false|false|||Abdomen
Finding|Finding|SIMPLE_SEGMENT|2932,2939|true|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2941,2946|false|false|false|C0028754|Obesity|obese
Event|Event|SIMPLE_SEGMENT|2941,2946|false|false|false|||obese
Finding|Finding|SIMPLE_SEGMENT|2941,2954|false|false|false|C0426650|Obese abdomen|obese abdomen
Anatomy|Body Location or Region|SIMPLE_SEGMENT|2947,2954|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|SIMPLE_SEGMENT|2947,2954|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|SIMPLE_SEGMENT|2947,2954|false|false|false|C0941288|Abdomen problem|abdomen
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|2956,2960|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|SIMPLE_SEGMENT|2956,2960|true|false|false|||soft
Event|Event|SIMPLE_SEGMENT|2993,3000|true|false|false|||rebound
Event|Event|SIMPLE_SEGMENT|3004,3012|true|false|false|||guarding
Finding|Finding|SIMPLE_SEGMENT|3004,3012|true|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|SIMPLE_SEGMENT|3016,3019|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|SIMPLE_SEGMENT|3016,3019|false|false|false|||Ext
Finding|Gene or Genome|SIMPLE_SEGMENT|3016,3019|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|SIMPLE_SEGMENT|3021,3025|false|false|false|||Warm
Finding|Finding|SIMPLE_SEGMENT|3021,3025|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|3021,3025|false|false|false|C0687712|warming process|Warm
Finding|Finding|SIMPLE_SEGMENT|3027,3031|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|3032,3040|false|false|false|||perfused
Drug|Food|SIMPLE_SEGMENT|3054,3060|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|3054,3060|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|3054,3060|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|3054,3060|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3090,3095|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|3090,3095|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|3090,3095|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3090,3095|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3090,3095|false|false|false|C0034107|Pulse taking|pulse
Event|Event|SIMPLE_SEGMENT|3099,3102|false|false|false|||LLE
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3119,3124|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|3119,3124|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|3119,3124|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3119,3124|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3119,3124|false|false|false|C0034107|Pulse taking|pulse
Event|Event|SIMPLE_SEGMENT|3128,3131|false|false|false|||LLE
Finding|Conceptual Entity|SIMPLE_SEGMENT|3136,3142|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3136,3148|false|false|false|C0232142||radial pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3136,3148|false|false|false|C2363059|examination of radial pulses|radial pulse
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3143,3148|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|3143,3148|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|3143,3148|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3143,3148|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3143,3148|false|false|false|C0034107|Pulse taking|pulse
Finding|Finding|SIMPLE_SEGMENT|3143,3151|false|false|false|C5238854|Pulse Wave Normal|pulse 2+
Finding|Conceptual Entity|SIMPLE_SEGMENT|3155,3161|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3155,3167|false|false|false|C0232142||radial pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3155,3167|false|false|false|C2363059|examination of radial pulses|radial pulse
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3162,3167|false|false|false|C0232117|Pulse Rate|pulse
Event|Event|SIMPLE_SEGMENT|3162,3167|false|false|false|||pulse
Finding|Physiologic Function|SIMPLE_SEGMENT|3162,3167|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|3162,3167|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|SIMPLE_SEGMENT|3162,3167|false|false|false|C0034107|Pulse taking|pulse
Finding|Finding|SIMPLE_SEGMENT|3162,3170|false|false|false|C5238852|Pulse Wave Decreased|pulse 1+
Finding|Intellectual Product|SIMPLE_SEGMENT|3172,3176|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|SIMPLE_SEGMENT|3177,3182|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3177,3187|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3183,3187|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3183,3187|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|SIMPLE_SEGMENT|3183,3196|false|false|false|C0238882|Swollen calf|calf swelling
Event|Event|SIMPLE_SEGMENT|3188,3196|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|3188,3196|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|3188,3196|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|SIMPLE_SEGMENT|3211,3215|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3211,3220|false|false|false|C0489800|Posterior part of left leg|left calf
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3216,3220|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3216,3220|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|SIMPLE_SEGMENT|3216,3229|false|false|false|C0238882|Swollen calf|calf swelling
Event|Event|SIMPLE_SEGMENT|3221,3229|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|3221,3229|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|3221,3229|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3234,3238|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3234,3238|true|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|SIMPLE_SEGMENT|3234,3249|true|false|false|C0238883|CALF TENDERNESS|calf tenderness
Event|Event|SIMPLE_SEGMENT|3239,3249|true|false|false|||tenderness
Finding|Mental Process|SIMPLE_SEGMENT|3239,3249|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|SIMPLE_SEGMENT|3239,3249|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|SIMPLE_SEGMENT|3254,3263|true|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3254,3263|true|false|false|C0030247|Palpation|palpation
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3268,3272|true|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|3268,3272|true|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|3268,3272|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|3268,3272|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|3276,3285|true|false|false|||palpation
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|3276,3285|true|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|SIMPLE_SEGMENT|3289,3293|true|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3313,3317|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|3313,3317|false|false|false|C0555980|Foot problem|foot
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|3321,3328|false|false|false|C0376154|Skin callus|callous
Event|Event|SIMPLE_SEGMENT|3321,3328|false|false|false|||callous
Event|Event|SIMPLE_SEGMENT|3329,3336|false|false|false|||present
Finding|Finding|SIMPLE_SEGMENT|3329,3336|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|SIMPLE_SEGMENT|3329,3336|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|SIMPLE_SEGMENT|3340,3344|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3353,3357|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|SIMPLE_SEGMENT|3353,3357|false|false|false|C0555980|Foot problem|foot
Finding|Finding|SIMPLE_SEGMENT|3359,3373|false|false|false|C4540337|Thick toenails|Thick toenails
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3365,3373|false|false|false|C0222007|Structure of nail of toe|toenails
Event|Event|SIMPLE_SEGMENT|3365,3373|false|false|false|||toenails
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3375,3383|false|false|false|C0043345|Xeroderma|dry skin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3375,3383|false|false|false|C0720057|Dry Skin brand of emollient|dry skin
Finding|Sign or Symptom|SIMPLE_SEGMENT|3375,3383|false|false|false|C0151908|Dry skin|dry skin
Anatomy|Body System|SIMPLE_SEGMENT|3379,3383|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3379,3383|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|3379,3383|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Event|Event|SIMPLE_SEGMENT|3379,3383|false|false|false|||skin
Finding|Body Substance|SIMPLE_SEGMENT|3379,3383|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|SIMPLE_SEGMENT|3379,3383|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3391,3395|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Finding|Functional Concept|SIMPLE_SEGMENT|3408,3417|false|false|false|C0702114|indurated|indurated
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3418,3422|false|false|false|C1550235|Cord - Body Parts|cord
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3418,3422|false|false|false|C3489532|Cone-Rod Dystrophy 2|cord
Finding|Functional Concept|SIMPLE_SEGMENT|3426,3430|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3426,3448|false|false|false|C0694648|left antecubital fossa|left antecubital fossa
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3431,3442|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3431,3448|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|3443,3448|false|false|false|C0836913|Fossa|fossa
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3457,3462|false|false|false|C5890168||alert
Drug|Organic Chemical|SIMPLE_SEGMENT|3457,3462|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3457,3462|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|SIMPLE_SEGMENT|3457,3462|false|false|false|||alert
Finding|Finding|SIMPLE_SEGMENT|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|SIMPLE_SEGMENT|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|SIMPLE_SEGMENT|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|SIMPLE_SEGMENT|3467,3475|false|false|false|||oriented
Finding|Finding|SIMPLE_SEGMENT|3467,3475|false|false|false|C1961028|Oriented to place|oriented
Event|Event|SIMPLE_SEGMENT|3490,3496|false|false|false|||intact
Finding|Finding|SIMPLE_SEGMENT|3490,3496|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Organic Chemical|SIMPLE_SEGMENT|3502,3505|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3502,3505|false|false|false|C0939812|Ruta graveolens preparation|RUE
Event|Event|SIMPLE_SEGMENT|3502,3505|false|false|false|||RUE
Finding|Idea or Concept|SIMPLE_SEGMENT|3512,3520|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|SIMPLE_SEGMENT|3521,3524|false|false|false|||LUE
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3530,3533|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|SIMPLE_SEGMENT|3530,3533|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3530,3533|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3534,3540|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Event|Event|SIMPLE_SEGMENT|3541,3549|false|false|false|||strength
Finding|Idea or Concept|SIMPLE_SEGMENT|3541,3549|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3565,3572|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|plantar
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3574,3581|false|false|false|C1525443|W flexion|flexion
Event|Event|SIMPLE_SEGMENT|3574,3581|false|false|false|||flexion
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3574,3581|false|false|false|C0231452||flexion
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3595,3600|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3595,3600|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3595,3612|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3601,3612|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Functional Concept|SIMPLE_SEGMENT|3622,3627|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|SIMPLE_SEGMENT|3628,3633|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|3628,3633|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3635,3644|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|3652,3655|false|false|false|||LLE
Event|Event|SIMPLE_SEGMENT|3663,3668|false|false|false|||touch
Finding|Mental Process|SIMPLE_SEGMENT|3663,3668|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3663,3668|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3663,3668|false|false|false|C0152054|Therapeutic Touch|touch
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3663,3678|false|false|false|C0702221|Touch sensation|touch sensation
Event|Event|SIMPLE_SEGMENT|3669,3678|false|false|false|||sensation
Finding|Finding|SIMPLE_SEGMENT|3669,3678|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|SIMPLE_SEGMENT|3669,3678|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|SIMPLE_SEGMENT|3669,3678|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|3682,3693|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Health Care Activity|SIMPLE_SEGMENT|3730,3739|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|SIMPLE_SEGMENT|3740,3744|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3740,3744|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3759,3764|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3759,3764|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3759,3764|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|3765,3768|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|3773,3776|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|3773,3776|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3773,3776|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|3783,3786|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|3783,3786|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|3783,3786|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3783,3786|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3792,3795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3792,3795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|3803,3806|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|3803,3806|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|3803,3806|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3803,3806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|3803,3806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|3810,3813|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|3810,3813|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|3810,3813|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|3810,3813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|3810,3813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3810,3813|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|3819,3823|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3819,3823|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|3850,3853|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3870,3875|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|3870,3875|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3870,3875|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|3888,3894|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|SIMPLE_SEGMENT|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|SIMPLE_SEGMENT|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|3912,3915|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|SIMPLE_SEGMENT|3912,3915|false|false|false|||Eos
Finding|Gene or Genome|SIMPLE_SEGMENT|3912,3915|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4014,4019|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4014,4019|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4014,4019|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4024,4027|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|4024,4027|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4024,4027|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4049,4054|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4049,4054|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4049,4054|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|4049,4062|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4049,4062|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4049,4062|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4055,4062|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|4055,4062|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4055,4062|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|4055,4062|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4055,4062|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4055,4062|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4110,4114|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4140,4145|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4140,4145|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4140,4145|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|SIMPLE_SEGMENT|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Event|Event|SIMPLE_SEGMENT|4171,4174|false|false|false|||TRF
Finding|Gene or Genome|SIMPLE_SEGMENT|4171,4174|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Event|Event|SIMPLE_SEGMENT|4190,4194|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4190,4194|false|false|false|C0587081|Laboratory test finding|LABS
Event|Event|SIMPLE_SEGMENT|4195,4202|false|false|false|||IMAGING
Finding|Finding|SIMPLE_SEGMENT|4195,4202|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4195,4202|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|SIMPLE_SEGMENT|4210,4218|false|false|false|||received
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4222,4227|false|false|false|C2316467|Packed red blood cells|pRBCs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4222,4227|false|false|false|C2316467|Packed red blood cells|pRBCs
Event|Event|SIMPLE_SEGMENT|4222,4227|false|false|false|||pRBCs
Event|Event|SIMPLE_SEGMENT|4231,4240|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|4231,4240|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4256,4261|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4256,4261|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4256,4261|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4262,4265|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4270,4273|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4270,4273|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4270,4273|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4280,4283|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4280,4283|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4280,4283|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4280,4283|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4289,4292|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4289,4292|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4300,4303|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4300,4303|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4300,4303|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4300,4303|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4300,4303|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4307,4310|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4307,4310|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4307,4310|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4307,4310|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4307,4310|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4307,4310|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4316,4320|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4316,4320|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4347,4350|false|false|false|C0201617|Primed lymphocyte test|Plt
Finding|Gene or Genome|SIMPLE_SEGMENT|4368,4373|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|4374,4381|false|false|false|||episode
Drug|Food|SIMPLE_SEGMENT|4385,4391|false|false|false|C0009237|Coffee|coffee
Event|Event|SIMPLE_SEGMENT|4385,4391|false|false|false|||coffee
Finding|Finding|SIMPLE_SEGMENT|4385,4405|false|false|false|C0278002;C1510416|Coffee ground vomiting;Vomit contains coffee grounds (finding)|coffee ground emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|4385,4405|false|false|false|C0278002;C1510416|Coffee ground vomiting;Vomit contains coffee grounds (finding)|coffee ground emesis
Event|Event|SIMPLE_SEGMENT|4399,4405|false|false|false|||emesis
Finding|Body Substance|SIMPLE_SEGMENT|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|SIMPLE_SEGMENT|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4419,4424|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4419,4424|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4419,4424|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4425,4428|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4433,4436|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4433,4436|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4433,4436|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4443,4446|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4443,4446|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4443,4446|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4443,4446|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4452,4455|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4452,4455|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4463,4466|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4463,4466|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4463,4466|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4463,4466|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4463,4466|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4470,4473|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4470,4473|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4470,4473|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4470,4473|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4470,4473|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4470,4473|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4479,4483|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4479,4483|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4510,4513|false|false|false|C0201617|Primed lymphocyte test|Plt
Event|Event|SIMPLE_SEGMENT|4523,4531|false|false|false|||received
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4566,4571|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|4566,4571|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|4566,4571|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|4572,4575|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|4580,4583|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4580,4583|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4580,4583|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|4591,4594|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4591,4594|false|false|false|C0019046|Hemoglobin|Hgb
Event|Event|SIMPLE_SEGMENT|4591,4594|false|false|false|||Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|4591,4594|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4591,4594|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4602,4605|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4602,4605|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|4613,4616|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|4613,4616|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|4613,4616|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4613,4616|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4613,4616|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|4620,4623|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|4620,4623|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|4620,4623|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|4620,4623|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|4620,4623|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4620,4623|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|4629,4633|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4629,4633|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|4660,4663|false|false|false|C0201617|Primed lymphocyte test|Plt
Anatomy|Body Location or Region|SIMPLE_SEGMENT|4683,4688|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|4683,4688|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4683,4698|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4689,4698|false|false|false|C0015385|Limb structure|extremity
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4699,4706|false|false|false|C0554756|Doppler studies|doppler
Event|Event|SIMPLE_SEGMENT|4707,4708|false|false|false|||U
Event|Event|SIMPLE_SEGMENT|4711,4721|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|4711,4721|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|4711,4721|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Attribute|Clinical Attribute|SIMPLE_SEGMENT|4729,4733|false|false|false|C4318566|Deep Resection Margin|Deep
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4729,4751|false|false|false|C0149871|Deep Vein Thrombosis|Deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4734,4740|false|false|false|C0042449|Veins|venous
Finding|Finding|SIMPLE_SEGMENT|4734,4751|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|4734,4751|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Event|Event|SIMPLE_SEGMENT|4741,4751|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|4741,4751|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4769,4778|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4779,4785|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4787,4792|false|false|false|C0042449|Veins|veins
Event|Event|SIMPLE_SEGMENT|4787,4792|false|false|false|||veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4787,4792|false|false|false|C0398102|Procedure on vein|veins
Finding|Functional Concept|SIMPLE_SEGMENT|4818,4823|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|4834,4838|false|false|false|C0010709|Cyst|cyst
Event|Event|SIMPLE_SEGMENT|4834,4838|false|false|false|||cyst
Finding|Body Substance|SIMPLE_SEGMENT|4834,4838|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|SIMPLE_SEGMENT|4834,4838|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Event|Event|SIMPLE_SEGMENT|4842,4845|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|4842,4845|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|4856,4862|true|false|false|||amount
Finding|Intellectual Product|SIMPLE_SEGMENT|4856,4862|true|false|false|C1561574|Amount class - Amount|amount
Drug|Biologically Active Substance|SIMPLE_SEGMENT|4866,4873|true|false|false|C0018927|Hematin|hematin
Drug|Organic Chemical|SIMPLE_SEGMENT|4866,4873|true|false|false|C0018927|Hematin|hematin
Event|Event|SIMPLE_SEGMENT|4866,4873|true|false|false|||hematin
Event|Event|SIMPLE_SEGMENT|4882,4890|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|4882,4890|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|4882,4893|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|4894,4904|true|false|false|||ulceration
Finding|Pathologic Function|SIMPLE_SEGMENT|4894,4904|true|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Event|Event|SIMPLE_SEGMENT|4908,4914|true|false|false|||active
Event|Event|SIMPLE_SEGMENT|4916,4924|true|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|4916,4924|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|4925,4929|false|false|false|||seen
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|4954,4961|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4954,4961|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|4954,4961|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Event|Event|SIMPLE_SEGMENT|4954,4961|false|false|false|||stomach
Finding|Finding|SIMPLE_SEGMENT|4954,4961|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|4954,4961|false|false|false|C0872393|Procedure on stomach|stomach
Event|Event|SIMPLE_SEGMENT|4979,4987|false|false|false|||deformed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|4997,5005|false|false|false|C0041834|Erythema|erythema
Event|Event|SIMPLE_SEGMENT|4997,5005|false|false|false|||erythema
Event|Event|SIMPLE_SEGMENT|5023,5034|false|false|false|||ulcerations
Finding|Pathologic Function|SIMPLE_SEGMENT|5023,5034|false|false|false|C0041582|Ulcer|ulcerations
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5042,5049|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5042,5049|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5042,5049|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|SIMPLE_SEGMENT|5042,5049|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5042,5049|false|false|false|C0872393|Procedure on stomach|stomach
Event|Event|SIMPLE_SEGMENT|5050,5060|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5050,5060|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5050,5065|false|false|false|C0332290|Consistent with|consistent with
Event|Event|SIMPLE_SEGMENT|5066,5072|false|false|false|||severe
Finding|Finding|SIMPLE_SEGMENT|5066,5072|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|SIMPLE_SEGMENT|5066,5072|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5074,5083|false|false|false|C0017152|Gastritis|gastritis
Event|Event|SIMPLE_SEGMENT|5074,5083|false|false|false|||gastritis
Event|Event|SIMPLE_SEGMENT|5095,5103|true|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|5095,5103|true|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|5104,5114|true|false|false|||identified
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5116,5122|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|Medium
Drug|Substance|SIMPLE_SEGMENT|5116,5122|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|Medium
Finding|Finding|SIMPLE_SEGMENT|5116,5122|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|Medium
Finding|Intellectual Product|SIMPLE_SEGMENT|5116,5122|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|Medium
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|5123,5136|false|false|false|C3489393|Hiatal Hernia|hiatal hernia
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|5130,5136|false|false|false|C0019270|Hernia|hernia
Event|Event|SIMPLE_SEGMENT|5130,5136|false|false|false|||hernia
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5137,5145|false|false|false|C0041834|Erythema|Erythema
Event|Event|SIMPLE_SEGMENT|5137,5145|false|false|false|||Erythema
Event|Event|SIMPLE_SEGMENT|5162,5173|false|false|false|||ulcerations
Finding|Pathologic Function|SIMPLE_SEGMENT|5162,5173|false|false|false|C0041582|Ulcer|ulcerations
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5181,5189|false|false|false|C0013303|Duodenum|duodenal
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5181,5194|false|false|false|C0227300|Duodenal ampulla|duodenal bulb
Anatomy|Anatomical Structure|SIMPLE_SEGMENT|5190,5194|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5190,5194|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Event|Event|SIMPLE_SEGMENT|5196,5206|false|false|false|||consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5196,5206|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|SIMPLE_SEGMENT|5196,5211|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5212,5222|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5212,5222|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Event|Event|SIMPLE_SEGMENT|5212,5222|false|false|false|||duodenitis
Event|Event|SIMPLE_SEGMENT|5241,5244|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5241,5244|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|5254,5258|false|false|false|||part
Finding|Idea or Concept|SIMPLE_SEGMENT|5254,5258|false|false|false|C1552020|Role Class - part|part
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5266,5274|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|SIMPLE_SEGMENT|5266,5274|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Finding|Functional Concept|SIMPLE_SEGMENT|5280,5284|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5280,5300|false|false|false|C0230330|Left upper extremity|Left upper extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5285,5300|false|false|false|C1140618|Upper Extremity|upper extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5291,5300|false|false|false|C0015385|Limb structure|extremity
Event|Event|SIMPLE_SEGMENT|5301,5311|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|5301,5311|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|5301,5311|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5301,5311|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Event|Event|SIMPLE_SEGMENT|5312,5322|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5312,5322|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5312,5322|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|5333,5341|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5333,5341|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5333,5344|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5345,5349|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5345,5354|true|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5345,5365|true|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5350,5354|true|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|5350,5365|true|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|5355,5365|true|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|5355,5365|true|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|SIMPLE_SEGMENT|5373,5377|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5385,5394|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|SIMPLE_SEGMENT|5401,5407|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|SIMPLE_SEGMENT|5401,5407|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Functional Concept|SIMPLE_SEGMENT|5408,5416|false|true|false|C0332253|Evolving|evolving
Event|Event|SIMPLE_SEGMENT|5417,5425|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|5417,5425|false|true|false|C0018944|Hematoma|hematoma
Finding|Functional Concept|SIMPLE_SEGMENT|5433,5437|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5433,5455|false|false|false|C0694648|left antecubital fossa|left antecubital fossa
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5438,5449|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5438,5455|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|5450,5455|false|false|false|C0836913|Fossa|fossa
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5463,5470|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5463,5470|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|SIMPLE_SEGMENT|5466,5470|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|5466,5470|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5466,5470|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5466,5470|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|5475,5483|false|false|false|C0009924|Contrast Media|contrast
Event|Event|SIMPLE_SEGMENT|5475,5483|false|false|false|||contrast
Event|Event|SIMPLE_SEGMENT|5484,5494|false|false|false|||IMPRESSION
Finding|Intellectual Product|SIMPLE_SEGMENT|5484,5494|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|SIMPLE_SEGMENT|5484,5494|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|SIMPLE_SEGMENT|5502,5510|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|5502,5510|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|5502,5513|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|SIMPLE_SEGMENT|5514,5519|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|5520,5530|true|false|false|||infarction
Finding|Pathologic Function|SIMPLE_SEGMENT|5520,5530|true|false|false|C0021308|Infarction|infarction
Event|Event|SIMPLE_SEGMENT|5532,5542|true|false|false|||hemorrhage
Finding|Pathologic Function|SIMPLE_SEGMENT|5532,5542|true|false|false|C0019080|Hemorrhage|hemorrhage
Disorder|Injury or Poisoning|SIMPLE_SEGMENT|5545,5554|false|false|false|C0016658|Fracture|fractures
Event|Event|SIMPLE_SEGMENT|5545,5554|false|false|false|||fractures
Finding|Finding|SIMPLE_SEGMENT|5545,5554|false|false|false|C4554413|Fractured|fractures
Finding|Body Substance|SIMPLE_SEGMENT|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|SIMPLE_SEGMENT|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|SIMPLE_SEGMENT|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|SIMPLE_SEGMENT|5558,5567|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|SIMPLE_SEGMENT|5568,5572|false|false|false|||LABS
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5568,5572|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5586,5591|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5586,5591|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5586,5591|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|SIMPLE_SEGMENT|5592,5595|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|SIMPLE_SEGMENT|5600,5603|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5600,5603|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5600,5603|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5610,5613|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5610,5613|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|SIMPLE_SEGMENT|5610,5613|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5610,5613|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5619,5622|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5619,5622|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|SIMPLE_SEGMENT|5630,5633|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|SIMPLE_SEGMENT|5630,5633|false|false|false|||MCV
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5630,5633|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5630,5633|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5630,5633|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|SIMPLE_SEGMENT|5637,5640|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5637,5640|false|false|false|C0600370|methacholine|MCH
Event|Event|SIMPLE_SEGMENT|5637,5640|false|false|false|||MCH
Finding|Gene or Genome|SIMPLE_SEGMENT|5637,5640|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|SIMPLE_SEGMENT|5637,5640|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5637,5640|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|SIMPLE_SEGMENT|5646,5650|false|false|false|||MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5646,5650|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5677,5680|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5697,5702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5697,5702|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5697,5702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5703,5706|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5723,5728|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5723,5728|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5723,5728|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5723,5736|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5723,5736|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5723,5736|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5729,5736|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|SIMPLE_SEGMENT|5729,5736|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5729,5736|false|false|false|C0017725|glucose|Glucose
Event|Event|SIMPLE_SEGMENT|5729,5736|false|false|false|||Glucose
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|5729,5736|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5729,5736|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5783,5787|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5783,5787|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5783,5787|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5810,5815|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5810,5815|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5810,5815|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5810,5823|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|SIMPLE_SEGMENT|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|SIMPLE_SEGMENT|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|SIMPLE_SEGMENT|5816,5823|false|false|false|||Calcium
Finding|Physiologic Function|SIMPLE_SEGMENT|5816,5823|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|5816,5823|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5856,5861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|SIMPLE_SEGMENT|5856,5861|false|false|false|||BLOOD
Finding|Body Substance|SIMPLE_SEGMENT|5856,5861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|SIMPLE_SEGMENT|5862,5866|false|false|false|C0013618|edetic acid|EDTA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|5862,5866|false|false|false|C0013618|edetic acid|EDTA
Event|Event|SIMPLE_SEGMENT|5862,5866|false|false|false|||EDTA
Finding|Intellectual Product|SIMPLE_SEGMENT|5873,5878|false|false|false|C4050216;C4724718|BRIEF Health Literacy Screening Tool;Behavior Rating Inventory of Executive Function|Brief
Finding|Idea or Concept|SIMPLE_SEGMENT|5879,5887|false|false|false|C1547192|Organization unit type - Hospital|Hospital
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5879,5894|false|false|false|C0488549||Hospital Course
Finding|Finding|SIMPLE_SEGMENT|5879,5894|false|false|false|C0489547|Hospital course|Hospital Course
Finding|Classification|SIMPLE_SEGMENT|5896,5906|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|5896,5906|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Event|Event|SIMPLE_SEGMENT|5907,5916|false|false|false|||Providers
Finding|Functional Concept|SIMPLE_SEGMENT|5907,5916|false|false|false|C1138603|Provider|Providers
Event|Event|SIMPLE_SEGMENT|5920,5921|false|false|false|||_
Event|Event|SIMPLE_SEGMENT|5932,5943|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|5932,5943|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5948,5951|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|5948,5951|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|5948,5951|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|5948,5951|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|5948,5951|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5953,5956|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|5953,5956|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|5959,5962|false|false|false|||HLD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5970,5973|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|5974,5979|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|5974,5982|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|5984,5987|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|SIMPLE_SEGMENT|5984,5987|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|5984,5987|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|SIMPLE_SEGMENT|6001,6005|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6019,6026|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6019,6033|false|false|false|C0015801;C4299099|Lower extremity>Femoral artery;Structure of femoral artery|femoral artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6027,6033|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|6027,6033|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|6036,6044|false|false|false|||presents
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6050,6055|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6050,6055|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6050,6064|false|false|false|C0230443|Structure of left lower leg|lower left leg
Finding|Functional Concept|SIMPLE_SEGMENT|6056,6060|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6056,6064|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|6056,6073|false|false|false|C2219779|numbness of left leg|left leg numbness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6061,6064|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|6061,6073|false|false|false|C0857160|Numbness in leg|leg numbness
Event|Event|SIMPLE_SEGMENT|6065,6073|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|6065,6073|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|6065,6073|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6078,6082|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|6078,6082|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|6078,6082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|6078,6082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|6085,6090|false|false|false|||found
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6120,6123|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6120,6123|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6120,6123|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|6120,6123|false|false|false|||DVT
Event|Event|SIMPLE_SEGMENT|6133,6140|false|false|false|||treated
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|6157,6161|false|false|false|||drip
Finding|Pathologic Function|SIMPLE_SEGMENT|6175,6183|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|6184,6190|false|false|false|||events
Event|Event|SIMPLE_SEGMENT|6184,6190|false|false|false|C0441471|Event|events
Event|Event|SIMPLE_SEGMENT|6213,6222|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|6232,6235|false|false|false|||GIB
Event|Event|SIMPLE_SEGMENT|6244,6247|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6244,6247|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|6257,6265|false|false|false|||followed
Event|Event|SIMPLE_SEGMENT|6284,6293|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6284,6293|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|6307,6311|false|false|false|||drip
Event|Event|SIMPLE_SEGMENT|6316,6323|false|false|false|||stopped
Finding|Intellectual Product|SIMPLE_SEGMENT|6328,6332|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|6334,6344|false|false|false|||re-started
Drug|Food|SIMPLE_SEGMENT|6354,6360|false|false|false|C0009237|Coffee|coffee
Event|Event|SIMPLE_SEGMENT|6368,6374|false|false|false|||emesis
Finding|Body Substance|SIMPLE_SEGMENT|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|SIMPLE_SEGMENT|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Event|Event|SIMPLE_SEGMENT|6375,6383|false|false|false|||resolved
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6389,6395|false|false|false|C0489144||stools
Finding|Body Substance|SIMPLE_SEGMENT|6389,6395|false|false|false|C0015733|Feces|stools
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|6408,6416|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|6408,6416|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|6408,6416|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|6408,6416|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|6436,6441|true|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|6436,6441|true|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|6436,6441|true|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|6446,6451|true|false|false|||found
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|6455,6461|true|false|false|C1272938|Rectal Dosage Form|rectal
Event|Event|SIMPLE_SEGMENT|6455,6461|true|false|false|||rectal
Finding|Finding|SIMPLE_SEGMENT|6455,6461|true|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Finding|Functional Concept|SIMPLE_SEGMENT|6455,6461|true|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Event|Event|SIMPLE_SEGMENT|6463,6467|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|6463,6467|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|6463,6467|false|false|false|C0582103|Medical Examination|exam
Event|Event|SIMPLE_SEGMENT|6472,6476|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|6482,6493|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6482,6493|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|6482,6493|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|SIMPLE_SEGMENT|6503,6511|false|false|false|||deferred
Finding|Body Substance|SIMPLE_SEGMENT|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6546,6555|false|false|false|||developed
Finding|Functional Concept|SIMPLE_SEGMENT|6558,6562|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6558,6566|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6563,6566|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6563,6566|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|6563,6566|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|6567,6575|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|6567,6575|false|false|false|C0018944|Hematoma|hematoma
Drug|Biologically Active Substance|SIMPLE_SEGMENT|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|6599,6606|false|false|false|||stopped
Finding|Intellectual Product|SIMPLE_SEGMENT|6611,6615|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|SIMPLE_SEGMENT|6616,6626|false|false|false|||re-started
Event|Event|SIMPLE_SEGMENT|6636,6644|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|6636,6644|false|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|6649,6653|false|false|false|||felt
Event|Event|SIMPLE_SEGMENT|6661,6667|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|6661,6667|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|SIMPLE_SEGMENT|6677,6681|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Event|Event|SIMPLE_SEGMENT|6682,6688|false|false|false|||radial
Finding|Conceptual Entity|SIMPLE_SEGMENT|6682,6688|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Finding|SIMPLE_SEGMENT|6692,6696|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|SIMPLE_SEGMENT|6710,6715|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|6710,6715|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6710,6725|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6716,6725|false|false|false|C0015385|Limb structure|extremity
Drug|Food|SIMPLE_SEGMENT|6743,6749|false|false|false|C5890763||pulses
Event|Event|SIMPLE_SEGMENT|6743,6749|false|false|false|||pulses
Finding|Physiologic Function|SIMPLE_SEGMENT|6743,6749|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|SIMPLE_SEGMENT|6743,6749|false|false|false|C0034107|Pulse taking|pulses
Event|Event|SIMPLE_SEGMENT|6761,6770|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|6761,6770|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|SIMPLE_SEGMENT|6772,6782|false|false|false|||Hematology
Finding|Intellectual Product|SIMPLE_SEGMENT|6772,6782|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|Hematology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6772,6782|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|Hematology
Event|Event|SIMPLE_SEGMENT|6788,6797|false|false|false|||consulted
Finding|Body Substance|SIMPLE_SEGMENT|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|6816,6825|false|false|false|||developed
Finding|Functional Concept|SIMPLE_SEGMENT|6828,6832|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6828,6836|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|6833,6836|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|6833,6836|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|6833,6836|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|6837,6845|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|6837,6845|false|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|6871,6881|false|false|false|||uptitrated
Event|Event|SIMPLE_SEGMENT|6895,6910|false|false|false|||recommendations
Finding|Idea or Concept|SIMPLE_SEGMENT|6895,6910|false|false|false|C0034866|Recommendation|recommendations
Event|Event|SIMPLE_SEGMENT|6934,6941|false|false|false|||bridged
Drug|Organic Chemical|SIMPLE_SEGMENT|6945,6953|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|6945,6953|false|false|false|C0699129|Coumadin|coumadin
Event|Event|SIMPLE_SEGMENT|6945,6953|false|false|false|||coumadin
Attribute|Clinical Attribute|SIMPLE_SEGMENT|6962,6965|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|6962,6965|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|6962,6965|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|6962,6965|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Event|Event|SIMPLE_SEGMENT|6969,6978|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|6969,6978|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|6996,7006|false|false|false|||discharged
Event|Event|SIMPLE_SEGMENT|7010,7015|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7010,7015|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|SIMPLE_SEGMENT|7042,7045|false|false|false|||see
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7063,7070|false|false|false|C3854081||problem
Event|Event|SIMPLE_SEGMENT|7063,7070|false|false|false|||problem
Finding|Finding|SIMPLE_SEGMENT|7063,7070|false|false|false|C0033213|Problem|problem
Event|Event|SIMPLE_SEGMENT|7086,7093|false|false|false|||summary
Finding|Intellectual Product|SIMPLE_SEGMENT|7086,7093|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|summary
Finding|Idea or Concept|SIMPLE_SEGMENT|7099,7111|false|false|false|C1548597|Marketing basis - Transitional|transitional
Event|Event|SIMPLE_SEGMENT|7112,7118|false|false|false|||issues
Event|Event|SIMPLE_SEGMENT|7248,7259|false|false|false|||significant
Finding|Idea or Concept|SIMPLE_SEGMENT|7248,7259|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7264,7267|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|7264,7267|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|7264,7267|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|7264,7267|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|7264,7267|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7269,7272|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|7269,7272|false|false|false|||HTN
Event|Event|SIMPLE_SEGMENT|7274,7277|false|false|false|||HLD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7285,7288|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|7285,7288|false|false|false|||CKD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7290,7295|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|SIMPLE_SEGMENT|7290,7298|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7300,7303|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Event|Event|SIMPLE_SEGMENT|7300,7303|false|false|false|||PVD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7300,7303|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|SIMPLE_SEGMENT|7317,7321|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7322,7348|false|false|false|C0447106|Superficial femoral artery|superficial femoral artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7334,7341|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7334,7348|false|false|false|C0015801;C4299099|Lower extremity>Femoral artery;Structure of femoral artery|femoral artery
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7342,7348|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|7342,7348|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Event|Event|SIMPLE_SEGMENT|7352,7361|false|false|false|||presented
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7367,7372|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|7367,7372|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7367,7381|false|false|false|C0230443|Structure of left lower leg|lower Left leg
Finding|Functional Concept|SIMPLE_SEGMENT|7373,7377|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7373,7381|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|Left leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|7373,7390|false|true|false|C2219779|numbness of left leg|Left leg numbness
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7378,7381|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|SIMPLE_SEGMENT|7378,7390|false|false|false|C0857160|Numbness in leg|leg numbness
Event|Event|SIMPLE_SEGMENT|7382,7390|false|false|false|||numbness
Finding|Finding|SIMPLE_SEGMENT|7382,7390|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|SIMPLE_SEGMENT|7382,7390|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7395,7399|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|7395,7399|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|7395,7399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7395,7399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|7406,7415|false|false|false|||yesterday
Event|Event|SIMPLE_SEGMENT|7431,7441|false|false|false|||ultrasound
Finding|Functional Concept|SIMPLE_SEGMENT|7431,7441|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|SIMPLE_SEGMENT|7431,7441|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|7431,7441|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7452,7457|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|SIMPLE_SEGMENT|7452,7457|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7452,7469|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7458,7469|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Event|Event|SIMPLE_SEGMENT|7470,7477|false|false|false|||showing
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7489,7498|false|false|false|C0751438|Posterior pituitary disease|posterior
Event|Event|SIMPLE_SEGMENT|7489,7498|false|false|false|||posterior
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7489,7511|false|false|false|C0226832|Structure of posterior tibial vein|posterior tibial veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7499,7505|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7499,7511|false|false|false|C0447138|Tibial vein structure|tibial veins
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|7506,7511|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7506,7511|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|SIMPLE_SEGMENT|7512,7515|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7512,7515|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7512,7515|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|SIMPLE_SEGMENT|7512,7517|false|false|false|||DVT's
Event|Event|SIMPLE_SEGMENT|7522,7532|false|false|false|||Unprovoked
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7543,7547|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|SIMPLE_SEGMENT|7543,7547|false|false|false|||DVTs
Finding|Intellectual Product|SIMPLE_SEGMENT|7552,7560|true|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Event|Event|SIMPLE_SEGMENT|7561,7566|true|false|false|||signs
Finding|Finding|SIMPLE_SEGMENT|7561,7566|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|SIMPLE_SEGMENT|7561,7566|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|SIMPLE_SEGMENT|7577,7586|true|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|7577,7586|true|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Cell or Molecular Dysfunction|SIMPLE_SEGMENT|7603,7611|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Event|Event|SIMPLE_SEGMENT|7603,7611|false|false|false|||positive
Finding|Classification|SIMPLE_SEGMENT|7603,7611|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|SIMPLE_SEGMENT|7603,7611|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|7622,7626|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Event|Event|SIMPLE_SEGMENT|7622,7626|false|false|false|||DVTs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7637,7641|false|false|false|C2598155||Pain
Finding|Functional Concept|SIMPLE_SEGMENT|7637,7641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|7637,7641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|SIMPLE_SEGMENT|7647,7655|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|7647,7655|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|SIMPLE_SEGMENT|7656,7664|false|false|false|||improved
Event|Event|SIMPLE_SEGMENT|7668,7683|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|7668,7683|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|7668,7683|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7668,7683|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Body Substance|SIMPLE_SEGMENT|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|7697,7704|false|false|false|||bridged
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|7719,7723|false|false|false|||drip
Drug|Organic Chemical|SIMPLE_SEGMENT|7727,7738|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7727,7738|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|SIMPLE_SEGMENT|7727,7738|false|false|false|||therapeutic
Finding|Functional Concept|SIMPLE_SEGMENT|7727,7738|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|SIMPLE_SEGMENT|7727,7738|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7727,7738|false|false|false|C0087111|Therapeutic procedure|therapeutic
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|7739,7747|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|7739,7747|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7739,7747|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|7739,7747|false|false|false|||warfarin
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7753,7756|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|7753,7756|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7753,7756|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|7753,7756|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Attribute|Clinical Attribute|SIMPLE_SEGMENT|7753,7761|false|false|false|C5142654|Coagulation tissue factor induced.INR goal|INR goal
Event|Event|SIMPLE_SEGMENT|7757,7761|false|false|false|||goal
Finding|Idea or Concept|SIMPLE_SEGMENT|7757,7761|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|SIMPLE_SEGMENT|7757,7761|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Functional Concept|SIMPLE_SEGMENT|7767,7770|false|false|false|C0678226;C3146286|Due;Due to|Due
Finding|Idea or Concept|SIMPLE_SEGMENT|7767,7770|false|false|false|C0678226;C3146286|Due;Due to|Due
Disorder|Neoplastic Process|SIMPLE_SEGMENT|7804,7807|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|7804,7807|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7804,7807|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|7832,7842|true|false|false|||hematology
Finding|Intellectual Product|SIMPLE_SEGMENT|7832,7842|true|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|7832,7842|true|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Event|Event|SIMPLE_SEGMENT|7847,7856|true|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|7872,7878|true|false|false|||workup
Event|Event|SIMPLE_SEGMENT|7883,7889|true|false|false|||deemed
Event|Event|SIMPLE_SEGMENT|7891,7900|true|false|false|||necessary
Drug|Biologically Active Substance|SIMPLE_SEGMENT|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|SIMPLE_SEGMENT|7929,7939|false|false|false|||uptitrated
Event|Event|SIMPLE_SEGMENT|7943,7949|false|false|false|||needed
Drug|Organic Chemical|SIMPLE_SEGMENT|7952,7963|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|7952,7963|false|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|SIMPLE_SEGMENT|7952,7963|false|false|false|||Clopidogrel
Event|Event|SIMPLE_SEGMENT|7968,7975|false|false|false|||stopped
Finding|Classification|SIMPLE_SEGMENT|7980,7990|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|7980,7990|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|7991,8003|false|false|false|||cardiologist
Finding|Body Substance|SIMPLE_SEGMENT|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8019,8023|false|false|false|||need
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8024,8027|false|false|false|C1114365||age
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8024,8027|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|SIMPLE_SEGMENT|8024,8027|false|false|false|C0162574|Glycation End Products, Advanced|age
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8040,8046|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8040,8056|false|false|false|C0199230|Screening for cancer|cancer screening
Event|Event|SIMPLE_SEGMENT|8047,8056|false|false|false|||screening
Finding|Finding|SIMPLE_SEGMENT|8047,8056|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|SIMPLE_SEGMENT|8047,8056|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|SIMPLE_SEGMENT|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|SIMPLE_SEGMENT|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Event|Event|SIMPLE_SEGMENT|8067,8078|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8067,8078|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|8067,8078|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|SIMPLE_SEGMENT|8084,8093|false|false|false|||mammogram
Finding|Finding|SIMPLE_SEGMENT|8084,8093|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8084,8093|false|false|false|C0024671|Mammography|mammogram
Finding|Body Substance|SIMPLE_SEGMENT|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8108,8114|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|8137,8152|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|8137,8152|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|8137,8152|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8137,8152|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|8153,8163|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|8153,8163|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|8153,8163|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|8175,8183|false|false|false|||continue
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8184,8195|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|8187,8195|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|8187,8195|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8187,8195|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|8187,8195|false|false|false|||warfarin
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8224,8232|false|false|false|C0203057|Upper gastrointestinal tract series|Upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|8224,8238|false|false|false|C0041909|Upper gastrointestinal hemorrhage|Upper GI bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|8230,8238|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|8233,8238|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|8233,8238|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|SIMPLE_SEGMENT|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8248,8257|false|false|false|||developed
Event|Event|SIMPLE_SEGMENT|8260,8267|false|false|false|||episode
Finding|Gene or Genome|SIMPLE_SEGMENT|8268,8273|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Food|SIMPLE_SEGMENT|8274,8280|false|false|false|C0009237|Coffee|coffee
Event|Event|SIMPLE_SEGMENT|8274,8280|false|false|false|||coffee
Event|Event|SIMPLE_SEGMENT|8289,8295|false|false|false|||emesis
Finding|Body Substance|SIMPLE_SEGMENT|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|SIMPLE_SEGMENT|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|SIMPLE_SEGMENT|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|8313,8317|false|false|false|||drip
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8323,8326|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|8323,8326|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8323,8326|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8347,8352|false|false|false|C2316467|Packed red blood cells|pRBCs
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8347,8352|false|false|false|C2316467|Packed red blood cells|pRBCs
Event|Event|SIMPLE_SEGMENT|8347,8352|false|false|false|||pRBCs
Event|Event|SIMPLE_SEGMENT|8357,8366|false|false|false|||consulted
Event|Event|SIMPLE_SEGMENT|8371,8374|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8371,8374|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|8375,8381|false|false|false|||showed
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8382,8391|false|false|false|C0017152|Gastritis|gastritis
Event|Event|SIMPLE_SEGMENT|8382,8391|false|false|false|||gastritis
Event|Event|SIMPLE_SEGMENT|8396,8407|false|false|false|||superficial
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8409,8417|false|false|false|C0333307|Superficial ulcer|erosions
Event|Event|SIMPLE_SEGMENT|8409,8417|false|false|false|||erosions
Finding|Pathologic Function|SIMPLE_SEGMENT|8409,8417|false|false|false|C1959609|Erosion lesion|erosions
Event|Event|SIMPLE_SEGMENT|8432,8440|true|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|8432,8440|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Functional Concept|SIMPLE_SEGMENT|8442,8452|false|false|false|C0444507|Incidental|Incidental
Finding|Finding|SIMPLE_SEGMENT|8442,8460|false|false|false|C0743997|Incidental Findings|Incidental finding
Event|Event|SIMPLE_SEGMENT|8453,8460|false|false|false|||finding
Finding|Finding|SIMPLE_SEGMENT|8453,8460|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|SIMPLE_SEGMENT|8453,8460|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|8464,8470|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Drug|Substance|SIMPLE_SEGMENT|8464,8470|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Event|Event|SIMPLE_SEGMENT|8464,8470|false|false|false|||medium
Finding|Finding|SIMPLE_SEGMENT|8464,8470|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Intellectual Product|SIMPLE_SEGMENT|8464,8470|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Disorder|Acquired Abnormality|SIMPLE_SEGMENT|8478,8491|false|false|false|C3489393|Hiatal Hernia|hiatal hernia
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|8485,8491|false|false|false|C0019270|Hernia|hernia
Event|Event|SIMPLE_SEGMENT|8485,8491|false|false|false|||hernia
Finding|Body Substance|SIMPLE_SEGMENT|8493,8498|false|false|false|C0015733|Feces|Stool
Drug|Immunologic Factor|SIMPLE_SEGMENT|8509,8516|false|false|false|C0003320|Antigens|antigen
Event|Event|SIMPLE_SEGMENT|8509,8516|false|false|false|||antigen
Event|Event|SIMPLE_SEGMENT|8521,8529|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|8521,8529|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|8521,8529|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|8521,8529|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|8535,8546|false|false|false|||recommended
Finding|Finding|SIMPLE_SEGMENT|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8568,8571|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|8568,8571|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|8568,8571|false|false|false|C0871125|Prepulse Inhibition|PPI
Finding|Functional Concept|SIMPLE_SEGMENT|8576,8580|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8581,8592|false|false|false|C1549091|Antecubital|antecubital
Event|Event|SIMPLE_SEGMENT|8593,8601|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|8593,8601|false|false|false|C0018944|Hematoma|hematoma
Finding|Body Substance|SIMPLE_SEGMENT|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|8611,8620|false|false|false|||developed
Finding|Gene or Genome|SIMPLE_SEGMENT|8621,8626|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|SIMPLE_SEGMENT|8627,8631|false|false|false|||left
Finding|Functional Concept|SIMPLE_SEGMENT|8627,8631|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|8633,8644|false|false|false|C1549091|Antecubital|antecubital
Event|Event|SIMPLE_SEGMENT|8645,8653|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|8645,8653|false|true|false|C0018944|Hematoma|hematoma
Finding|Mental Process|SIMPLE_SEGMENT|8657,8664|false|false|false|C0542559|contextual factors|setting
Event|Event|SIMPLE_SEGMENT|8668,8678|false|false|false|||phlebotomy
Finding|Finding|SIMPLE_SEGMENT|8668,8678|false|false|false|C2183248|diagnostic service sources phlebotomy|phlebotomy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|8668,8678|false|false|false|C0031555;C0190979;C0684257|Phlebotomy, therapeutic (separate procedure);Venesection;Venous blood sampling|phlebotomy
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|8668,8678|false|false|false|C0031555;C0190979;C0684257|Phlebotomy, therapeutic (separate procedure);Venesection;Venous blood sampling|phlebotomy
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8683,8686|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|SIMPLE_SEGMENT|8683,8686|false|false|false|||PTT
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8683,8686|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Event|Event|SIMPLE_SEGMENT|8697,8704|false|false|false|||heparin
Disorder|Neoplastic Process|SIMPLE_SEGMENT|8705,8708|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8705,8708|false|false|false|C0991568|Drops - Drug Form|gtt
Event|Event|SIMPLE_SEGMENT|8705,8708|false|false|false|||gtt
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8705,8708|false|false|false|C0017741|Glucose tolerance test|gtt
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|SIMPLE_SEGMENT|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Event|Event|SIMPLE_SEGMENT|8722,8726|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|8733,8741|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|8733,8741|false|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|8742,8750|false|false|false|||improved
Finding|Functional Concept|SIMPLE_SEGMENT|8752,8758|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Event|Event|SIMPLE_SEGMENT|8769,8775|false|false|false|||stable
Finding|Intellectual Product|SIMPLE_SEGMENT|8769,8775|false|false|false|C1547311|Patient Condition Code - Stable|stable
Event|Event|SIMPLE_SEGMENT|8781,8786|false|false|false|||Acute
Finding|Intellectual Product|SIMPLE_SEGMENT|8781,8786|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|8790,8793|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|8790,8793|false|false|false|||CKD
Attribute|Clinical Attribute|SIMPLE_SEGMENT|8794,8799|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|SIMPLE_SEGMENT|8794,8802|false|false|false|C0441772|Stage level 4|Stage IV
Finding|Body Substance|SIMPLE_SEGMENT|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|SIMPLE_SEGMENT|8817,8827|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|SIMPLE_SEGMENT|8817,8827|false|false|false|C0010294|creatinine|creatinine
Event|Event|SIMPLE_SEGMENT|8817,8827|false|false|false|||creatinine
Finding|Physiologic Function|SIMPLE_SEGMENT|8817,8827|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|8817,8827|false|false|false|C0201975|Creatinine measurement|creatinine
Event|Event|SIMPLE_SEGMENT|8839,8848|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|8839,8848|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|8854,8862|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|SIMPLE_SEGMENT|8854,8862|false|false|false|||baseline
Finding|Idea or Concept|SIMPLE_SEGMENT|8854,8862|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|SIMPLE_SEGMENT|8872,8880|false|false|false|||Improved
Event|Event|SIMPLE_SEGMENT|8886,8895|false|false|false|||hydration
Finding|Finding|SIMPLE_SEGMENT|8886,8895|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|SIMPLE_SEGMENT|8886,8895|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Event|Event|SIMPLE_SEGMENT|8897,8901|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8897,8901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8897,8901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8897,8901|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|8903,8908|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8903,8908|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8903,8908|false|false|false|||lasix
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|8913,8923|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8913,8923|false|false|false|C0065374|lisinopril|lisinopril
Event|Event|SIMPLE_SEGMENT|8913,8923|false|false|false|||lisinopril
Event|Event|SIMPLE_SEGMENT|8939,8943|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|8945,8949|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|8945,8949|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|8945,8949|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|8945,8949|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|8950,8955|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|8950,8955|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|8956,8965|false|false|false|||restarted
Event|Event|SIMPLE_SEGMENT|8970,8979|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|8970,8979|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9010,9016|false|false|false|C0002871|Anemia|Anemia
Event|Event|SIMPLE_SEGMENT|9010,9016|false|false|false|||Anemia
Finding|Body Substance|SIMPLE_SEGMENT|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|SIMPLE_SEGMENT|9018,9029|false|false|false|C0332310|Has patient|Patient has
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9041,9047|false|false|false|C0002871|Anemia|anemia
Event|Event|SIMPLE_SEGMENT|9041,9047|false|false|false|||anemia
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|9049,9055|false|false|false|C1272938|Rectal Dosage Form|Rectal
Finding|Finding|SIMPLE_SEGMENT|9049,9055|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Finding|Functional Concept|SIMPLE_SEGMENT|9049,9055|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9049,9060|false|false|false|C0199900|Rectal examination|Rectal exam
Event|Event|SIMPLE_SEGMENT|9056,9060|false|false|false|||exam
Finding|Functional Concept|SIMPLE_SEGMENT|9056,9060|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|SIMPLE_SEGMENT|9056,9060|false|false|false|C0582103|Medical Examination|exam
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|9072,9078|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|SIMPLE_SEGMENT|9072,9078|false|false|false|C0018302|guaiac|guaiac
Event|Event|SIMPLE_SEGMENT|9072,9078|false|false|false|||guaiac
Event|Event|SIMPLE_SEGMENT|9079,9087|false|false|false|||negative
Finding|Classification|SIMPLE_SEGMENT|9079,9087|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|SIMPLE_SEGMENT|9079,9087|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|SIMPLE_SEGMENT|9079,9087|false|false|false|C5237010|Expression Negative|negative
Event|Event|SIMPLE_SEGMENT|9097,9104|false|false|false|||treated
Event|Event|SIMPLE_SEGMENT|9110,9117|false|false|false|||aransep
Finding|Finding|SIMPLE_SEGMENT|9121,9125|false|false|false|C5575035|Well (answer to question)|well
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Hormone|SIMPLE_SEGMENT|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Event|Event|SIMPLE_SEGMENT|9130,9133|false|false|false|||EPO
Finding|Gene or Genome|SIMPLE_SEGMENT|9130,9133|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|EPO
Finding|Intellectual Product|SIMPLE_SEGMENT|9130,9133|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|EPO
Event|Event|SIMPLE_SEGMENT|9135,9143|false|false|false|||Etiology
Finding|Conceptual Entity|SIMPLE_SEGMENT|9135,9143|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|SIMPLE_SEGMENT|9135,9143|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Finding|SIMPLE_SEGMENT|9144,9150|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|9144,9150|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|SIMPLE_SEGMENT|9151,9158|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|SIMPLE_SEGMENT|9151,9158|false|false|false|||related
Finding|Finding|SIMPLE_SEGMENT|9151,9158|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|SIMPLE_SEGMENT|9151,9158|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Event|Event|SIMPLE_SEGMENT|9162,9172|false|false|false|||underlying
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9173,9176|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Event|Event|SIMPLE_SEGMENT|9173,9176|false|false|false|||CKD
Event|Event|SIMPLE_SEGMENT|9197,9205|false|false|false|||consider
Finding|Pathologic Function|SIMPLE_SEGMENT|9211,9219|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|9214,9219|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|9214,9219|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|9221,9232|false|false|false|C0332310|Has patient|patient has
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9233,9242|false|false|false|C0017152|Gastritis|gastritis
Event|Event|SIMPLE_SEGMENT|9233,9242|false|false|false|||gastritis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9243,9253|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Disorder|Neoplastic Process|SIMPLE_SEGMENT|9243,9253|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Event|Event|SIMPLE_SEGMENT|9243,9253|false|false|false|||duodenitis
Event|Event|SIMPLE_SEGMENT|9258,9261|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9258,9261|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|9269,9277|true|false|false|||evidence
Finding|Idea or Concept|SIMPLE_SEGMENT|9269,9277|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|SIMPLE_SEGMENT|9269,9280|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|SIMPLE_SEGMENT|9288,9296|true|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|9288,9296|true|false|false|C0019080|Hemorrhage|bleeding
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9298,9302|false|false|false|C0337439|Iron measurement|Iron
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|9298,9310|false|false|false|C2079295|iron studies|Iron studies
Event|Event|SIMPLE_SEGMENT|9303,9310|false|false|false|||studies
Procedure|Research Activity|SIMPLE_SEGMENT|9303,9310|false|false|false|C0947630|Scientific Study|studies
Event|Event|SIMPLE_SEGMENT|9317,9323|false|false|false|||normal
Event|Event|SIMPLE_SEGMENT|9336,9340|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9336,9340|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9336,9340|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9336,9340|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|9341,9351|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9341,9351|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|9341,9351|false|false|false|||furosemide
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9356,9366|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9356,9366|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|SIMPLE_SEGMENT|9356,9366|false|false|false|||Lisinopril
Event|Event|SIMPLE_SEGMENT|9372,9376|false|false|false|||held
Event|Event|SIMPLE_SEGMENT|9380,9389|false|false|false|||admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|9380,9389|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Pathologic Function|SIMPLE_SEGMENT|9411,9419|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|9414,9419|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|9414,9419|false|false|false|C0019080|Hemorrhage|bleed
Drug|Organic Chemical|SIMPLE_SEGMENT|9421,9431|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9421,9431|false|false|false|C0054836|carvedilol|Carvedilol
Event|Event|SIMPLE_SEGMENT|9421,9431|false|false|false|||Carvedilol
Event|Event|SIMPLE_SEGMENT|9436,9444|false|false|false|||nifedine
Event|Event|SIMPLE_SEGMENT|9450,9454|false|false|false|||held
Finding|Mental Process|SIMPLE_SEGMENT|9459,9466|false|false|false|C0542559|contextual factors|setting
Finding|Idea or Concept|SIMPLE_SEGMENT|9479,9484|false|false|false|C1552828|Table Frame - above|above
Drug|Organic Chemical|SIMPLE_SEGMENT|9487,9497|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9487,9497|false|false|false|C0028066|nifedipine|Nifedipine
Event|Event|SIMPLE_SEGMENT|9502,9511|false|false|false|||restarted
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9521,9524|false|false|false|C4546282|Body integrity dysphoria|bid
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9521,9524|false|false|false|C1530795|BID protein, human|bid
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9521,9524|false|false|false|C1530795|BID protein, human|bid
Event|Event|SIMPLE_SEGMENT|9521,9524|false|false|false|||bid
Finding|Gene or Genome|SIMPLE_SEGMENT|9521,9524|false|false|false|C1332410|BID gene|bid
Drug|Organic Chemical|SIMPLE_SEGMENT|9529,9534|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9529,9534|false|false|false|C0699992|Lasix|lasix
Event|Event|SIMPLE_SEGMENT|9529,9534|false|false|false|||lasix
Event|Event|SIMPLE_SEGMENT|9539,9548|false|false|false|||decreased
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9577,9580|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9577,9580|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|SIMPLE_SEGMENT|9577,9580|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|SIMPLE_SEGMENT|9577,9580|false|false|false|||CAD
Finding|Gene or Genome|SIMPLE_SEGMENT|9577,9580|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|SIMPLE_SEGMENT|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9598,9601|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Event|Event|SIMPLE_SEGMENT|9598,9601|false|false|false|||BMS
Anatomy|Body Location or Region|SIMPLE_SEGMENT|9630,9633|false|false|false|C0449201|PER (body structure)|Per
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9630,9633|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Per
Event|Event|SIMPLE_SEGMENT|9630,9633|false|false|false|||Per
Finding|Functional Concept|SIMPLE_SEGMENT|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Gene or Genome|SIMPLE_SEGMENT|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Intellectual Product|SIMPLE_SEGMENT|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Event|Event|SIMPLE_SEGMENT|9635,9646|false|false|false|||discussions
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|9635,9646|false|false|false|C0557061|Discussion (procedure)|discussions
Finding|Body Substance|SIMPLE_SEGMENT|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|SIMPLE_SEGMENT|9686,9697|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9686,9697|false|false|false|C0070166|clopidogrel|clopidogrel
Event|Event|SIMPLE_SEGMENT|9686,9697|false|false|false|||clopidogrel
Event|Event|SIMPLE_SEGMENT|9702,9706|false|false|false|||held
Finding|Pathologic Function|SIMPLE_SEGMENT|9713,9721|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|9716,9721|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|9716,9721|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|SIMPLE_SEGMENT|9726,9736|false|false|false|||initiation
Finding|Functional Concept|SIMPLE_SEGMENT|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|SIMPLE_SEGMENT|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|SIMPLE_SEGMENT|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|9740,9748|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9740,9748|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9740,9748|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|9740,9748|false|false|false|||warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|9751,9756|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9751,9756|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|9767,9771|false|false|false|||held
Finding|Idea or Concept|SIMPLE_SEGMENT|9775,9780|false|false|false|C1552828|Table Frame - above|above
Event|Event|SIMPLE_SEGMENT|9786,9795|false|false|false|||restarted
Event|Event|SIMPLE_SEGMENT|9799,9808|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|9799,9808|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|9825,9829|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9825,9829|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9825,9829|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9825,9829|false|false|false|C1553498|home health encounter|Home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|SIMPLE_SEGMENT|9830,9833|false|false|false|||ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|9830,9833|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|9835,9841|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9835,9841|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Event|Event|SIMPLE_SEGMENT|9835,9841|false|false|false|||statin
Finding|Gene or Genome|SIMPLE_SEGMENT|9835,9841|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Organic Chemical|SIMPLE_SEGMENT|9847,9857|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9847,9857|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|SIMPLE_SEGMENT|9847,9857|false|false|false|||carvedilol
Event|Event|SIMPLE_SEGMENT|9863,9872|false|false|false|||continued
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9878,9881|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|SIMPLE_SEGMENT|9878,9881|false|false|false|||HTN
Drug|Organic Chemical|SIMPLE_SEGMENT|9883,9893|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|9883,9893|false|false|false|C0028066|nifedipine|Nifedipine
Event|Event|SIMPLE_SEGMENT|9883,9893|false|false|false|||Nifedipine
Event|Event|SIMPLE_SEGMENT|9898,9907|false|false|false|||decreased
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9916,9919|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9916,9919|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9916,9919|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9916,9919|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9916,9919|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|9930,9933|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|9930,9933|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|9930,9933|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|9930,9933|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|9930,9933|false|false|false|C1332410|BID gene|BID
Finding|Pathologic Function|SIMPLE_SEGMENT|9950,9958|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|SIMPLE_SEGMENT|9950,9967|false|false|false|C1970394|Bleeding episodes|bleeding episodes
Event|Event|SIMPLE_SEGMENT|9959,9967|false|false|false|||episodes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|9979,9984|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|9979,9984|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|9979,9984|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|SIMPLE_SEGMENT|9979,9994|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Event|Event|SIMPLE_SEGMENT|9985,9994|false|false|false|||pressures
Finding|Finding|SIMPLE_SEGMENT|9985,9994|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|9985,9994|false|false|false|C0033095||pressures
Event|Event|SIMPLE_SEGMENT|9996,10000|false|false|false|||Home
Finding|Idea or Concept|SIMPLE_SEGMENT|9996,10000|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|SIMPLE_SEGMENT|9996,10000|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|SIMPLE_SEGMENT|9996,10000|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|SIMPLE_SEGMENT|10002,10012|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10002,10012|false|false|false|C0054836|carvedilol|carvedilol
Event|Event|SIMPLE_SEGMENT|10002,10012|false|false|false|||carvedilol
Event|Event|SIMPLE_SEGMENT|10013,10022|false|false|false|||continued
Finding|Body Substance|SIMPLE_SEGMENT|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|10034,10044|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10034,10044|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|10034,10044|false|false|false|||nifedipine
Event|Event|SIMPLE_SEGMENT|10049,10058|false|false|false|||decreased
Finding|Intellectual Product|SIMPLE_SEGMENT|10080,10085|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|SIMPLE_SEGMENT|10080,10091|false|false|false|C0333276|Acute hemorrhage|acute bleed
Event|Event|SIMPLE_SEGMENT|10086,10091|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10086,10091|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10096,10100|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Drug|Organic Chemical|SIMPLE_SEGMENT|10112,10117|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10112,10117|false|false|false|C0699992|Lasix|Lasix
Event|Event|SIMPLE_SEGMENT|10112,10117|false|false|false|||Lasix
Event|Event|SIMPLE_SEGMENT|10122,10131|false|false|false|||decreased
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10163,10171|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10163,10180|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Event|Event|SIMPLE_SEGMENT|10172,10180|false|false|false|||Mellitus
Event|Event|SIMPLE_SEGMENT|10182,10188|false|false|false|||Stable
Finding|Intellectual Product|SIMPLE_SEGMENT|10182,10188|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Event|Event|SIMPLE_SEGMENT|10192,10196|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|10192,10196|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10192,10196|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10192,10196|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|SIMPLE_SEGMENT|10212,10219|false|false|false|||insulin
Finding|Gene or Genome|SIMPLE_SEGMENT|10212,10219|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|10212,10219|false|false|false|C0202098|Insulin measurement|insulin
Event|Event|SIMPLE_SEGMENT|10224,10231|false|false|false|||bedtime
Finding|Idea or Concept|SIMPLE_SEGMENT|10236,10248|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|SIMPLE_SEGMENT|10249,10255|false|false|false|||ISSUES
Finding|Body Substance|SIMPLE_SEGMENT|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|SIMPLE_SEGMENT|10289,10293|false|false|false|||work
Event|Occupational Activity|SIMPLE_SEGMENT|10289,10293|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10289,10296|false|false|false|C0750430|Work-up|work up
Event|Event|SIMPLE_SEGMENT|10307,10316|false|false|false|||screening
Finding|Finding|SIMPLE_SEGMENT|10307,10316|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|SIMPLE_SEGMENT|10307,10316|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|SIMPLE_SEGMENT|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|SIMPLE_SEGMENT|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Event|Event|SIMPLE_SEGMENT|10318,10329|false|false|false|||colonoscopy
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10318,10329|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|SIMPLE_SEGMENT|10318,10329|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Event|Event|SIMPLE_SEGMENT|10347,10356|false|false|false|||mammogram
Finding|Finding|SIMPLE_SEGMENT|10347,10356|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10347,10356|false|false|false|C0024671|Mammography|mammogram
Finding|Body Substance|SIMPLE_SEGMENT|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10372,10376|false|false|false|||need
Event|Event|SIMPLE_SEGMENT|10380,10388|false|false|false|||complete
Finding|Intellectual Product|SIMPLE_SEGMENT|10394,10398|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|SIMPLE_SEGMENT|10399,10405|false|false|false|||course
Finding|Finding|SIMPLE_SEGMENT|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|SIMPLE_SEGMENT|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|SIMPLE_SEGMENT|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Event|Event|SIMPLE_SEGMENT|10414,10418|false|false|false|||dose
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10420,10423|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Event|Event|SIMPLE_SEGMENT|10420,10423|false|false|false|||PPI
Finding|Physiologic Function|SIMPLE_SEGMENT|10420,10423|false|false|false|C0871125|Prepulse Inhibition|PPI
Event|Event|SIMPLE_SEGMENT|10425,10432|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|10438,10450|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10438,10450|false|false|false|C0081876|pantoprazole|pantoprazole
Event|Event|SIMPLE_SEGMENT|10438,10450|false|false|false|||pantoprazole
Event|Event|SIMPLE_SEGMENT|10479,10488|false|false|false|||projected
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10489,10492|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|SIMPLE_SEGMENT|10489,10492|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|SIMPLE_SEGMENT|10489,10492|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|SIMPLE_SEGMENT|10489,10492|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10506,10514|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|10506,10520|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10512,10520|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|10515,10520|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10515,10520|false|false|false|C0019080|Hemorrhage|bleed
Finding|Finding|SIMPLE_SEGMENT|10521,10527|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|SIMPLE_SEGMENT|10521,10527|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10534,10543|false|false|false|C0017152|Gastritis|gastritis
Event|Event|SIMPLE_SEGMENT|10534,10543|false|false|false|||gastritis
Finding|Body Substance|SIMPLE_SEGMENT|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|10557,10569|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|SIMPLE_SEGMENT|10557,10569|false|false|false|||hypertension
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10557,10581|false|false|false|C0684167|hypertensive agents|hypertension medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10570,10581|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10570,10581|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|10570,10581|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|10570,10581|false|false|false|C4284232|Medications|medications
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10583,10593|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10583,10593|false|false|false|C0065374|lisinopril|Lisinopril
Event|Event|SIMPLE_SEGMENT|10583,10593|false|false|false|||Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|10598,10608|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10598,10608|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|10598,10608|false|false|false|||nifedipine
Event|Event|SIMPLE_SEGMENT|10616,10620|false|false|false|||held
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|10628,10636|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|10628,10642|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10634,10642|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|10637,10642|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10637,10642|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|SIMPLE_SEGMENT|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|10656,10666|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10656,10666|false|false|false|C0016860|furosemide|furosemide
Event|Event|SIMPLE_SEGMENT|10656,10666|false|false|false|||furosemide
Event|Event|SIMPLE_SEGMENT|10671,10680|false|false|false|||decreased
Finding|Body Substance|SIMPLE_SEGMENT|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|SIMPLE_SEGMENT|10707,10717|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10707,10717|false|false|false|C0028066|nifedipine|nifedipine
Event|Event|SIMPLE_SEGMENT|10707,10717|false|false|false|||nifedipine
Event|Event|SIMPLE_SEGMENT|10722,10731|false|false|false|||decreased
Event|Event|SIMPLE_SEGMENT|10752,10757|false|false|false|||acute
Finding|Intellectual Product|SIMPLE_SEGMENT|10752,10757|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|SIMPLE_SEGMENT|10759,10764|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|10759,10764|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|10769,10773|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Finding|Body Substance|SIMPLE_SEGMENT|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|SIMPLE_SEGMENT|10799,10806|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|10810,10818|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10810,10818|false|false|false|C0699129|Coumadin|Coumadin
Event|Event|SIMPLE_SEGMENT|10810,10818|false|false|false|||Coumadin
Drug|Organic Chemical|SIMPLE_SEGMENT|10820,10831|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10820,10831|false|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|SIMPLE_SEGMENT|10820,10831|false|false|false|||Clopidogrel
Event|Event|SIMPLE_SEGMENT|10836,10843|false|false|false|||stopped
Anatomy|Body System|SIMPLE_SEGMENT|10849,10859|false|false|false|C0007226|Cardiovascular system|cardiology
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|SIMPLE_SEGMENT|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|SIMPLE_SEGMENT|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|SIMPLE_SEGMENT|10861,10864|false|false|false|C1412553|ARSA gene|ASA
Event|Event|SIMPLE_SEGMENT|10874,10883|false|false|false|||continued
Attribute|Clinical Attribute|SIMPLE_SEGMENT|10894,10901|false|false|false|C2741676||address
Event|Event|SIMPLE_SEGMENT|10894,10901|false|false|false|||address
Finding|Intellectual Product|SIMPLE_SEGMENT|10894,10901|false|false|false|C0376649;C1442065;C1547327;C1578436;C1578437;C4319699|Address;Address (property);Address Data Type;Addresses (publication format);MDF Attribute Type - Address;Value type - Address|address
Finding|Body Substance|SIMPLE_SEGMENT|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|10912,10916|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10912,10916|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10912,10916|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|10912,10928|false|false|false|C2242846|home environment (history)|home environment
Event|Event|SIMPLE_SEGMENT|10917,10928|false|false|false|||environment
Finding|Finding|SIMPLE_SEGMENT|10933,10937|false|false|false|C0085639|Falls|fall
Finding|Finding|SIMPLE_SEGMENT|10933,10942|false|false|false|C1268740|At increased risk for falls|fall risk
Event|Event|SIMPLE_SEGMENT|10938,10942|false|false|false|||risk
Finding|Idea or Concept|SIMPLE_SEGMENT|10938,10942|false|false|false|C0035647|Risk|risk
Event|Event|SIMPLE_SEGMENT|10950,10956|false|false|false|||recent
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|10958,10962|false|false|false|C0077275|triptorelin|trip
Drug|Hormone|SIMPLE_SEGMENT|10958,10962|false|false|false|C0077275|triptorelin|trip
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|10958,10962|false|false|false|C0077275|triptorelin|trip
Event|Event|SIMPLE_SEGMENT|10958,10962|false|false|false|||trip
Finding|Gene or Genome|SIMPLE_SEGMENT|10958,10962|false|false|false|C1416921;C2239819;C2608049;C4085339|LRRFIP1 gene;PIK3IP1 gene;TRAIP gene;TRAIP wt Allele|trip
Phenomenon|Phenomenon or Process|SIMPLE_SEGMENT|10958,10962|false|false|false|C0221188|Tripping|trip
Finding|Finding|SIMPLE_SEGMENT|10964,10971|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|SIMPLE_SEGMENT|10967,10971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|10967,10971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|10967,10971|false|false|false|C1553498|home health encounter|home
Finding|Finding|SIMPLE_SEGMENT|10976,10979|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|10976,10979|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Event|Event|SIMPLE_SEGMENT|10980,10995|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|10980,10995|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|10980,10995|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|10980,10995|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|11006,11012|false|false|false|||ensure
Finding|Body Substance|SIMPLE_SEGMENT|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|SIMPLE_SEGMENT|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|SIMPLE_SEGMENT|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|SIMPLE_SEGMENT|11013,11024|false|false|false|C0332310|Has patient|patient has
Finding|Classification|SIMPLE_SEGMENT|11025,11035|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|11025,11035|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|SIMPLE_SEGMENT|11036,11051|false|false|false|||anticoagulation
Finding|Finding|SIMPLE_SEGMENT|11036,11051|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|SIMPLE_SEGMENT|11036,11051|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11036,11051|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|SIMPLE_SEGMENT|11052,11058|false|false|false|||follow
Event|Event|SIMPLE_SEGMENT|11067,11077|false|false|false|||management
Event|Occupational Activity|SIMPLE_SEGMENT|11067,11077|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|SIMPLE_SEGMENT|11067,11077|false|false|false|C0376636|Disease Management|management
Event|Event|SIMPLE_SEGMENT|11083,11092|false|false|false|||discharge
Finding|Body Substance|SIMPLE_SEGMENT|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11083,11092|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|SIMPLE_SEGMENT|11098,11103|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|11098,11103|false|false|false|C0034991|Rehabilitation therapy|rehab
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11109,11120|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11109,11120|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|11109,11120|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11109,11120|false|false|false|C4284232|Medications|Medications
Finding|Finding|SIMPLE_SEGMENT|11109,11133|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|SIMPLE_SEGMENT|11124,11133|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|11124,11133|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11152,11162|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11152,11162|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|SIMPLE_SEGMENT|11152,11167|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|SIMPLE_SEGMENT|11163,11167|false|false|false|||list
Finding|Intellectual Product|SIMPLE_SEGMENT|11163,11167|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|SIMPLE_SEGMENT|11171,11179|false|false|false|||accurate
Drug|Organic Chemical|SIMPLE_SEGMENT|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|SIMPLE_SEGMENT|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|SIMPLE_SEGMENT|11184,11192|false|false|false|||complete
Finding|Functional Concept|SIMPLE_SEGMENT|11184,11192|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|SIMPLE_SEGMENT|11184,11192|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11197,11207|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11197,11207|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|11227,11238|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11227,11238|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Organic Chemical|SIMPLE_SEGMENT|11259,11271|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11259,11271|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|11281,11284|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|11289,11299|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11289,11299|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11311,11314|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11311,11314|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11311,11314|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11311,11314|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11311,11314|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11319,11330|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11319,11330|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|11350,11360|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11350,11360|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|SIMPLE_SEGMENT|11380,11390|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11380,11390|false|false|false|C0034665|ranitidine|Ranitidine
Finding|Gene or Genome|SIMPLE_SEGMENT|11407,11410|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|SIMPLE_SEGMENT|11411,11417|false|false|false|||reflux
Finding|Pathologic Function|SIMPLE_SEGMENT|11411,11417|false|false|false|C0232483|Reflux|reflux
Drug|Organic Chemical|SIMPLE_SEGMENT|11422,11429|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11422,11429|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|11449,11462|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11465,11468|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|11465,11468|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11483,11492|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|11497,11501|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|11516,11526|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11516,11526|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|SIMPLE_SEGMENT|11516,11526|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11539,11542|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11539,11542|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11539,11542|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11539,11542|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11539,11542|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11548,11561|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11548,11561|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Event|Event|SIMPLE_SEGMENT|11548,11561|false|false|false|||Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|11581,11584|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|11585,11590|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|11585,11590|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11585,11595|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11585,11595|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11591,11595|false|true|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|11591,11595|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|11591,11595|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11591,11595|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|11616,11622|false|false|false|||Dinner
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11616,11622|false|false|false|C4048877|Dinner|Dinner
Event|Event|SIMPLE_SEGMENT|11626,11635|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|11626,11635|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|11626,11647|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|SIMPLE_SEGMENT|11636,11647|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11636,11647|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|SIMPLE_SEGMENT|11636,11647|false|false|false|||Medications
Finding|Intellectual Product|SIMPLE_SEGMENT|11636,11647|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|SIMPLE_SEGMENT|11652,11663|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11652,11663|false|false|false|C0002144|allopurinol|Allopurinol
Event|Event|SIMPLE_SEGMENT|11686,11689|false|false|false|||DAY
Finding|Idea or Concept|SIMPLE_SEGMENT|11686,11689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|SIMPLE_SEGMENT|11686,11689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|SIMPLE_SEGMENT|11694,11701|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11694,11701|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|SIMPLE_SEGMENT|11721,11733|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11721,11733|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|SIMPLE_SEGMENT|11743,11746|false|false|false|||QPM
Drug|Organic Chemical|SIMPLE_SEGMENT|11751,11761|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11751,11761|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11773,11776|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11773,11776|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11773,11776|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11773,11776|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11773,11776|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|11796,11802|false|false|false|||Dinner
Finding|Daily or Recreational Activity|SIMPLE_SEGMENT|11796,11802|false|false|false|C4048877|Dinner|Dinner
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11806,11816|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11806,11816|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|SIMPLE_SEGMENT|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|SIMPLE_SEGMENT|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|SIMPLE_SEGMENT|11836,11849|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|11852,11855|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|SIMPLE_SEGMENT|11852,11855|false|false|false|||TAB
Drug|Organic Chemical|SIMPLE_SEGMENT|11869,11879|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11869,11879|false|false|false|C0028066|nifedipine|NIFEdipine
Event|Event|SIMPLE_SEGMENT|11869,11879|false|false|false|||NIFEdipine
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11892,11895|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11892,11895|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11892,11895|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11892,11895|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11892,11895|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|SIMPLE_SEGMENT|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|SIMPLE_SEGMENT|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|SIMPLE_SEGMENT|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|SIMPLE_SEGMENT|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11900,11909|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|SIMPLE_SEGMENT|11908,11909|false|false|false|||D
Event|Event|SIMPLE_SEGMENT|11914,11918|false|false|false|||UNIT
Drug|Organic Chemical|SIMPLE_SEGMENT|11933,11941|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11933,11941|false|false|false|C1692318|docusate|Docusate
Event|Event|SIMPLE_SEGMENT|11933,11941|false|false|false|||Docusate
Drug|Organic Chemical|SIMPLE_SEGMENT|11933,11948|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11933,11948|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|SIMPLE_SEGMENT|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|SIMPLE_SEGMENT|11942,11948|false|false|false|||Sodium
Finding|Physiologic Function|SIMPLE_SEGMENT|11942,11948|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|11942,11948|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|11959,11962|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|11959,11962|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|11959,11962|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|11959,11962|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|11959,11962|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|SIMPLE_SEGMENT|11968,11978|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|11968,11978|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|SIMPLE_SEGMENT|11993,12009|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|11993,12009|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12005,12009|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12005,12009|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12005,12009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12005,12009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|12015,12027|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12015,12027|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|SIMPLE_SEGMENT|12047,12052|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12047,12052|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|SIMPLE_SEGMENT|12063,12066|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|SIMPLE_SEGMENT|12063,12066|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|SIMPLE_SEGMENT|12063,12066|false|false|false|C1530795|BID protein, human|BID
Event|Event|SIMPLE_SEGMENT|12063,12066|false|false|false|||BID
Finding|Gene or Genome|SIMPLE_SEGMENT|12063,12066|false|false|false|C1332410|BID gene|BID
Event|Event|SIMPLE_SEGMENT|12067,12079|false|false|false|||constipation
Finding|Sign or Symptom|SIMPLE_SEGMENT|12067,12079|false|false|false|C0009806|Constipation|constipation
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Event|Event|SIMPLE_SEGMENT|12118,12122|false|false|false|||dose
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12138,12141|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|SIMPLE_SEGMENT|12138,12141|false|false|false|||INR
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12138,12141|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12138,12141|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|SIMPLE_SEGMENT|12147,12160|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12147,12160|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|SIMPLE_SEGMENT|12180,12183|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12184,12189|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|SIMPLE_SEGMENT|12184,12189|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12184,12194|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12184,12194|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12190,12194|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12190,12194|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12190,12194|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12190,12194|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|SIMPLE_SEGMENT|12200,12210|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12200,12210|false|false|false|C0016860|furosemide|Furosemide
Drug|Biomedical or Dental Material|SIMPLE_SEGMENT|12231,12243|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|12231,12243|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Event|Event|SIMPLE_SEGMENT|12231,12243|false|false|false|||Polyethylene
Drug|Organic Chemical|SIMPLE_SEGMENT|12231,12250|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12231,12250|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|12244,12250|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|12244,12250|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Event|Event|SIMPLE_SEGMENT|12244,12250|false|false|false|||Glycol
Drug|Organic Chemical|SIMPLE_SEGMENT|12270,12283|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12270,12283|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|SIMPLE_SEGMENT|12270,12283|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12270,12283|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|SIMPLE_SEGMENT|12302,12305|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12306,12310|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12306,12310|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12306,12310|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12306,12310|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|SIMPLE_SEGMENT|12314,12319|false|false|false|||fever
Finding|Finding|SIMPLE_SEGMENT|12314,12319|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|SIMPLE_SEGMENT|12314,12319|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|SIMPLE_SEGMENT|12324,12333|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12324,12333|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12324,12345|false|false|false|C4019243||Discharge Disposition
Finding|Finding|SIMPLE_SEGMENT|12324,12345|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12334,12345|false|false|false|C2926604||Disposition
Event|Event|SIMPLE_SEGMENT|12334,12345|false|false|false|||Disposition
Procedure|Health Care Activity|SIMPLE_SEGMENT|12334,12345|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|SIMPLE_SEGMENT|12347,12355|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|SIMPLE_SEGMENT|12347,12355|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|SIMPLE_SEGMENT|12347,12360|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|SIMPLE_SEGMENT|12356,12360|false|false|false|C1947933|care activity|Care
Event|Event|SIMPLE_SEGMENT|12356,12360|false|false|false|||Care
Finding|Finding|SIMPLE_SEGMENT|12356,12360|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|12356,12360|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|SIMPLE_SEGMENT|12363,12371|false|false|false|||Facility
Finding|Intellectual Product|SIMPLE_SEGMENT|12363,12371|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|SIMPLE_SEGMENT|12379,12388|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12379,12388|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|SIMPLE_SEGMENT|12379,12398|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12389,12398|false|false|false|C0945731||Diagnosis
Event|Event|SIMPLE_SEGMENT|12389,12398|false|false|false|||Diagnosis
Finding|Classification|SIMPLE_SEGMENT|12389,12398|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|SIMPLE_SEGMENT|12389,12398|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12389,12398|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12409,12413|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12409,12418|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12409,12429|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12409,12435|false|false|false|C0149871|Deep Vein Thrombosis|Deep vein thrombosis (DVT)
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12414,12418|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|12414,12429|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|12419,12429|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|12419,12429|false|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Location or Region|SIMPLE_SEGMENT|12431,12434|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12431,12434|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12431,12434|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12437,12446|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|SIMPLE_SEGMENT|12437,12446|false|false|false|||Secondary
Finding|Functional Concept|SIMPLE_SEGMENT|12437,12446|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12448,12456|false|false|false|C0203057|Upper gastrointestinal tract series|Upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|12448,12462|false|false|false|C0041909|Upper gastrointestinal hemorrhage|Upper GI bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|12454,12462|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|12457,12462|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|12457,12462|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12463,12468|false|false|false|C5779993|Left arm|L arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12465,12468|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|12465,12468|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|12465,12468|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|12469,12477|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|12469,12477|false|false|false|C0018944|Hematoma|hematoma
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12478,12506|false|false|false|C1510431|Superficial Thrombophlebitis|Superficial thrombophlebitis
Event|Event|SIMPLE_SEGMENT|12490,12506|false|false|false|||thrombophlebitis
Finding|Pathologic Function|SIMPLE_SEGMENT|12490,12506|false|false|false|C0040046|Thrombophlebitis|thrombophlebitis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12510,12521|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12510,12527|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|SIMPLE_SEGMENT|12522,12527|false|false|false|C0836913|Fossa|fossa
Event|Event|SIMPLE_SEGMENT|12528,12535|false|false|false|||Chronic
Finding|Intellectual Product|SIMPLE_SEGMENT|12528,12535|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|SIMPLE_SEGMENT|12528,12535|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12528,12550|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12536,12542|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|SIMPLE_SEGMENT|12536,12542|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|SIMPLE_SEGMENT|12536,12542|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12536,12542|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|12536,12542|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12536,12550|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12543,12550|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|12543,12550|false|false|false|||disease
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12552,12557|false|true|false|C1300072|Tumor stage|Stage
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12562,12589|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12573,12581|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12573,12589|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12582,12589|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|12582,12589|false|false|false|||disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12590,12598|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12590,12607|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12590,12615|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes mellitus type II
Finding|Gene or Genome|SIMPLE_SEGMENT|12608,12612|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|SIMPLE_SEGMENT|12608,12612|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12616,12624|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12616,12631|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12616,12639|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12625,12631|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|SIMPLE_SEGMENT|12625,12631|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12625,12639|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12632,12639|false|false|false|C0012634|Disease|disease
Event|Event|SIMPLE_SEGMENT|12632,12639|false|false|false|||disease
Event|Event|SIMPLE_SEGMENT|12643,12652|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12643,12652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12643,12652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12643,12652|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12643,12652|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12653,12662|false|false|false|C3864998||Condition
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12653,12662|false|false|false|C0012634|Disease|Condition
Event|Event|SIMPLE_SEGMENT|12653,12662|false|false|false|||Condition
Finding|Conceptual Entity|SIMPLE_SEGMENT|12653,12662|false|false|false|C1705253|Logical Condition|Condition
Finding|Mental Process|SIMPLE_SEGMENT|12664,12670|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12664,12677|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|SIMPLE_SEGMENT|12664,12677|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12671,12677|false|false|false|C5889824||Status
Finding|Idea or Concept|SIMPLE_SEGMENT|12671,12677|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|SIMPLE_SEGMENT|12679,12684|false|false|false|||Clear
Finding|Idea or Concept|SIMPLE_SEGMENT|12679,12684|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|SIMPLE_SEGMENT|12689,12697|false|false|false|||coherent
Finding|Finding|SIMPLE_SEGMENT|12689,12697|false|false|false|C4068804|Coherent|coherent
Event|Event|SIMPLE_SEGMENT|12699,12704|false|false|false|||Level
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12699,12721|false|false|false|C4050479||Level of Consciousness
Finding|Finding|SIMPLE_SEGMENT|12699,12721|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|SIMPLE_SEGMENT|12708,12721|false|false|false|||Consciousness
Finding|Finding|SIMPLE_SEGMENT|12708,12721|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|SIMPLE_SEGMENT|12708,12721|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12723,12728|false|false|false|C5890168||Alert
Drug|Organic Chemical|SIMPLE_SEGMENT|12723,12728|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|12723,12728|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|SIMPLE_SEGMENT|12723,12728|false|false|false|||Alert
Finding|Finding|SIMPLE_SEGMENT|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|SIMPLE_SEGMENT|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|SIMPLE_SEGMENT|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|SIMPLE_SEGMENT|12733,12744|false|false|false|||interactive
Finding|Functional Concept|SIMPLE_SEGMENT|12733,12744|false|false|false|C1704675|Interaction|interactive
Event|Event|SIMPLE_SEGMENT|12749,12758|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|12749,12758|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|12749,12758|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|12749,12758|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|12749,12758|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12749,12771|false|false|false|C3669312||Discharge Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12749,12771|false|false|false|C4282220|Discharge instructions|Discharge Instructions
Procedure|Health Care Activity|SIMPLE_SEGMENT|12749,12771|false|false|false|C2266673|hospital discharge instructions (treatment)|Discharge Instructions
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12759,12771|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|12759,12771|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|12759,12771|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions
Finding|Gene or Genome|SIMPLE_SEGMENT|12773,12777|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|SIMPLE_SEGMENT|12793,12801|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|12793,12801|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|12793,12801|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Event|SIMPLE_SEGMENT|12802,12808|false|false|false|||caring
Event|Event|SIMPLE_SEGMENT|12834,12842|false|false|false|||admitted
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12848,12851|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|SIMPLE_SEGMENT|12848,12860|false|true|false|C0581394|Swelling of lower limb|leg swelling
Event|Event|SIMPLE_SEGMENT|12852,12860|false|false|false|||swelling
Finding|Finding|SIMPLE_SEGMENT|12852,12860|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|SIMPLE_SEGMENT|12852,12860|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12865,12869|false|false|false|C2598155||pain
Event|Event|SIMPLE_SEGMENT|12865,12869|false|false|false|||pain
Finding|Functional Concept|SIMPLE_SEGMENT|12865,12869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|SIMPLE_SEGMENT|12865,12869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Indicator, Reagent, or Diagnostic Aid|SIMPLE_SEGMENT|12871,12881|false|false|false|C0358514|Diagnostic agents|Diagnostic
Finding|Functional Concept|SIMPLE_SEGMENT|12871,12881|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Finding|Intellectual Product|SIMPLE_SEGMENT|12871,12881|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12871,12881|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|Diagnostic
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|12871,12887|false|false|false|C0086143|Diagnostic tests|Diagnostic tests
Event|Event|SIMPLE_SEGMENT|12882,12887|false|false|false|||tests
Finding|Intellectual Product|SIMPLE_SEGMENT|12882,12887|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|SIMPLE_SEGMENT|12882,12887|false|false|false|C0022885|Laboratory Procedures|tests
Event|Event|SIMPLE_SEGMENT|12917,12926|false|false|false|||diagnosed
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12932,12936|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12932,12941|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12932,12952|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12937,12941|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|SIMPLE_SEGMENT|12937,12952|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Event|Event|SIMPLE_SEGMENT|12942,12952|false|false|false|||thrombosis
Finding|Pathologic Function|SIMPLE_SEGMENT|12942,12952|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|12954,12959|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|12954,12959|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|12954,12959|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|12954,12965|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clots
Event|Event|SIMPLE_SEGMENT|12960,12965|false|false|false|||clots
Finding|Pathologic Function|SIMPLE_SEGMENT|12960,12965|false|false|false|C0302148|Blood Clot|clots
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|12975,12979|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|SIMPLE_SEGMENT|12975,12979|false|false|false|C5781420||legs
Event|Event|SIMPLE_SEGMENT|12990,12997|false|false|false|||treated
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13003,13008|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13003,13008|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13003,13008|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Sign or Symptom|SIMPLE_SEGMENT|13009,13017|false|false|false|C0851184|Thinning Weight Loss|thinning
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13018,13029|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13018,13029|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|SIMPLE_SEGMENT|13018,13029|false|false|false|||medications
Finding|Intellectual Product|SIMPLE_SEGMENT|13018,13029|false|false|false|C4284232|Medications|medications
Event|Event|SIMPLE_SEGMENT|13045,13053|false|false|false|||continue
Finding|Finding|SIMPLE_SEGMENT|13054,13061|false|false|false|C4534363|At home|at home
Event|Event|SIMPLE_SEGMENT|13057,13061|false|false|false|||home
Finding|Idea or Concept|SIMPLE_SEGMENT|13057,13061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|SIMPLE_SEGMENT|13057,13061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|SIMPLE_SEGMENT|13057,13061|false|false|false|C1553498|home health encounter|home
Event|Event|SIMPLE_SEGMENT|13074,13081|false|false|false|||episode
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13085,13093|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|13085,13102|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|13091,13102|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleeding
Event|Event|SIMPLE_SEGMENT|13094,13102|false|false|false|||bleeding
Finding|Pathologic Function|SIMPLE_SEGMENT|13094,13102|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|SIMPLE_SEGMENT|13116,13120|false|false|false|||stay
Event|Event|SIMPLE_SEGMENT|13145,13152|false|false|false|||treated
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13158,13168|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|SIMPLE_SEGMENT|13158,13168|false|false|false|||medication
Finding|Intellectual Product|SIMPLE_SEGMENT|13158,13168|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|SIMPLE_SEGMENT|13178,13187|false|false|false|||underwent
Event|Event|SIMPLE_SEGMENT|13191,13194|false|false|false|||EGD
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13191,13194|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Event|Event|SIMPLE_SEGMENT|13200,13209|false|false|false|||developed
Finding|Functional Concept|SIMPLE_SEGMENT|13212,13216|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13212,13220|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|SIMPLE_SEGMENT|13217,13220|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|SIMPLE_SEGMENT|13217,13220|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|SIMPLE_SEGMENT|13217,13220|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|SIMPLE_SEGMENT|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|SIMPLE_SEGMENT|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|SIMPLE_SEGMENT|13221,13229|false|false|false|||hematoma
Finding|Pathologic Function|SIMPLE_SEGMENT|13221,13229|false|false|false|C0018944|Hematoma|hematoma
Event|Event|SIMPLE_SEGMENT|13234,13238|false|false|false|||well
Finding|Finding|SIMPLE_SEGMENT|13234,13238|false|false|false|C5575035|Well (answer to question)|well
Event|Event|SIMPLE_SEGMENT|13251,13255|false|false|false|||stay
Event|Event|SIMPLE_SEGMENT|13267,13274|false|false|false|||resolve
Event|Event|SIMPLE_SEGMENT|13282,13285|false|false|false|||own
Finding|Finding|SIMPLE_SEGMENT|13282,13285|false|false|false|C5939094|Own|own
Finding|Finding|SIMPLE_SEGMENT|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|SIMPLE_SEGMENT|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|SIMPLE_SEGMENT|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13307,13312|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13307,13312|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13307,13312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|SIMPLE_SEGMENT|13307,13318|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clots
Event|Event|SIMPLE_SEGMENT|13313,13318|false|false|false|||clots
Finding|Pathologic Function|SIMPLE_SEGMENT|13313,13318|false|false|false|C0302148|Blood Clot|clots
Event|Event|SIMPLE_SEGMENT|13329,13336|false|false|false|||started
Finding|Finding|SIMPLE_SEGMENT|13342,13345|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|SIMPLE_SEGMENT|13342,13345|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13346,13350|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Event|Event|SIMPLE_SEGMENT|13346,13350|false|false|false|||drug
Finding|Finding|SIMPLE_SEGMENT|13346,13350|false|false|false|C0740721|Drug problem|drug
Event|Event|SIMPLE_SEGMENT|13351,13357|false|false|false|||called
Drug|Hazardous or Poisonous Substance|SIMPLE_SEGMENT|13359,13367|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|SIMPLE_SEGMENT|13359,13367|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13359,13367|false|false|false|C0043031|warfarin|warfarin
Event|Event|SIMPLE_SEGMENT|13359,13367|false|false|false|||warfarin
Event|Event|SIMPLE_SEGMENT|13378,13382|false|false|false|||need
Disorder|Disease or Syndrome|SIMPLE_SEGMENT|13396,13401|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|SIMPLE_SEGMENT|13396,13401|false|false|false|||blood
Finding|Body Substance|SIMPLE_SEGMENT|13396,13401|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|SIMPLE_SEGMENT|13402,13409|false|false|false|||checked
Event|Event|SIMPLE_SEGMENT|13413,13419|false|false|false|||adjust
Event|Event|SIMPLE_SEGMENT|13425,13431|false|false|false|||dosing
Procedure|Diagnostic Procedure|SIMPLE_SEGMENT|13442,13450|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|SIMPLE_SEGMENT|13442,13456|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|13448,13456|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Event|Event|SIMPLE_SEGMENT|13451,13456|false|false|false|||bleed
Finding|Pathologic Function|SIMPLE_SEGMENT|13451,13456|false|false|false|C0019080|Hemorrhage|bleed
Event|Event|SIMPLE_SEGMENT|13467,13474|false|false|false|||started
Drug|Organic Chemical|SIMPLE_SEGMENT|13479,13491|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13479,13491|false|false|false|C0081876|pantoprazole|Pantoprazole
Event|Event|SIMPLE_SEGMENT|13519,13527|false|false|false|||continue
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13533,13537|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Event|Event|SIMPLE_SEGMENT|13533,13537|false|false|false|||drug
Finding|Finding|SIMPLE_SEGMENT|13533,13537|false|false|false|C0740721|Drug problem|drug
Event|Event|SIMPLE_SEGMENT|13545,13555|false|false|false|||outpatient
Finding|Classification|SIMPLE_SEGMENT|13545,13555|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|SIMPLE_SEGMENT|13545,13555|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|SIMPLE_SEGMENT|13622,13633|true|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13622,13633|true|false|false|C0070166|clopidogrel|Clopidogrel
Event|Event|SIMPLE_SEGMENT|13622,13633|true|false|false|||Clopidogrel
Drug|Organic Chemical|SIMPLE_SEGMENT|13635,13641|true|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|13635,13641|true|false|false|C0633084|Plavix|Plavix
Event|Event|SIMPLE_SEGMENT|13635,13641|true|false|false|||Plavix
Event|Event|SIMPLE_SEGMENT|13671,13683|false|false|false|||cardiologist
Event|Event|SIMPLE_SEGMENT|13695,13703|false|false|false|||pleasure
Finding|Intellectual Product|SIMPLE_SEGMENT|13695,13703|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|SIMPLE_SEGMENT|13695,13703|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|SIMPLE_SEGMENT|13711,13715|false|false|false|C1947933|care activity|care
Event|Event|SIMPLE_SEGMENT|13711,13715|false|false|false|||care
Finding|Finding|SIMPLE_SEGMENT|13711,13715|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|SIMPLE_SEGMENT|13711,13715|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|SIMPLE_SEGMENT|13732,13740|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|SIMPLE_SEGMENT|13741,13745|false|false|false|||stay
Event|Activity|SIMPLE_SEGMENT|13771,13775|false|false|false|C1947933|care activity|Care
Finding|Finding|SIMPLE_SEGMENT|13771,13775|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|SIMPLE_SEGMENT|13771,13775|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13771,13780|false|false|false|C4321316||Care Team
Finding|Finding|SIMPLE_SEGMENT|13771,13780|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|SIMPLE_SEGMENT|13783,13791|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|SIMPLE_SEGMENT|13792,13804|false|false|false|C3263700||Instructions
Event|Event|SIMPLE_SEGMENT|13792,13804|false|false|false|||Instructions
Finding|Intellectual Product|SIMPLE_SEGMENT|13792,13804|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

