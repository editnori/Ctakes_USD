 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|42,51|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|42,51|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|42,56|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|76,85|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|76,85|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|76,85|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|76,90|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|108,113|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|132,135|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|132,135|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|143,150|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|143,150|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|152,160|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|178,181|false|false|false|C0013343|Dyes|Dye
Event|Event|Allergies|178,181|false|false|false|||Dye
Drug|Biologically Active Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Element, Ion, or Isotope|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Drug|Pharmacologic Substance|Allergies|183,189|false|false|false|C0021968;C0885449|Iodine, Homeopathic preparation;iodine|Iodine
Event|Activity|Allergies|190,200|false|false|false|C2700400|Contain (action)|Containing
Finding|Functional Concept|Allergies|190,200|false|false|false|C0332256|Containing (qualifier value)|Containing
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,209|false|false|false|C0009924|Contrast Media|Contrast
Drug|Indicator, Reagent, or Diagnostic Aid|Allergies|201,215|false|false|false|C0009924|Contrast Media|Contrast Media
Anatomy|Tissue|Allergies|210,215|false|false|false|C0162867;C1254021|Media layer;Tunica Media|Media
Finding|Intellectual Product|Allergies|210,215|false|false|false|C0009458;C0677540|Communications Media;PAMS Media|Media
Drug|Organic Chemical|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Drug|Pharmacologic Substance|Allergies|218,227|false|false|false|C0030049|oxycodone|Oxycodone
Event|Event|Allergies|218,227|false|false|false|||Oxycodone
Procedure|Laboratory Procedure|Allergies|218,227|false|false|false|C0524222|Oxycodone measurement|Oxycodone
Drug|Organic Chemical|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Drug|Pharmacologic Substance|Allergies|231,241|false|false|false|C0055729|cilostazol|cilostazol
Event|Event|Allergies|231,241|false|false|false|||cilostazol
Drug|Organic Chemical|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Drug|Pharmacologic Substance|Allergies|244,255|false|false|false|C1569608|varenicline|Varenicline
Event|Event|Allergies|244,255|false|false|false|||Varenicline
Event|Event|Allergies|258,267|false|false|false|||Attending
Finding|Functional Concept|Allergies|258,267|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|293,302|false|false|false|||Shortness
Attribute|Clinical Attribute|Chief Complaint|293,312|false|false|false|C2707305||Shortness of Breath
Finding|Sign or Symptom|Chief Complaint|293,312|false|false|false|C0013404|Dyspnea|Shortness of Breath
Event|Event|Chief Complaint|306,312|false|false|false|||Breath
Finding|Body Substance|Chief Complaint|306,312|false|false|false|C0225386|Breath|Breath
Finding|Classification|Chief Complaint|316,321|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|322,330|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|334,352|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|343,352|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|343,352|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|343,352|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|343,352|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|343,352|false|false|false|C0184661|Interventional procedure|Procedure
Event|Event|Chief Complaint|354,355|false|false|false|||N
Event|Event|History of Present Illness|418,425|false|false|false|||history
Finding|Conceptual Entity|History of Present Illness|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|History of Present Illness|418,425|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|History of Present Illness|418,428|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|History of Present Illness|430,434|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|430,434|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|430,434|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|430,434|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|438,442|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|438,442|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|438,442|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|438,442|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|447,453|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|History of Present Illness|447,466|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|447,466|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|History of Present Illness|447,466|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|454,466|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|History of Present Illness|454,466|false|false|false|||fibrillation
Drug|Organic Chemical|History of Present Illness|470,478|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|History of Present Illness|470,478|false|false|false|C1831808|apixaban|apixaban
Event|Event|History of Present Illness|470,478|false|false|false|||apixaban
Disorder|Disease or Syndrome|History of Present Illness|480,492|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|480,492|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|495,498|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|495,498|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|495,498|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|History of Present Illness|495,498|false|false|false|||CAD
Finding|Gene or Genome|History of Present Illness|495,498|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|495,498|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|504,518|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|History of Present Illness|504,518|false|false|false|||hyperlipidemia
Finding|Finding|History of Present Illness|504,518|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|History of Present Illness|523,531|false|false|false|||presents
Event|Event|History of Present Illness|537,546|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|537,556|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|537,556|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|550,556|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|History of Present Illness|559,564|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|559,564|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|559,564|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|559,564|false|false|false|C0010200|Coughing|cough
Event|Event|History of Present Illness|570,578|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|570,578|false|false|false|C0043144|Wheezing|wheezing
Finding|Idea or Concept|History of Present Illness|587,590|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|History of Present Illness|587,590|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Body Substance|History of Present Illness|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|597,604|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|605,612|false|false|false|||reports
Finding|Finding|History of Present Illness|605,632|false|false|false|C4718286|Reports shortness of breath|reports shortness of breath
Event|Event|History of Present Illness|613,622|false|false|false|||shortness
Attribute|Clinical Attribute|History of Present Illness|613,632|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|613,632|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|626,632|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|History of Present Illness|644,649|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|644,649|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|644,649|false|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|644,649|false|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|669,672|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Finding|Gene or Genome|History of Present Illness|669,672|false|false|false|C0332575;C1414207;C1416378|DYRK3 gene;IK gene;Redness|red
Event|Event|History of Present Illness|681,687|false|false|false|||sputum
Finding|Body Substance|History of Present Illness|681,687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Intellectual Product|History of Present Illness|681,687|false|false|false|C0038056;C1546789;C1576419|Specimen Type - Sputum;Sputum|sputum
Finding|Sign or Symptom|History of Present Illness|693,701|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|719,726|false|false|false|||evening
Drug|Organic Chemical|History of Present Illness|748,757|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|History of Present Illness|748,757|false|false|false|C0001927|albuterol|albuterol
Event|Event|History of Present Illness|748,757|false|false|false|||albuterol
Drug|Organic Chemical|History of Present Illness|789,800|false|false|false|C0027235|ipratropium|ipratropium
Drug|Pharmacologic Substance|History of Present Illness|789,800|false|false|false|C0027235|ipratropium|ipratropium
Drug|Biomedical or Dental Material|History of Present Illness|801,805|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|History of Present Illness|801,805|false|false|false|||nebs
Drug|Organic Chemical|History of Present Illness|834,840|false|false|false|C0723011|Relief brand of phenylephrine|relief
Drug|Pharmacologic Substance|History of Present Illness|834,840|false|false|false|C0723011|Relief brand of phenylephrine|relief
Event|Event|History of Present Illness|834,840|false|false|false|||relief
Finding|Finding|History of Present Illness|834,840|false|false|false|C0564405|Feeling relief|relief
Event|Event|History of Present Illness|853,861|false|false|false|||increase
Event|Event|History of Present Illness|869,873|false|false|false|||flow
Phenomenon|Natural Phenomenon or Process|History of Present Illness|869,873|false|false|false|C0806140|Flow|flow
Finding|Idea or Concept|History of Present Illness|892,903|false|false|false|C0750502|Significant|significant
Event|Event|History of Present Illness|904,915|false|false|false|||improvement
Finding|Conceptual Entity|History of Present Illness|904,915|false|false|false|C2986411|Improvement|improvement
Finding|Finding|History of Present Illness|925,941|false|false|false|C3843777|Currently taking|currently taking
Event|Event|History of Present Illness|935,941|false|false|false|||taking
Drug|Hormone|History of Present Illness|951,961|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|951,961|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|951,961|false|false|false|C0032952|prednisone|prednisone
Event|Event|History of Present Illness|951,961|false|false|false|||prednisone
Event|Event|History of Present Illness|981,987|false|false|false|||taking
Drug|Organic Chemical|History of Present Illness|988,998|false|false|false|C0213771|tiotropium|tiotropium
Drug|Pharmacologic Substance|History of Present Illness|988,998|false|false|false|C0213771|tiotropium|tiotropium
Event|Event|History of Present Illness|988,998|false|false|false|||tiotropium
Drug|Organic Chemical|History of Present Illness|1004,1016|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|1004,1016|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|1004,1016|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|1004,1016|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|History of Present Illness|1018,1024|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|History of Present Illness|1018,1024|false|false|false|C0965130|Advair|advair
Event|Event|History of Present Illness|1018,1024|false|false|false|||advair
Finding|Finding|History of Present Illness|1028,1035|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|History of Present Illness|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1031,1035|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1031,1035|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|1039,1049|false|false|false|||prescribed
Event|Event|History of Present Illness|1055,1061|false|false|false|||denies
Event|Event|History of Present Illness|1062,1066|false|false|false|||sick
Finding|Sign or Symptom|History of Present Illness|1062,1066|false|false|false|C0221423|Illness (finding)|sick
Event|Event|History of Present Illness|1068,1076|false|false|false|||contacts
Procedure|Health Care Activity|History of Present Illness|1068,1076|false|false|false|C4036459|Contacts|contacts
Event|Event|History of Present Illness|1082,1086|false|false|false|||quit
Event|Event|History of Present Illness|1087,1094|false|false|false|||smoking
Finding|Idea or Concept|History of Present Illness|1111,1116|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|1111,1116|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Gene or Genome|History of Present Illness|1117,1120|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|1127,1134|false|false|false|||reports
Event|Event|History of Present Illness|1138,1145|false|false|false|||episode
Anatomy|Body Location or Region|History of Present Illness|1149,1154|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1149,1154|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1149,1159|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1149,1159|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1155,1159|false|false|false|C2598155||pain
Event|Event|History of Present Illness|1155,1159|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1155,1159|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1155,1159|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1183,1190|false|false|false|||sitting
Event|Event|History of Present Illness|1213,1221|false|false|false|||resolved
Event|Event|History of Present Illness|1244,1250|false|false|false|||denies
Event|Event|History of Present Illness|1251,1256|false|false|false|||fever
Finding|Finding|History of Present Illness|1251,1256|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1251,1256|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|History of Present Illness|1257,1263|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1257,1263|true|false|false|C0085593|Chills|chills
Anatomy|Body Location or Region|History of Present Illness|1265,1274|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1265,1279|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1275,1279|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1275,1279|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1275,1279|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1275,1279|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1281,1287|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|1281,1287|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1281,1287|false|false|false|C0027497|Nausea|nausea
Finding|Sign or Symptom|History of Present Illness|1281,1296|true|false|false|C0027498|Nausea and vomiting|nausea/vomiting
Event|Event|History of Present Illness|1288,1296|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1288,1296|true|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|1299,1311|false|false|false|||palpitations
Finding|Finding|History of Present Illness|1299,1311|false|false|false|C0030252|Palpitations|palpitations
Event|Event|History of Present Illness|1317,1328|false|false|false|||diaphoresis
Finding|Finding|History of Present Illness|1317,1328|false|false|false|C0700590|Increased sweating|diaphoresis
Event|Event|History of Present Illness|1350,1358|false|false|false|||admitted
Event|Event|History of Present Illness|1379,1386|false|false|false|||dyspnea
Finding|Finding|History of Present Illness|1379,1386|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|History of Present Illness|1379,1386|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|History of Present Illness|1397,1404|false|false|false|||thought
Disorder|Neoplastic Process|History of Present Illness|1411,1420|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|History of Present Illness|1411,1420|false|false|false|||secondary
Finding|Functional Concept|History of Present Illness|1411,1420|false|false|false|C1522484|metastatic qualifier|secondary
Drug|Organic Chemical|History of Present Illness|1424,1431|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|History of Present Illness|1424,1431|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|History of Present Illness|1432,1437|false|false|false|||taper
Procedure|Health Care Activity|History of Present Illness|1432,1437|false|false|false|C0441640||taper
Disorder|Disease or Syndrome|History of Present Illness|1449,1453|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|1449,1453|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|1449,1453|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|1449,1453|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|1455,1467|false|false|false|||exacerbation
Finding|Finding|History of Present Illness|1455,1467|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1475,1484|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|History of Present Illness|1475,1484|false|false|false|C1179435|Protein Component|component
Event|Event|History of Present Illness|1475,1484|false|false|false|||component
Finding|Conceptual Entity|History of Present Illness|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|History of Present Illness|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|History of Present Illness|1475,1484|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1488,1495|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|History of Present Illness|1488,1495|false|false|false|||anxiety
Finding|Sign or Symptom|History of Present Illness|1488,1495|false|false|false|C0860603|Anxiety symptoms|anxiety
Finding|Intellectual Product|History of Present Illness|1504,1509|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Disorder|Disease or Syndrome|History of Present Illness|1510,1514|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|1510,1514|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|1510,1514|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|1510,1514|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|History of Present Illness|1516,1528|false|false|false|||exacerbation
Finding|Finding|History of Present Illness|1516,1528|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|History of Present Illness|1538,1545|false|false|false|||treated
Drug|Organic Chemical|History of Present Illness|1551,1559|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|History of Present Illness|1551,1559|false|false|false|C0038317|Steroids|steroids
Event|Event|History of Present Illness|1551,1559|false|false|false|||steroids
Event|Event|History of Present Illness|1564,1571|false|false|false|||duonebs
Drug|Antibiotic|History of Present Illness|1580,1591|false|false|false|C0003232;C0003237;C3540704;C3540705;C3540706;C3540707;C3540708;C3540709;C3540710|Antibiotic throat preparations;Antibiotics;Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE;Antibiotics for systemic use;Antibiotics, Antitubercular;Antibiotics, Gynecological;Antibiotics, ophthalmologic;Antifungal Antibiotics, Topical;antibiotics, intestinal|antibiotics
Event|Event|History of Present Illness|1580,1591|false|false|false|||antibiotics
Event|Event|History of Present Illness|1603,1605|false|false|false|||CT
Event|Event|History of Present Illness|1611,1617|false|false|false|||showed
Disorder|Disease or Syndrome|History of Present Illness|1618,1627|false|false|false|C0034067|Pulmonary Emphysema|emphysema
Event|Event|History of Present Illness|1618,1627|false|false|false|||emphysema
Finding|Pathologic Function|History of Present Illness|1618,1627|false|false|false|C0013990|Pathological accumulation of air in tissues|emphysema
Event|Event|History of Present Illness|1635,1643|false|false|false|||evidence
Finding|Idea or Concept|History of Present Illness|1635,1643|true|false|false|C3887511|Evidence|evidence
Disorder|Disease or Syndrome|History of Present Illness|1648,1657|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|History of Present Illness|1648,1657|false|false|false|||infection
Finding|Pathologic Function|History of Present Illness|1648,1657|false|false|false|C3714514|Infection|infection
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1671,1680|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|History of Present Illness|1671,1680|false|false|false|C2707265||Pulmonary
Finding|Finding|History of Present Illness|1671,1680|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|History of Present Illness|1685,1694|false|false|false|||consulted
Event|Event|History of Present Illness|1700,1711|false|false|false|||recommended
Event|Event|History of Present Illness|1712,1722|false|false|false|||increasing
Drug|Organic Chemical|History of Present Illness|1727,1733|false|false|false|C0965130|Advair|Advair
Drug|Pharmacologic Substance|History of Present Illness|1727,1733|false|false|false|C0965130|Advair|Advair
Event|Event|History of Present Illness|1734,1738|false|false|false|||dose
Event|Event|History of Present Illness|1771,1780|false|false|false|||switching
Drug|Organic Chemical|History of Present Illness|1786,1798|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|History of Present Illness|1786,1798|false|false|false|C0039771|theophylline|theophylline
Event|Event|History of Present Illness|1786,1798|false|false|false|||theophylline
Procedure|Laboratory Procedure|History of Present Illness|1786,1798|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|History of Present Illness|1803,1814|false|false|false|C0965618|roflumilast|roflumilast
Drug|Pharmacologic Substance|History of Present Illness|1803,1814|false|false|false|C0965618|roflumilast|roflumilast
Event|Event|History of Present Illness|1803,1814|false|false|false|||roflumilast
Event|Event|History of Present Illness|1819,1829|false|false|false|||initiation
Finding|Functional Concept|History of Present Illness|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|History of Present Illness|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|History of Present Illness|1819,1829|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Idea or Concept|History of Present Illness|1838,1842|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Finding|Organism Function|History of Present Illness|1838,1842|false|false|false|C0233324;C1705313|Term (lexical);Term Birth|term
Drug|Antibiotic|History of Present Illness|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|History of Present Illness|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|History of Present Illness|1843,1855|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|History of Present Illness|1856,1863|false|false|false|||therapy
Finding|Finding|History of Present Illness|1856,1863|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|History of Present Illness|1856,1863|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1856,1863|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|History of Present Illness|1876,1884|false|false|false|||deferred
Finding|Classification|History of Present Illness|1889,1899|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|History of Present Illness|1889,1899|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|History of Present Illness|1900,1906|false|false|false|||follow
Finding|Functional Concept|History of Present Illness|1900,1906|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|History of Present Illness|1900,1906|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|History of Present Illness|1900,1909|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|History of Present Illness|1900,1909|false|false|false|C1522577|follow-up|follow-up
Event|Event|History of Present Illness|1919,1928|false|false|false|||initiated
Drug|Organic Chemical|History of Present Illness|1935,1942|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|History of Present Illness|1935,1942|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|History of Present Illness|1935,1942|false|false|false|||steroid
Event|Event|History of Present Illness|1944,1949|false|false|false|||taper
Drug|Hormone|History of Present Illness|1960,1970|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|History of Present Illness|1960,1970|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|History of Present Illness|1960,1970|false|false|false|C0032952|prednisone|prednisone
Finding|Intellectual Product|History of Present Illness|1989,1993|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Intellectual Product|History of Present Illness|2013,2017|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Classification|History of Present Illness|2030,2040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|History of Present Illness|2030,2040|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|History of Present Illness|2041,2047|false|false|false|||follow
Finding|Functional Concept|History of Present Illness|2041,2047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|History of Present Illness|2041,2047|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Finding|History of Present Illness|2041,2050|false|false|false|C0589120|Follow-up status|follow-up
Procedure|Health Care Activity|History of Present Illness|2041,2050|false|false|false|C1522577|follow-up|follow-up
Finding|Idea or Concept|History of Present Illness|2064,2071|false|false|false|C1555582|Initial (abbreviation)|initial
Drug|Food|History of Present Illness|2072,2077|false|false|false|C1875856|Vital High Nitrogen Enteral Nutrition|vital
Attribute|Clinical Attribute|History of Present Illness|2072,2083|false|false|false|C0488614;C0518766|Vital signs|vital signs
Procedure|Health Care Activity|History of Present Illness|2072,2083|false|false|false|C0150404|Taking vital signs|vital signs
Event|Event|History of Present Illness|2078,2083|false|false|false|||signs
Finding|Finding|History of Present Illness|2078,2083|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|History of Present Illness|2078,2083|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Event|Event|History of Present Illness|2117,2121|false|false|false|||Exam
Finding|Functional Concept|History of Present Illness|2117,2121|false|false|false|C4284036|Exam|Exam
Procedure|Health Care Activity|History of Present Illness|2117,2121|false|false|false|C0582103|Medical Examination|Exam
Event|Event|History of Present Illness|2126,2133|false|false|false|||notable
Finding|Functional Concept|History of Present Illness|2138,2145|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Finding|Intellectual Product|History of Present Illness|2138,2145|false|false|false|C0439801;C3542948|Limited (extensiveness);Limited component (foundation metadata concept)|limited
Drug|Inorganic Chemical|History of Present Illness|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|History of Present Illness|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|History of Present Illness|2146,2149|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|History of Present Illness|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|History of Present Illness|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|History of Present Illness|2146,2149|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|History of Present Illness|2146,2158|false|false|false|C0001868|Air Movements|air movement
Event|Event|History of Present Illness|2150,2158|false|false|false|||movement
Finding|Organism Function|History of Present Illness|2150,2158|false|false|false|C0026649|Movement|movement
Event|Event|History of Present Illness|2164,2172|false|false|false|||wheezing
Finding|Sign or Symptom|History of Present Illness|2164,2172|false|false|false|C0043144|Wheezing|wheezing
Event|Event|History of Present Illness|2187,2191|false|false|false|||Labs
Lab|Laboratory or Test Result|History of Present Illness|2187,2191|false|false|false|C0587081|Laboratory test finding|Labs
Event|Event|History of Present Illness|2197,2204|false|false|false|||notable
Anatomy|Cell|History of Present Illness|2209,2212|false|false|false|C0023516|Leukocytes|WBC
Event|Event|History of Present Illness|2233,2236|false|false|false|||Plt
Procedure|Laboratory Procedure|History of Present Illness|2233,2236|false|false|false|C0201617|Primed lymphocyte test|Plt
Drug|Biologically Active Substance|History of Present Illness|2258,2261|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Drug|Inorganic Chemical|History of Present Illness|2258,2261|false|false|false|C0600137|Blood Urea Nitrogen|BUN
Event|Event|History of Present Illness|2258,2261|false|false|false|||BUN
Procedure|Laboratory Procedure|History of Present Illness|2258,2261|false|false|false|C0005845|Blood urea nitrogen measurement|BUN
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Hormone|History of Present Illness|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Drug|Pharmacologic Substance|History of Present Illness|2283,2286|false|false|false|C0054015;C5442037|NPPB protein, human;nesiritide|BNP
Event|Event|History of Present Illness|2283,2286|false|false|false|||BNP
Finding|Gene or Genome|History of Present Illness|2283,2286|false|false|false|C1417808;C2982014|NPPB gene;NPPB wt Allele|BNP
Procedure|Laboratory Procedure|History of Present Illness|2283,2286|false|false|false|C1095989|Brain natriuretic peptide measurement|BNP
Drug|Organic Chemical|History of Present Illness|2292,2299|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Drug|Pharmacologic Substance|History of Present Illness|2292,2299|false|false|false|C0022924;C0376261|Lactates;lactate|lactate
Event|Event|History of Present Illness|2292,2299|false|false|false|||lactate
Procedure|Laboratory Procedure|History of Present Illness|2292,2299|false|false|false|C0202115|Lactic acid measurement|lactate
Event|Event|History of Present Illness|2306,2309|false|false|false|||VBG
Event|Event|History of Present Illness|2320,2327|false|false|false|||Imaging
Finding|Finding|History of Present Illness|2320,2327|false|false|false|C0740845|Imaging problem|Imaging
Procedure|Diagnostic Procedure|History of Present Illness|2320,2327|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|Imaging
Event|Event|History of Present Illness|2333,2336|false|false|false|||CXR
Procedure|Diagnostic Procedure|History of Present Illness|2333,2336|false|false|false|C0039985|Plain chest X-ray|CXR
Event|Event|History of Present Illness|2337,2343|false|false|false|||showed
Finding|Intellectual Product|History of Present Illness|2344,2348|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|History of Present Illness|2349,2356|false|false|false|||basilar
Event|Event|History of Present Illness|2358,2369|false|false|false|||atelectasis
Finding|Pathologic Function|History of Present Illness|2358,2369|false|false|false|C0004144|Atelectasis|atelectasis
Disorder|Disease or Syndrome|History of Present Illness|2393,2406|true|false|false|C0521530|Lung consolidation|consolidation
Event|Event|History of Present Illness|2393,2406|false|false|false|||consolidation
Finding|Body Substance|History of Present Illness|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|2412,2419|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|History of Present Illness|2443,2453|false|false|false|C0701466|Solu-Medrol|solumedrol
Drug|Pharmacologic Substance|History of Present Illness|2443,2453|false|false|false|C0701466|Solu-Medrol|solumedrol
Event|Event|History of Present Illness|2481,2489|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|2481,2489|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|2481,2489|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|2481,2489|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Activity|History of Present Illness|2502,2509|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|2502,2509|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|2502,2509|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Anatomy|Anatomical Structure|History of Present Illness|2517,2522|false|false|false|C3714591|Floor (anatomic)|floor
Event|Event|History of Present Illness|2528,2535|false|false|false|||reports
Attribute|Clinical Attribute|History of Present Illness|2540,2549|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|2540,2549|false|false|false|||breathing
Finding|Finding|History of Present Illness|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|2540,2549|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|2540,2549|false|false|false|C1160636|respiratory system process|breathing
Event|Event|History of Present Illness|2554,2562|false|false|false|||improved
Event|Event|History of Present Illness|2565,2571|false|false|false|||REVIEW
Finding|Idea or Concept|History of Present Illness|2565,2571|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Intellectual Product|History of Present Illness|2565,2571|false|false|false|C0282443;C1552617|Act Class - review;Review (Publication Type)|REVIEW
Finding|Functional Concept|History of Present Illness|2565,2574|false|false|false|C0699752|Review of|REVIEW OF
Attribute|Clinical Attribute|History of Present Illness|2565,2582|false|false|false|C0488564;C0488565||REVIEW OF SYSTEMS
Procedure|Health Care Activity|History of Present Illness|2565,2582|false|false|false|C0489633|Review of systems (procedure)|REVIEW OF SYSTEMS
Event|Event|History of Present Illness|2575,2582|false|false|false|||SYSTEMS
Finding|Functional Concept|History of Present Illness|2575,2582|false|false|false|C0449913|System|SYSTEMS
Disorder|Disease or Syndrome|History of Present Illness|2588,2591|false|false|false|C0268529|Proline dehydrogenase deficiency|HPI
Event|Event|History of Present Illness|2588,2591|false|false|false|||HPI
Finding|Finding|History of Present Illness|2588,2591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Finding|Molecular Function|History of Present Illness|2588,2591|false|false|false|C0262512;C1323983|History of present illness (finding);allene oxide synthase activity|HPI
Event|Event|History of Present Illness|2593,2599|false|false|false|||Denies
Event|Event|History of Present Illness|2600,2608|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2600,2608|true|false|false|C0018681|Headache|headache
Finding|Functional Concept|History of Present Illness|2610,2616|false|false|false|C0234621|Visual|visual
Finding|Finding|History of Present Illness|2610,2624|true|false|false|C0750280|Visual changes|visual changes
Event|Event|History of Present Illness|2617,2624|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|2617,2624|false|false|false|C0392747|Changing|changes
Disorder|Disease or Syndrome|History of Present Illness|2627,2638|false|false|false|C0031350|Pharyngitis|pharyngitis
Event|Event|History of Present Illness|2627,2638|false|false|false|||pharyngitis
Event|Event|History of Present Illness|2640,2650|false|false|false|||rhinorrhea
Finding|Sign or Symptom|History of Present Illness|2640,2650|false|false|false|C1260880|Rhinorrhea|rhinorrhea
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|2652,2657|false|false|false|C0028429||nasal
Drug|Biomedical or Dental Material|History of Present Illness|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Organic Chemical|History of Present Illness|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Drug|Pharmacologic Substance|History of Present Illness|2652,2657|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|nasal
Finding|Finding|History of Present Illness|2652,2657|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Functional Concept|History of Present Illness|2652,2657|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|nasal
Finding|Sign or Symptom|History of Present Illness|2652,2668|false|false|false|C0027424|Nasal congestion (finding)|nasal congestion
Event|Event|History of Present Illness|2658,2668|false|false|false|||congestion
Finding|Pathologic Function|History of Present Illness|2658,2668|false|false|false|C0700148|Congestion|congestion
Event|Event|History of Present Illness|2670,2676|false|false|false|||fevers
Finding|Sign or Symptom|History of Present Illness|2670,2676|false|false|false|C0015967|Fever|fevers
Event|Event|History of Present Illness|2678,2684|false|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|2678,2684|false|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|2687,2693|false|false|false|||sweats
Finding|Body Substance|History of Present Illness|2687,2693|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Finding|Finding|History of Present Illness|2687,2693|false|false|false|C0038984;C0038990|Sweat;Sweating|sweats
Attribute|Clinical Attribute|History of Present Illness|2695,2701|false|false|false|C0944911||weight
Event|Event|History of Present Illness|2695,2701|false|false|false|||weight
Finding|Finding|History of Present Illness|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2695,2701|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2695,2701|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|2695,2706|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|2695,2706|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|2702,2706|false|false|false|||loss
Finding|Finding|History of Present Illness|2702,2706|false|false|false|C5890125|Loss (adaptation)|loss
Anatomy|Body Location or Region|History of Present Illness|2708,2717|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|2708,2722|false|false|true|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|2718,2722|false|false|true|C2598155||pain
Event|Event|History of Present Illness|2718,2722|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|2718,2722|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|2718,2722|false|false|true|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|2724,2730|false|false|false|C4255480||nausea
Event|Event|History of Present Illness|2724,2730|false|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|2724,2730|false|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|2732,2740|false|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|2732,2740|false|false|false|C0042963|Vomiting|vomiting
Event|Event|History of Present Illness|2742,2750|false|false|false|||diarrhea
Finding|Finding|History of Present Illness|2742,2750|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|2742,2750|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Event|Event|History of Present Illness|2753,2765|false|false|false|||constipation
Finding|Sign or Symptom|History of Present Illness|2753,2765|false|false|false|C0009806|Constipation|constipation
Disorder|Disease or Syndrome|History of Present Illness|2767,2779|false|false|false|C0018932|Hematochezia|hematochezia
Event|Event|History of Present Illness|2767,2779|false|false|false|||hematochezia
Finding|Sign or Symptom|History of Present Illness|2767,2779|false|false|false|C1321898|Blood in stool|hematochezia
Event|Event|History of Present Illness|2781,2788|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2781,2788|false|false|false|C0013428|Dysuria|dysuria
Disorder|Disease or Syndrome|History of Present Illness|2790,2794|false|false|false|C5779629|Eruption of skin (disorder)|rash
Event|Event|History of Present Illness|2790,2794|false|false|false|||rash
Finding|Pathologic Function|History of Present Illness|2790,2794|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Finding|Sign or Symptom|History of Present Illness|2790,2794|false|false|false|C0015230;C0302295;C5779628|Eruptions;Exanthema;Skin rash|rash
Disorder|Disease or Syndrome|History of Present Illness|2796,2808|false|false|false|C0030554|Paresthesia|paresthesias
Event|Event|History of Present Illness|2796,2808|false|false|false|||paresthesias
Event|Event|History of Present Illness|2815,2823|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|2815,2823|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Disorder|Disease or Syndrome|Past Medical History|2851,2855|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2851,2855|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2851,2855|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2851,2855|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Past Medical History|2856,2862|false|false|false|C0004096|Asthma|Asthma
Event|Event|Past Medical History|2856,2862|false|false|false|||Asthma
Event|Event|Past Medical History|2866,2870|false|false|false|||home
Finding|Idea or Concept|Past Medical History|2866,2870|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Past Medical History|2866,2870|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Past Medical History|2866,2870|false|false|false|C1553498|home health encounter|home
Finding|Finding|Past Medical History|2879,2887|false|false|false|C0741302|atypia morphology|Atypical
Finding|Sign or Symptom|Past Medical History|2879,2898|false|false|false|C0262384|Atypical chest pain|Atypical Chest Pain
Anatomy|Body Location or Region|Past Medical History|2888,2893|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|Chest
Finding|Finding|Past Medical History|2888,2893|false|false|false|C0741025|Chest problem|Chest
Attribute|Clinical Attribute|Past Medical History|2888,2898|false|false|false|C2926613||Chest Pain
Finding|Sign or Symptom|Past Medical History|2888,2898|false|false|false|C0008031|Chest Pain|Chest Pain
Attribute|Clinical Attribute|Past Medical History|2894,2898|false|true|false|C2598155||Pain
Event|Event|Past Medical History|2894,2898|false|false|false|||Pain
Finding|Functional Concept|Past Medical History|2894,2898|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Past Medical History|2894,2898|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Disorder|Disease or Syndrome|Past Medical History|2901,2913|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|2901,2913|false|false|false|||Hypertension
Disorder|Disease or Syndrome|Past Medical History|2916,2930|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Past Medical History|2916,2930|false|false|false|||Hyperlipidemia
Finding|Finding|Past Medical History|2916,2930|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|2951,2957|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Past Medical History|2951,2970|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2951,2970|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Past Medical History|2951,2970|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Past Medical History|2958,2970|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Past Medical History|2958,2970|false|false|false|||Fibrillation
Drug|Organic Chemical|Past Medical History|2974,2982|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Past Medical History|2974,2982|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2985,2992|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Past Medical History|2985,2992|false|false|false|||Anxiety
Finding|Sign or Symptom|Past Medical History|2985,2992|false|false|false|C0860603|Anxiety symptoms|Anxiety
Anatomy|Body Location or Region|Past Medical History|2995,3003|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|2995,3015|false|false|false|C0263884|Cervical radiculitis|Cervical Radiculitis
Disorder|Disease or Syndrome|Past Medical History|3004,3015|false|false|false|C0034544|Radiculitis|Radiculitis
Event|Event|Past Medical History|3004,3015|false|false|false|||Radiculitis
Anatomy|Body Location or Region|Past Medical History|3018,3026|false|false|false|C0027530|Neck|Cervical
Disorder|Disease or Syndrome|Past Medical History|3018,3038|false|false|false|C0158241;C1384641|Cervical spondylosis;Cervical spondylosis without myelopathy|Cervical Spondylosis
Disorder|Disease or Syndrome|Past Medical History|3027,3038|false|false|false|C0038019|Spondylosis|Spondylosis
Event|Event|Past Medical History|3027,3038|false|false|false|||Spondylosis
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3041,3049|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3041,3056|false|false|false|C0205042|Coronary artery|Coronary Artery
Disorder|Disease or Syndrome|Past Medical History|3041,3064|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary Artery Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3050,3056|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Anatomy|Body System|Past Medical History|3050,3056|false|false|false|C0003842;C0226004|Arterial system;Arteries|Artery
Disorder|Disease or Syndrome|Past Medical History|3050,3064|false|false|false|C0852949|Arteriopathic disease|Artery Disease
Disorder|Disease or Syndrome|Past Medical History|3057,3064|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|3057,3064|false|false|false|||Disease
Finding|Sign or Symptom|Past Medical History|3067,3075|false|false|false|C0018681|Headache|Headache
Disorder|Disease or Syndrome|Past Medical History|3078,3084|false|false|false|C0019340;C0854331|Herpes simplex dermatitis|Herpes
Disorder|Disease or Syndrome|Past Medical History|3078,3091|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Virus|Past Medical History|3078,3091|false|false|false|C0019360;C0042338|Herpes zoster (disorder);herpesvirus 3, human|Herpes Zoster
Disorder|Disease or Syndrome|Past Medical History|3085,3091|false|false|false|C0019360|Herpes zoster (disorder)|Zoster
Event|Event|Past Medical History|3085,3091|false|false|false|||Zoster
Finding|Pathologic Function|Past Medical History|3094,3105|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI Bleeding
Event|Event|Past Medical History|3097,3105|false|false|false|||Bleeding
Finding|Pathologic Function|Past Medical History|3097,3105|false|false|false|C0019080|Hemorrhage|Bleeding
Disorder|Disease or Syndrome|Past Medical History|3108,3135|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral Vascular Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3119,3127|false|false|false|C0005847|Blood Vessel|Vascular
Disorder|Disease or Syndrome|Past Medical History|3119,3135|false|false|false|C0042373|Vascular Diseases|Vascular Disease
Disorder|Disease or Syndrome|Past Medical History|3128,3135|false|false|false|C0012634|Disease|Disease
Event|Event|Past Medical History|3128,3135|false|false|false|||Disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3150,3155|false|false|false|C0020889|Bone structure of ilium|iliac
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3150,3162|false|false|false|C0850459|iliac stents|iliac stents
Event|Event|Past Medical History|3156,3162|false|false|false|||stents
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3169,3172|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|Past Medical History|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|Past Medical History|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|Past Medical History|3169,3172|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|Past Medical History|3169,3172|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3169,3172|false|false|false|C1292890|Procedure on hip|hip
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3169,3184|false|false|false|C0392806|Prosthetic arthroplasty of hip (procedure)|hip replacement
Event|Event|Past Medical History|3173,3184|false|false|false|||replacement
Finding|Functional Concept|Past Medical History|3173,3184|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|Past Medical History|3173,3184|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|Past Medical History|3173,3184|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|Family Medical History|3223,3229|false|false|false|||Mother
Finding|Idea or Concept|Family Medical History|3223,3229|false|false|false|C1546508|Relationship - Mother|Mother
Disorder|Disease or Syndrome|Family Medical History|3235,3241|false|false|false|C0004096|Asthma|asthma
Event|Event|Family Medical History|3235,3241|false|false|false|||asthma
Disorder|Disease or Syndrome|Family Medical History|3246,3258|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Family Medical History|3246,3258|false|false|false|||hypertension
Finding|Conceptual Entity|Family Medical History|3260,3266|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|3260,3266|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3272,3277|false|false|false|C0009368;C4071907|Abdomen+Pelvis>Colon;Colon structure (body structure)|colon
Disorder|Disease or Syndrome|Family Medical History|3272,3277|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Disorder|Neoplastic Process|Family Medical History|3272,3277|false|false|false|C0009373;C0154061;C0496907|Carcinoma in situ of colon;Colonic Diseases;Neoplasm of uncertain or unknown behavior of colon|colon
Finding|Finding|Family Medical History|3272,3277|false|false|false|C0750873|COLON PROBLEM|colon
Disorder|Neoplastic Process|Family Medical History|3272,3284|false|false|false|C0007102;C0346629;C0699790|Colon Carcinoma;Malignant neoplasm of large intestine;Malignant tumor of colon|colon cancer
Disorder|Neoplastic Process|Family Medical History|3278,3284|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Family Medical History|3278,3284|false|false|false|||cancer
Event|Event|Family Medical History|3287,3294|false|false|false|||Brother
Finding|Conceptual Entity|Family Medical History|3287,3294|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|3287,3294|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Neoplastic Process|Family Medical History|3300,3308|false|false|false|C0023418|leukemia|leukemia
Event|Event|Family Medical History|3300,3308|false|false|false|||leukemia
Procedure|Health Care Activity|General Exam|3328,3337|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3338,3346|false|false|false|||PHYSICAL
Finding|Finding|General Exam|3338,3346|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3338,3346|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3338,3346|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3338,3351|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3338,3351|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|3347,3351|false|false|false|||EXAM
Finding|Functional Concept|General Exam|3347,3351|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3347,3351|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3380,3386|false|false|false|||VITALS
Event|Event|General Exam|3388,3392|false|false|false|||Temp
Finding|Gene or Genome|General Exam|3388,3392|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|3388,3392|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|3399,3401|false|false|false|||HR
Event|Event|General Exam|3442,3449|false|false|false|||GENERAL
Finding|Classification|General Exam|3442,3449|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|3442,3449|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|3457,3465|false|false|false|||speaking
Event|Event|General Exam|3474,3483|false|false|false|||sentences
Finding|Intellectual Product|General Exam|3474,3483|false|false|true|C0876929|Sentence|sentences
Disorder|Disease or Syndrome|General Exam|3485,3488|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3485,3488|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3485,3488|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|3485,3488|false|false|false|||NAD
Finding|Finding|General Exam|3485,3488|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|3490,3497|false|false|false|||resting
Disorder|Disease or Syndrome|General Exam|3501,3504|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|3501,3504|false|false|false|||bed
Finding|Intellectual Product|General Exam|3501,3504|false|false|false|C2346952|Bachelor of Education|bed
Anatomy|Body Location or Region|General Exam|3519,3524|false|false|false|C1512338|HEENT|HEENT
Event|Event|General Exam|3526,3530|false|false|false|||NCAT
Event|Event|General Exam|3532,3537|false|false|false|||PERRL
Finding|Finding|General Exam|3532,3537|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|3539,3543|false|false|false|||EOMI
Anatomy|Body Part, Organ, or Organ Component|General Exam|3545,3551|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3545,3551|false|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3545,3551|false|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3545,3551|false|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3552,3561|false|false|false|||anicteric
Finding|Finding|General Exam|3552,3561|false|false|false|C0205180|Anicteric|anicteric
Event|Event|General Exam|3570,3578|false|false|false|||injected
Anatomy|Body Part, Organ, or Organ Component|General Exam|3581,3584|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3581,3584|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3581,3584|false|false|false|||MMM
Anatomy|Body Location or Region|General Exam|3586,3596|false|false|false|C0521367|Oropharyngeal|Oropharynx
Event|Event|General Exam|3600,3605|false|false|false|||clear
Finding|Idea or Concept|General Exam|3600,3605|false|false|false|C1550016|Remote control command - Clear|clear
Anatomy|Body Location or Region|General Exam|3607,3611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Anatomy|Cell Component|General Exam|3607,3611|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|NECK
Finding|Finding|General Exam|3607,3611|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|NECK
Event|Event|General Exam|3613,3619|false|false|false|||Supple
Finding|Functional Concept|General Exam|3613,3619|false|false|false|C0332254|Supple|Supple
Anatomy|Body Part, Organ, or Organ Component|General Exam|3624,3627|false|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3624,3627|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3624,3627|false|false|false|||LAD
Finding|Gene or Genome|General Exam|3624,3627|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Event|Event|General Exam|3629,3632|false|false|false|||JVP
Finding|Finding|General Exam|3629,3632|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|3637,3648|false|false|false|||appreciated
Event|Event|General Exam|3655,3662|false|false|false|||degrees
Finding|Intellectual Product|General Exam|3655,3662|false|false|false|C0542560|Academic degree|degrees
Anatomy|Body Part, Organ, or Organ Component|General Exam|3664,3671|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|3664,3671|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Event|General Exam|3685,3694|false|false|false|||irregular
Event|Activity|General Exam|3703,3707|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3703,3707|false|false|false|||rate
Finding|Idea or Concept|General Exam|3703,3707|false|false|false|C1549480|Amount type - Rate|rate
Finding|Organ or Tissue Function|General Exam|3713,3721|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|3713,3728|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|General Exam|3722,3728|false|false|false|||murmur
Finding|Finding|General Exam|3722,3728|false|false|false|C0018808|Heart murmur|murmur
Event|Event|General Exam|3738,3742|false|false|false|||RUSB
Event|Event|General Exam|3747,3751|false|false|false|||rubs
Finding|Finding|General Exam|3747,3751|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3755,3762|false|false|false|||gallops
Anatomy|Body Part, Organ, or Organ Component|General Exam|3764,3769|false|false|false|C0024109|Lung|LUNGS
Finding|Organism Function|General Exam|3771,3781|false|false|false|C0231800|Expiration, Respiratory|Expiratory
Finding|Sign or Symptom|General Exam|3771,3789|false|false|false|C0231875|Expiratory wheezing|Expiratory wheezes
Event|Event|General Exam|3782,3789|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3782,3789|false|false|false|C0043144|Wheezing|wheezes
Finding|Intellectual Product|General Exam|3806,3810|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|General Exam|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|3811,3814|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|General Exam|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|3811,3814|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|General Exam|3811,3823|false|false|false|C0001868|Air Movements|air movement
Event|Event|General Exam|3815,3823|false|false|false|||movement
Finding|Organism Function|General Exam|3815,3823|false|false|false|C0026649|Movement|movement
Anatomy|Body Location or Region|General Exam|3825,3832|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|3825,3832|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|3825,3832|false|false|false|||ABDOMEN
Finding|Finding|General Exam|3825,3832|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|3839,3843|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|3839,3843|false|false|false|||soft
Event|Event|General Exam|3845,3854|false|false|false|||nontender
Event|Event|General Exam|3860,3872|false|false|false|||nondistended
Anatomy|Body Part, Organ, or Organ Component|General Exam|3874,3885|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|3887,3891|false|false|false|||Warm
Finding|Finding|General Exam|3887,3891|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3887,3891|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3896,3900|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3901,3909|false|false|false|||perfused
Attribute|Clinical Attribute|General Exam|3914,3919|true|false|false|C1717255||edema
Event|Event|General Exam|3914,3919|false|false|false|||edema
Finding|Pathologic Function|General Exam|3914,3919|true|false|false|C0013604|Edema|edema
Drug|Food|General Exam|3927,3933|false|false|false|C5890763||pulses
Event|Event|General Exam|3927,3933|false|false|false|||pulses
Finding|Physiologic Function|General Exam|3927,3933|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3927,3933|false|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|3949,3959|false|false|false|||NEUROLOGIC
Event|Event|General Exam|3977,3983|false|false|false|||intact
Finding|Finding|General Exam|3977,3983|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|3985,3993|false|false|false|||strength
Finding|Idea or Concept|General Exam|3985,3993|false|false|false|C0808080|Strength (attribute)|strength
Event|Event|General Exam|3998,4007|false|false|false|||sensation
Finding|Finding|General Exam|3998,4007|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3998,4007|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3998,4007|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|4017,4023|false|false|false|||intact
Finding|Finding|General Exam|4017,4023|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Body Substance|General Exam|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4038,4047|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4038,4047|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4048,4056|false|false|false|||PHYSICAL
Finding|Finding|General Exam|4048,4056|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|4048,4056|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|4048,4056|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|4048,4061|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|4048,4061|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|4057,4061|false|false|false|||EXAM
Finding|Functional Concept|General Exam|4057,4061|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|4057,4061|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|4091,4097|false|false|false|||VITALS
Event|Event|General Exam|4151,4158|false|false|false|||GENERAL
Finding|Classification|General Exam|4151,4158|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|4151,4158|false|false|false|C3812897|General medical service|GENERAL
Event|Event|General Exam|4160,4168|false|false|false|||speaking
Event|Event|General Exam|4177,4186|false|false|false|||sentences
Finding|Intellectual Product|General Exam|4177,4186|false|false|false|C0876929|Sentence|sentences
Disorder|Disease or Syndrome|General Exam|4188,4191|false|false|true|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|4188,4191|false|false|true|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|4188,4191|false|false|true|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|4188,4191|false|false|false|||NAD
Finding|Finding|General Exam|4188,4191|false|false|true|C2051415|patient appears in no acute distress (physical finding)|NAD
Event|Event|General Exam|4193,4200|false|false|false|||resting
Disorder|Disease or Syndrome|General Exam|4204,4207|false|false|true|C3159311|BORNHOLM EYE DISEASE|bed
Event|Event|General Exam|4204,4207|false|false|false|||bed
Finding|Intellectual Product|General Exam|4204,4207|false|false|true|C2346952|Bachelor of Education|bed
Anatomy|Body Part, Organ, or Organ Component|General Exam|4222,4229|false|false|false|C0018787|Heart|CARDIAC
Finding|Intellectual Product|General Exam|4222,4229|false|false|false|C1314974|Cardiac attachment|CARDIAC
Event|Activity|General Exam|4243,4247|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|4243,4247|false|false|false|||rate
Finding|Idea or Concept|General Exam|4243,4247|false|false|false|C1549480|Amount type - Rate|rate
Finding|Organ or Tissue Function|General Exam|4253,4261|false|false|false|C0039155|Systole|systolic
Finding|Finding|General Exam|4253,4268|false|false|false|C0232257|Systolic Murmurs|systolic murmur
Event|Event|General Exam|4262,4268|false|false|false|||murmur
Finding|Finding|General Exam|4262,4268|false|false|false|C0018808|Heart murmur|murmur
Anatomy|Body Part, Organ, or Organ Component|General Exam|4281,4286|false|false|false|C0024109|Lung|LUNGS
Finding|Intellectual Product|General Exam|4289,4293|false|false|false|C1547225|Mild Severity of Illness Code|mild
Event|Event|General Exam|4294,4301|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|4294,4301|false|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|4313,4320|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|ABDOMEN
Disorder|Neoplastic Process|General Exam|4313,4320|false|false|false|C0153662|Malignant neoplasm of abdomen|ABDOMEN
Event|Event|General Exam|4313,4320|false|false|false|||ABDOMEN
Finding|Finding|General Exam|4313,4320|false|false|false|C0941288|Abdomen problem|ABDOMEN
Disorder|Disease or Syndrome|General Exam|4327,4331|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Event|Event|General Exam|4327,4331|false|false|false|||soft
Event|Event|General Exam|4333,4342|false|false|false|||nontender
Event|Event|General Exam|4348,4360|false|false|false|||nondistended
Anatomy|Body Part, Organ, or Organ Component|General Exam|4362,4373|false|false|false|C0015385;C0278454|All extremities;Limb structure|EXTREMITIES
Event|Event|General Exam|4375,4379|false|false|false|||Warm
Finding|Finding|General Exam|4375,4379|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|4375,4379|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|4384,4388|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4389,4397|false|false|false|||perfused
Attribute|Clinical Attribute|General Exam|4410,4415|false|false|false|C1717255||edema
Event|Event|General Exam|4410,4415|false|false|false|||edema
Finding|Pathologic Function|General Exam|4410,4415|false|false|false|C0013604|Edema|edema
Event|Event|General Exam|4418,4428|false|false|false|||NEUROLOGIC
Procedure|Health Care Activity|General Exam|4475,4484|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|4485,4489|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4485,4489|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4530,4535|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4530,4535|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4530,4535|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4536,4539|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4544,4547|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4544,4547|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4544,4547|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4553,4556|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4553,4556|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4553,4556|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4553,4556|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4562,4565|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4562,4565|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4571,4574|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4571,4574|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4571,4574|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4571,4574|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4579,4582|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4579,4582|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4579,4582|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4579,4582|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4579,4582|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4579,4582|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|4588,4592|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|4588,4592|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4621,4624|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4641,4646|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4641,4646|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4641,4646|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|4659,4665|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|4671,4676|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|4682,4685|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|4682,4685|false|false|false|||Eos
Finding|Gene or Genome|General Exam|4682,4685|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4786,4791|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4786,4791|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4786,4791|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4786,4799|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4792,4799|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|4792,4799|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|4792,4799|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4792,4799|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|4832,4837|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4832,4837|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4832,4837|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4842,4845|false|false|false|||pO2
Finding|Classification|General Exam|4842,4845|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Finding|Molecular Function|General Exam|4842,4845|false|false|false|C0391840;C4521535|Partial pressure of Oxygen;US Military enlisted E5|pO2
Procedure|Laboratory Procedure|General Exam|4842,4845|false|false|false|C1283004|PO2 measurement|pO2
Lab|Laboratory or Test Result|General Exam|4850,4854|false|false|false|C0391839|Carbon dioxide, partial pressure|pCO2
Procedure|Laboratory Procedure|General Exam|4850,4854|false|false|false|C0201931|Carbon dioxide measurement, partial pressure|pCO2
Anatomy|Body Location or Region|General Exam|4880,4884|false|false|false|C2987514|Anatomical base|Base
Drug|Biomedical or Dental Material|General Exam|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Chemical Viewed Functionally|General Exam|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|4880,4884|false|false|false|C0178499;C1550601;C1704464;C1880279|Base;Dental Base;base - RoleClass;nitrogenous base|Base
Finding|Gene or Genome|General Exam|4880,4884|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Finding|Idea or Concept|General Exam|4880,4884|false|false|false|C1549548;C1705938;C1843354|BPIFA4P gene;Base - General Qualifier;Base - RX Component Type|Base
Disorder|Disease or Syndrome|General Exam|4902,4907|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4902,4907|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4902,4907|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4902,4915|false|false|false|C3824990|lactate in blood (lab test)|BLOOD Lactate
Drug|Organic Chemical|General Exam|4908,4915|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Drug|Pharmacologic Substance|General Exam|4908,4915|false|false|false|C0022924;C0376261|Lactates;lactate|Lactate
Event|Event|General Exam|4908,4915|false|false|false|||Lactate
Procedure|Laboratory Procedure|General Exam|4908,4915|false|false|false|C0202115|Lactic acid measurement|Lactate
Disorder|Disease or Syndrome|General Exam|4932,4937|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4932,4937|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4932,4937|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4938,4944|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Drug|Hormone|General Exam|4938,4944|false|false|false|C5574646|Natriuretic Peptides B, human|proBNP
Disorder|Disease or Syndrome|General Exam|4961,4966|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4961,4966|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4961,4966|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|4982,4989|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|4982,4989|false|false|false|C0947630|Scientific Study|STUDIES
Event|Event|General Exam|5020,5023|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|5020,5023|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|5031,5035|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Finding|Pathologic Function|General Exam|5036,5055|false|false|false|C4049574|Basilar atelectasis|basilar atelectasis
Event|Event|General Exam|5044,5055|false|false|false|||atelectasis
Finding|Pathologic Function|General Exam|5044,5055|false|false|false|C0004144|Atelectasis|atelectasis
Disorder|Disease or Syndrome|General Exam|5080,5093|false|false|false|C0521530|Lung consolidation|consolidation
Event|Event|General Exam|5080,5093|false|false|false|||consolidation
Event|Event|General Exam|5097,5100|false|false|false|||EKG
Finding|Intellectual Product|General Exam|5097,5100|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|5097,5100|false|false|false|C1623258|Electrocardiography|EKG
Anatomy|Body Space or Junction|General Exam|5102,5107|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|Sinus
Disorder|Anatomical Abnormality|General Exam|5102,5107|false|false|false|C0016169|pathologic fistula|Sinus
Drug|Organic Chemical|General Exam|5102,5107|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Drug|Pharmacologic Substance|General Exam|5102,5107|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|Sinus
Finding|Finding|General Exam|5102,5114|false|false|false|C0232201;C2041122|Sinus rhythm|Sinus rhythm
Event|Event|General Exam|5108,5114|false|false|false|||rhythm
Finding|Finding|General Exam|5108,5114|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|5108,5114|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Functional Concept|General Exam|5122,5126|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|5122,5140|false|false|false|C0459156|Left bundle branch structure|left bundle branch
Disorder|Disease or Syndrome|General Exam|5122,5146|false|false|false|C0023211|Left Bundle-Branch Block|left bundle branch block
Finding|Idea or Concept|General Exam|5122,5146|false|false|false|C2828132|Left Bundle Branch Block Artifact|left bundle branch block
Lab|Laboratory or Test Result|General Exam|5122,5146|false|false|false|C0344420||left bundle branch block
Disorder|Disease or Syndrome|General Exam|5127,5146|false|false|false|C0006384;C1879286|Bundle-Branch Block;Hereditary bundle branch system defect|bundle branch block
Drug|Chemical Viewed Structurally|General Exam|5134,5140|false|false|false|C1881507|Macromolecular Branch|branch
Drug|Biomedical or Dental Material|General Exam|5141,5146|false|false|false|C1706085|Block Dosage Form|block
Event|Event|General Exam|5141,5146|false|false|false|||block
Finding|Body Substance|General Exam|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Finding|General Exam|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Functional Concept|General Exam|5141,5146|false|false|false|C0028778;C0332206;C1533157|Blocking;Fixed Block;Obstruction|block
Finding|Intellectual Product|General Exam|5151,5156|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Finding|General Exam|5164,5170|false|false|false|C0429103|T wave feature|T wave
Finding|Finding|General Exam|5164,5178|false|false|false|C5780423|T wave changes|T wave changes
Finding|Gene or Genome|General Exam|5166,5170|false|false|false|C1421479|WASF1 gene|wave
Phenomenon|Natural Phenomenon or Process|General Exam|5166,5170|false|false|false|C0678544||wave
Event|Event|General Exam|5171,5178|false|false|false|||changes
Finding|Functional Concept|General Exam|5171,5178|false|false|false|C0392747|Changing|changes
Finding|Body Substance|General Exam|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5181,5190|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5181,5190|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|5191,5195|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|5191,5195|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|5236,5241|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5236,5241|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5236,5241|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|5242,5245|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|5253,5256|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|5253,5256|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|5253,5256|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|5262,5265|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|5262,5265|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|5262,5265|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|5262,5265|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|5271,5274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|5271,5274|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|5281,5284|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|5281,5284|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|5281,5284|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|5281,5284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|5281,5284|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|5288,5291|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|5288,5291|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|5288,5291|false|false|false|||MCH
Finding|Gene or Genome|General Exam|5288,5291|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|5288,5291|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|5288,5291|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|5297,5301|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|5297,5301|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|5330,5333|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|5350,5355|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|5350,5355|false|false|false|||BLOOD
Finding|Body Substance|General Exam|5350,5355|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|5350,5363|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|5350,5363|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|5350,5363|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|5356,5363|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|5356,5363|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|5356,5363|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|5356,5363|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|5356,5363|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|5356,5363|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|Hospital Course|5492,5499|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|5492,5499|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|5492,5502|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|5504,5508|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5504,5508|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5504,5508|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5504,5508|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|5512,5516|false|false|false|||home
Finding|Idea or Concept|Hospital Course|5512,5516|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|5512,5516|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|5512,5516|false|false|false|C1553498|home health encounter|home
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|5521,5527|false|false|false|C0018792|Heart Atrium|atrial
Attribute|Clinical Attribute|Hospital Course|5521,5540|false|false|false|C2926591||atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5521,5540|false|false|false|C0004238|Atrial Fibrillation|atrial fibrillation
Lab|Laboratory or Test Result|Hospital Course|5521,5540|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|atrial fibrillation
Disorder|Disease or Syndrome|Hospital Course|5528,5540|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Hospital Course|5528,5540|false|false|false|||fibrillation
Drug|Organic Chemical|Hospital Course|5544,5552|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|5544,5552|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|5544,5552|false|false|false|||apixaban
Disorder|Disease or Syndrome|Hospital Course|5554,5566|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|Hospital Course|5554,5566|false|false|false|||hypertension
Disorder|Disease or Syndrome|Hospital Course|5569,5572|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5569,5572|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5569,5572|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|5569,5572|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|5569,5572|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5569,5572|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|5578,5592|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Hospital Course|5578,5592|false|false|false|||hyperlipidemia
Finding|Finding|Hospital Course|5578,5592|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Event|Event|Hospital Course|5597,5605|false|false|false|||presents
Event|Event|Hospital Course|5611,5620|false|false|false|||shortness
Attribute|Clinical Attribute|Hospital Course|5611,5630|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Hospital Course|5611,5630|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Hospital Course|5624,5630|false|false|false|C0225386|Breath|breath
Drug|Organic Chemical|Hospital Course|5633,5638|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|5633,5638|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|5633,5638|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|5633,5638|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|5644,5652|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5644,5652|false|false|false|C0043144|Wheezing|wheezing
Finding|Idea or Concept|Hospital Course|5661,5664|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|5661,5664|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|5678,5680|false|false|false|||DC
Finding|Idea or Concept|Hospital Course|5688,5696|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Hospital Course|5702,5709|false|false|false|||dyspnea
Finding|Finding|Hospital Course|5702,5709|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|5702,5709|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Event|Event|Hospital Course|5711,5718|false|false|false|||treated
Drug|Biomedical or Dental Material|Hospital Course|5726,5730|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|Hospital Course|5726,5730|false|false|false|||nebs
Drug|Organic Chemical|Hospital Course|5735,5743|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|5735,5743|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|5735,5743|false|false|false|||steroids
Event|Event|Hospital Course|5751,5758|false|false|false|||thought
Disorder|Disease or Syndrome|Hospital Course|5769,5773|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5769,5773|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5769,5773|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5769,5773|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5769,5786|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|5774,5786|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5774,5786|false|false|false|C4086268|Exacerbation|exacerbation
Disorder|Mental or Behavioral Dysfunction|Hospital Course|5792,5799|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|5792,5799|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|5792,5799|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5800,5809|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|5800,5809|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|5800,5809|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|5800,5809|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|Hospital Course|5841,5848|false|false|false|||thought
Finding|Idea or Concept|Hospital Course|5841,5848|false|false|false|C0039869;C4319827|Thought|thought
Finding|Mental Process|Hospital Course|5841,5848|false|false|false|C0039869;C4319827|Thought|thought
Disorder|Disease or Syndrome|Hospital Course|5853,5857|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|5853,5857|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|5853,5857|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|5853,5857|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|5853,5870|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Hospital Course|5858,5870|false|false|false|||exacerbation
Finding|Finding|Hospital Course|5858,5870|false|false|false|C4086268|Exacerbation|exacerbation
Drug|Biomedical or Dental Material|Hospital Course|5881,5885|false|false|false|C1300458|Nebulizer solution|nebs
Event|Event|Hospital Course|5881,5885|false|false|false|||nebs
Drug|Organic Chemical|Hospital Course|5888,5896|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|5888,5896|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|5888,5896|false|false|false|||steroids
Drug|Antibiotic|Hospital Course|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|5898,5910|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|5898,5910|false|false|false|||azithromycin
Event|Event|Hospital Course|5917,5925|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|5917,5925|false|false|false|C0043144|Wheezing|wheezing
Drug|Organic Chemical|Hospital Course|5927,5932|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|5927,5932|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|5927,5932|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|5927,5932|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|5934,5937|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|5934,5937|false|false|false|C0013404|Dyspnea|SOB
Event|Event|Hospital Course|5938,5946|false|false|false|||improved
Finding|Finding|Hospital Course|5938,5946|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|Hospital Course|5938,5946|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Event|Event|Hospital Course|5962,5971|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|5962,5971|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|5976,5984|false|false|false|||titrated
Event|Event|Hospital Course|6000,6004|false|false|false|||well
Finding|Finding|Hospital Course|6000,6004|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Hospital Course|6008,6010|false|false|false|||2L
Drug|Biomedical or Dental Material|Hospital Course|6032,6040|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|6032,6040|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|6032,6040|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|6042,6051|false|false|false|||Evaluated
Event|Event|Hospital Course|6060,6071|false|false|false|||recommended
Event|Event|Hospital Course|6072,6074|false|false|false|||DC
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6079,6088|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6079,6088|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6079,6088|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Hospital Course|6089,6094|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6089,6094|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|6103,6112|false|false|false|||agreeable
Attribute|Clinical Attribute|Hospital Course|6150,6169|false|false|false|C2707305||Shortness of Breath
Finding|Sign or Symptom|Hospital Course|6150,6169|false|false|false|C0013404|Dyspnea|Shortness of Breath
Finding|Body Substance|Hospital Course|6163,6169|false|false|false|C0225386|Breath|Breath
Finding|Body Substance|Hospital Course|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|6171,6178|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|Hospital Course|6184,6191|false|false|false|||history
Finding|Conceptual Entity|Hospital Course|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Hospital Course|6184,6191|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Hospital Course|6184,6194|false|false|false|C0262926|Medical History|history of
Disorder|Disease or Syndrome|Hospital Course|6195,6199|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6195,6199|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6195,6199|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6195,6199|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|6212,6221|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|6212,6221|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|6226,6233|false|false|false|||dyspnea
Finding|Finding|Hospital Course|6226,6233|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Sign or Symptom|Hospital Course|6226,6233|false|false|false|C0013404;C2024878|Dyspnea|dyspnea
Finding|Mental Process|Hospital Course|6241,6248|false|false|false|C0542559|contextual factors|setting
Drug|Organic Chemical|Hospital Course|6252,6259|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Drug|Pharmacologic Substance|Hospital Course|6252,6259|false|false|false|C0038317;C5782153|Steroid [EPC];Steroids|steroid
Event|Event|Hospital Course|6260,6265|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|6260,6265|false|false|false|C0441640||taper
Event|Event|Hospital Course|6272,6280|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|6272,6280|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|6272,6280|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|6284,6296|false|false|false|||presentation
Finding|Idea or Concept|Hospital Course|6284,6296|false|false|false|C0449450|Presentation|presentation
Event|Event|Hospital Course|6302,6312|false|false|false|||consistent
Finding|Idea or Concept|Hospital Course|6302,6312|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Hospital Course|6302,6317|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|Hospital Course|6318,6324|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Hospital Course|6318,6324|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Hospital Course|6325,6329|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|6325,6329|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|6325,6329|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|6325,6329|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Finding|Hospital Course|6337,6353|false|false|false|C2089439|diffuse wheezing|diffuse wheezing
Event|Event|Hospital Course|6345,6353|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|6345,6353|false|false|false|C0043144|Wheezing|wheezing
Finding|Intellectual Product|Hospital Course|6358,6362|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Inorganic Chemical|Hospital Course|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|Hospital Course|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|Hospital Course|6363,6366|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|Hospital Course|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|Hospital Course|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|Hospital Course|6363,6366|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|Hospital Course|6363,6375|false|false|false|C0001868|Air Movements|air movement
Event|Event|Hospital Course|6367,6375|false|false|false|||movement
Finding|Organism Function|Hospital Course|6367,6375|false|false|false|C0026649|Movement|movement
Finding|Finding|Hospital Course|6381,6387|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|6381,6387|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|Hospital Course|6396,6408|false|false|false|||exacerbation
Finding|Finding|Hospital Course|6396,6408|false|false|false|C4086268|Exacerbation|exacerbation
Finding|Mental Process|Hospital Course|6416,6423|false|false|false|C0542559|contextual factors|setting
Event|Event|Hospital Course|6429,6437|false|false|false|||decrease
Finding|Finding|Hospital Course|6429,6437|false|false|false|C0392756|Reduced|decrease
Drug|Organic Chemical|Hospital Course|6445,6453|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|6445,6453|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|6445,6453|false|false|false|||steroids
Drug|Amino Acid, Peptide, or Protein|Hospital Course|6476,6485|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|6476,6485|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|6476,6485|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|6476,6485|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Disorder|Mental or Behavioral Dysfunction|Hospital Course|6489,6496|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|6489,6496|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|6489,6496|false|false|false|C0860603|Anxiety symptoms|anxiety
Event|Event|Hospital Course|6521,6530|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|6521,6530|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|6540,6548|false|false|false|||negative
Finding|Classification|Hospital Course|6540,6548|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|6540,6548|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|6540,6548|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|6540,6552|false|false|false|C0205160|Negative|negative for
Disorder|Disease or Syndrome|Hospital Course|6553,6563|false|false|false|C0851162|Infection of musculoskeletal system|infections
Event|Event|Hospital Course|6553,6563|false|false|false|||infections
Finding|Pathologic Function|Hospital Course|6553,6563|false|false|false|C3714514|Infection|infections
Event|Event|Hospital Course|6586,6595|false|false|false|||continued
Finding|Idea or Concept|Hospital Course|6599,6603|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|6599,6603|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|6599,6603|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|6604,6611|false|false|false|C0905678|Spiriva|spiriva
Drug|Pharmacologic Substance|Hospital Course|6604,6611|false|false|false|C0905678|Spiriva|spiriva
Event|Event|Hospital Course|6604,6611|false|false|false|||spiriva
Drug|Organic Chemical|Hospital Course|6613,6625|false|false|false|C0039771|theophylline|theophylline
Drug|Pharmacologic Substance|Hospital Course|6613,6625|false|false|false|C0039771|theophylline|theophylline
Event|Event|Hospital Course|6613,6625|false|false|false|||theophylline
Procedure|Laboratory Procedure|Hospital Course|6613,6625|false|false|false|C0039773|Assay of theophylline|theophylline
Drug|Organic Chemical|Hospital Course|6627,6633|false|false|false|C0965130|Advair|advair
Drug|Pharmacologic Substance|Hospital Course|6627,6633|false|false|false|C0965130|Advair|advair
Event|Event|Hospital Course|6627,6633|false|false|false|||advair
Event|Event|Hospital Course|6643,6650|false|false|false|||started
Event|Event|Hospital Course|6672,6675|false|false|false|||q6h
Drug|Organic Chemical|Hospital Course|6680,6689|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|6680,6689|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|6680,6689|false|false|false|||albuterol
Event|Event|Hospital Course|6694,6697|false|false|false|||prn
Finding|Gene or Genome|Hospital Course|6694,6697|false|false|false|C1422467|CIAO3 gene|prn
Drug|Hormone|Hospital Course|6702,6712|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|6702,6712|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|6702,6712|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|6702,6712|false|false|false|||prednisone
Event|Event|Hospital Course|6718,6725|false|false|false|||started
Event|Event|Hospital Course|6750,6755|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|6750,6755|false|false|false|C0441640||taper
Event|Event|Hospital Course|6770,6775|false|false|false|||given
Drug|Antibiotic|Hospital Course|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Clinical Drug|Hospital Course|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Drug|Organic Chemical|Hospital Course|6777,6789|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|azithromycin
Event|Event|Hospital Course|6777,6789|false|false|false|||azithromycin
Drug|Organic Chemical|Hospital Course|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|6793,6801|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|6793,6801|false|false|false|||complete
Finding|Functional Concept|Hospital Course|6793,6801|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6793,6801|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|6804,6807|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Hospital Course|6804,6807|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|Hospital Course|6824,6835|false|false|false|||improvement
Finding|Conceptual Entity|Hospital Course|6824,6835|false|false|false|C2986411|Improvement|improvement
Event|Event|Hospital Course|6844,6852|false|false|false|||wheezing
Finding|Sign or Symptom|Hospital Course|6844,6852|false|false|false|C0043144|Wheezing|wheezing
Event|Event|Hospital Course|6857,6865|false|false|false|||returned
Drug|Biomedical or Dental Material|Hospital Course|6869,6877|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|6869,6877|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|6869,6877|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|Hospital Course|6881,6892|false|false|false|||requirement
Finding|Functional Concept|Hospital Course|6881,6892|false|false|false|C1514873|Requirement|requirement
Event|Event|Hospital Course|6903,6908|false|false|false|||hours
Event|Event|Hospital Course|6918,6922|false|false|false|||seen
Event|Event|Hospital Course|6934,6938|false|false|false|||felt
Event|Event|Hospital Course|6954,6961|false|false|false|||benefit
Event|Event|Hospital Course|6968,6977|false|false|false|||discharge
Finding|Body Substance|Hospital Course|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6968,6977|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6968,6977|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Hospital Course|6981,6990|false|false|false|||inpatient
Finding|Idea or Concept|Hospital Course|6981,6990|false|false|false|C1548438;C1549404|Patient Class - Inpatient;Referral category - Inpatient|inpatient
Procedure|Health Care Activity|Hospital Course|6981,6990|false|false|false|C1555324|inpatient encounter|inpatient
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6991,7000|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Hospital Course|6991,7000|false|false|false|C2707265||pulmonary
Finding|Finding|Hospital Course|6991,7000|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6991,7015|false|false|false|C0199529|Pulmonary rehabilitation (procedure)|pulmonary rehabilitation
Event|Event|Hospital Course|7001,7015|false|false|false|||rehabilitation
Finding|Finding|Hospital Course|7001,7015|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Finding|Functional Concept|Hospital Course|7001,7015|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7001,7015|false|false|false|C0034991|Rehabilitation therapy|rehabilitation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7001,7023|false|false|false|C0034991|Rehabilitation therapy|rehabilitation program
Drug|Organic Chemical|Hospital Course|7016,7023|false|false|false|C2728259|Program|program
Drug|Pharmacologic Substance|Hospital Course|7016,7023|false|false|false|C2728259|Program|program
Event|Event|Hospital Course|7016,7023|false|false|false|||program
Finding|Conceptual Entity|Hospital Course|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Functional Concept|Hospital Course|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Finding|Intellectual Product|Hospital Course|7016,7023|false|false|false|C0376691;C1709697;C3484370|Program - framework of goals;Programs;Programs - Publication Format|program
Event|Event|Hospital Course|7039,7044|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7039,7044|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Hospital Course|7046,7057|false|false|false|||recommended
Event|Event|Hospital Course|7058,7067|false|false|false|||continued
Finding|Intellectual Product|Hospital Course|7098,7102|false|false|false|C1561540|Transaction counts and value totals - week|week
Event|Event|Hospital Course|7113,7118|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|7113,7118|false|false|false|C0441640||taper
Event|Event|Hospital Course|7150,7158|false|false|false|||consider
Finding|Idea or Concept|Hospital Course|7150,7158|false|false|false|C0750591|consider|consider
Drug|Organic Chemical|Hospital Course|7168,7175|false|false|false|C0591139|Bactrim|bactrim
Drug|Pharmacologic Substance|Hospital Course|7168,7175|false|false|false|C0591139|Bactrim|bactrim
Event|Event|Hospital Course|7176,7179|false|false|false|||ppx
Finding|Gene or Genome|Hospital Course|7176,7179|false|false|false|C1418850|PPP4C gene|ppx
Finding|Finding|Hospital Course|7185,7193|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|Hospital Course|7185,7193|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Drug|Pharmacologic Substance|Hospital Course|7194,7202|false|false|false|C0720099|Duration brand of oxymetazoline|duration
Event|Event|Hospital Course|7194,7202|false|false|false|||duration
Drug|Organic Chemical|Hospital Course|7206,7214|false|false|false|C0038317|Steroids|steroids
Drug|Pharmacologic Substance|Hospital Course|7206,7214|false|false|false|C0038317|Steroids|steroids
Event|Event|Hospital Course|7206,7214|false|false|false|||steroids
Event|Event|Hospital Course|7219,7225|false|false|false|||unable
Finding|Finding|Hospital Course|7219,7225|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|7229,7233|false|false|false|||wean
Event|Event|Hospital Course|7263,7264|false|false|false|||f
Event|Event|Hospital Course|7270,7280|false|false|false|||outpatient
Finding|Classification|Hospital Course|7270,7280|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7270,7280|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Hospital Course|7287,7291|false|false|false|||pulm
Procedure|Health Care Activity|Hospital Course|7287,7291|false|false|false|C1315068|Pulmonary ventilator management|pulm
Event|Event|Hospital Course|7294,7301|false|false|false|||CHRONIC
Finding|Intellectual Product|Hospital Course|7294,7301|false|false|false|C1547296|Chronic - Admission Level of Care Code|CHRONIC
Procedure|Health Care Activity|Hospital Course|7294,7301|false|false|false|C1555457|Provision of recurring care for chronic illness|CHRONIC
Disorder|Mental or Behavioral Dysfunction|Hospital Course|7332,7339|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|7332,7339|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|7332,7339|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Pharmacologic Substance|Hospital Course|7340,7348|false|false|false|C1950154|Insomnia homeopathic medication|Insomnia
Event|Event|Hospital Course|7340,7348|false|false|false|||Insomnia
Finding|Sign or Symptom|Hospital Course|7340,7348|false|false|false|C0917801|Sleeplessness|Insomnia
Event|Event|Hospital Course|7350,7359|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7360,7364|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7360,7364|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7360,7364|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7365,7374|false|false|false|C0024002|lorazepam|lorazepam
Drug|Pharmacologic Substance|Hospital Course|7365,7374|false|false|false|C0024002|lorazepam|lorazepam
Event|Event|Hospital Course|7365,7374|false|false|false|||lorazepam
Finding|Idea or Concept|Hospital Course|7376,7384|false|false|false|C0750591|consider|Consider
Event|Event|Hospital Course|7395,7399|false|false|false|||SRRI
Event|Event|Hospital Course|7406,7416|false|false|false|||outpatient
Finding|Classification|Hospital Course|7406,7416|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7406,7416|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7421,7427|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Hospital Course|7421,7440|false|false|false|C2926591||Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|7421,7440|false|false|false|C0004238|Atrial Fibrillation|Atrial Fibrillation
Lab|Laboratory or Test Result|Hospital Course|7421,7440|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial Fibrillation
Disorder|Disease or Syndrome|Hospital Course|7428,7440|false|false|false|C0232197|Fibrillation|Fibrillation
Event|Event|Hospital Course|7428,7440|false|false|false|||Fibrillation
Drug|Organic Chemical|Hospital Course|7452,7456|false|false|false|C1601858|Dilt|dilt
Drug|Pharmacologic Substance|Hospital Course|7452,7456|false|false|false|C1601858|Dilt|dilt
Event|Event|Hospital Course|7452,7456|false|false|false|||dilt
Event|Activity|Hospital Course|7461,7465|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|Hospital Course|7461,7465|false|false|false|C1549480|Amount type - Rate|rate
Finding|Functional Concept|Hospital Course|7461,7473|false|false|false|C0489879|rate control|rate control
Drug|Organic Chemical|Hospital Course|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Pharmacologic Substance|Hospital Course|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Drug|Substance|Hospital Course|7466,7473|false|false|false|C0308718;C0728976;C1550141|CONTROL veterinary product;Control brand of phenylpropanolamine;control substance|control
Event|Event|Hospital Course|7466,7473|false|false|false|||control
Finding|Conceptual Entity|Hospital Course|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Functional Concept|Hospital Course|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Finding|Idea or Concept|Hospital Course|7466,7473|false|false|false|C1547100;C1882979;C2587213|Control - Relationship modifier;Control function;Scientific Control|control
Drug|Organic Chemical|Hospital Course|7479,7487|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|7479,7487|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|7479,7487|false|false|false|||apixaban
Event|Event|Hospital Course|7492,7507|false|false|false|||anticoagulation
Finding|Finding|Hospital Course|7492,7507|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|7492,7507|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7492,7507|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Disorder|Disease or Syndrome|Hospital Course|7511,7523|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Hospital Course|7511,7523|false|false|false|||Hypertension
Event|Event|Hospital Course|7525,7534|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7535,7539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7535,7539|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7535,7539|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7540,7545|false|false|false|C0590690|Imdur|imdur
Drug|Pharmacologic Substance|Hospital Course|7540,7545|false|false|false|C0590690|Imdur|imdur
Event|Event|Hospital Course|7540,7545|false|false|false|||imdur
Drug|Organic Chemical|Hospital Course|7547,7566|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|7547,7566|false|false|false|C0020261|hydrochlorothiazide|hydrochlorothiazide
Event|Event|Hospital Course|7547,7566|false|false|false|||hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|7573,7582|false|false|false|C0012373|diltiazem|diltiazem
Drug|Pharmacologic Substance|Hospital Course|7573,7582|false|false|false|C0012373|diltiazem|diltiazem
Event|Event|Hospital Course|7573,7582|false|false|false|||diltiazem
Disorder|Disease or Syndrome|Hospital Course|7586,7589|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7586,7589|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7586,7589|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|7586,7589|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|7586,7589|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7586,7589|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7591,7598|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|Hospital Course|7591,7598|false|false|false|C1314974|Cardiac attachment|Cardiac
Disorder|Injury or Poisoning|Hospital Course|7591,7614|false|false|false|C0261588|Cardiac catheterisation as the cause of abnormal reaction of the patient, or of later complication, without mention of misadventure at the time of the procedure|Cardiac catheterization
Finding|Intellectual Product|Hospital Course|7591,7614|false|false|false|C1547981|Diagnostic Service Section ID - Cardiac Catheterization|Cardiac catheterization
Procedure|Diagnostic Procedure|Hospital Course|7591,7614|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Procedure|Health Care Activity|Hospital Course|7591,7614|false|false|false|C0018795;C1548828|Cardiac Catheterization Procedures;Consent Type - Cardiac Catheterization|Cardiac catheterization
Event|Event|Hospital Course|7599,7614|false|false|false|||catheterization
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7599,7614|false|false|false|C0007430|Catheterization|catheterization
Event|Event|Hospital Course|7630,7638|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|7630,7638|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|7630,7641|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Idea or Concept|Hospital Course|7643,7654|false|false|false|C0750502|Significant|significant
Event|Event|Hospital Course|7655,7663|false|false|false|||stenosis
Finding|Pathologic Function|Hospital Course|7655,7663|false|false|false|C1261287|Stenosis|stenosis
Event|Event|Hospital Course|7667,7677|false|false|false|||coronaries
Event|Event|Hospital Course|7679,7683|false|false|false|||ECHO
Procedure|Health Care Activity|Hospital Course|7679,7683|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7679,7683|false|false|false|C0058928;C5575284|ECHO protocol;Extension for Community Healthcare Outcomes|ECHO
Attribute|Clinical Attribute|Hospital Course|7732,7743|false|false|false|C1980023|Wall motion|wall motion
Phenomenon|Natural Phenomenon or Process|Hospital Course|7737,7743|false|false|false|C0026597|Motion|motion
Disorder|Congenital Abnormality|Hospital Course|7744,7757|false|false|false|C0000768|Congenital Abnormality|abnormalities
Event|Event|Hospital Course|7744,7757|false|false|false|||abnormalities
Finding|Functional Concept|Hospital Course|7744,7757|false|false|false|C0000769|teratologic|abnormalities
Event|Event|Hospital Course|7760,7769|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7770,7774|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7770,7774|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7770,7774|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|7775,7782|false|false|false|C0004057|aspirin|aspirin
Drug|Pharmacologic Substance|Hospital Course|7775,7782|false|false|false|C0004057|aspirin|aspirin
Event|Event|Hospital Course|7775,7782|false|false|false|||aspirin
Drug|Organic Chemical|Hospital Course|7787,7799|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|7787,7799|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|7787,7799|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|Hospital Course|7803,7809|false|false|false|C0002871|Anemia|Anemia
Event|Event|Hospital Course|7803,7809|false|false|false|||Anemia
Event|Event|Hospital Course|7811,7820|false|false|false|||Continued
Finding|Idea or Concept|Hospital Course|7821,7825|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|7821,7825|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|7821,7825|false|false|false|C1553498|home health encounter|home
Drug|Biologically Active Substance|Hospital Course|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Element, Ion, or Isotope|Hospital Course|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Drug|Pharmacologic Substance|Hospital Course|7826,7830|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|iron
Procedure|Laboratory Procedure|Hospital Course|7826,7830|false|false|false|C0337439|Iron measurement|iron
Drug|Inorganic Chemical|Hospital Course|7826,7842|false|false|false|C0721124|Iron Supplement|iron supplements
Drug|Pharmacologic Substance|Hospital Course|7826,7842|false|false|false|C0721124|Iron Supplement|iron supplements
Event|Event|Hospital Course|7831,7842|false|false|false|||supplements
Finding|Idea or Concept|Hospital Course|7845,7857|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|Hospital Course|7858,7864|false|false|false|||ISSUES
Finding|Idea or Concept|Hospital Course|7905,7914|false|false|false|C0549178|Continuous|continued
Disorder|Disease or Syndrome|Hospital Course|7915,7919|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|7915,7919|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|7915,7919|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|7915,7919|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|Hospital Course|7920,7933|false|false|false|||exacerbations
Event|Event|Hospital Course|7935,7944|false|false|false|||recommend
Event|Event|Hospital Course|7945,7954|false|false|false|||finishing
Event|Event|Hospital Course|7959,7965|false|false|false|||course
Drug|Antibiotic|Hospital Course|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Hospital Course|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|7969,7981|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Event|Event|Hospital Course|7969,7981|false|false|false|||Azithromycin
Event|Event|Hospital Course|8005,8014|false|false|false|||Recommend
Finding|Finding|Hospital Course|8015,8023|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Finding|Functional Concept|Hospital Course|8015,8023|false|false|false|C0231448;C5781021|Extended (finding);Extension|extended
Drug|Hormone|Hospital Course|8024,8034|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|8024,8034|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|8024,8034|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|8035,8040|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|8035,8040|false|false|false|C0441640||taper
Drug|Hormone|Hospital Course|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Drug|Organic Chemical|Hospital Course|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Drug|Pharmacologic Substance|Hospital Course|8058,8068|false|false|false|C0032952|prednisone|Prednisone
Finding|Functional Concept|Hospital Course|8073,8079|false|false|false|C1706059|Finish - dosing instruction imperative|finish
Event|Event|Hospital Course|8101,8106|false|false|false|||taper
Procedure|Health Care Activity|Hospital Course|8101,8106|false|false|false|C0441640||taper
Finding|Idea or Concept|Hospital Course|8147,8150|false|false|false|C1548556|Etc.|etc
Event|Event|Hospital Course|8166,8174|false|false|false|||consider
Disorder|Disease or Syndrome|Hospital Course|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|8175,8178|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|8175,8178|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|8175,8178|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|8175,8178|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|8175,8178|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8175,8190|false|false|false|C0747314|pcp prophylaxis|PCP prophylaxis
Event|Event|Hospital Course|8179,8190|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8179,8190|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|Hospital Course|8203,8209|false|false|false|||unable
Finding|Finding|Hospital Course|8203,8209|false|false|false|C1299582|Unable|unable
Event|Event|Hospital Course|8213,8217|false|false|false|||wean
Finding|Finding|Hospital Course|8213,8217|false|false|false|C0043084|Weaning|wean
Drug|Hormone|Hospital Course|8219,8229|false|false|false|C0032952|prednisone|prednisone
Drug|Organic Chemical|Hospital Course|8219,8229|false|false|false|C0032952|prednisone|prednisone
Drug|Pharmacologic Substance|Hospital Course|8219,8229|false|false|false|C0032952|prednisone|prednisone
Event|Event|Hospital Course|8219,8229|false|false|false|||prednisone
Event|Event|Hospital Course|8264,8267|false|false|false|||SOB
Finding|Sign or Symptom|Hospital Course|8264,8267|false|false|false|C0013404|Dyspnea|SOB
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8280,8287|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|anxiety
Event|Event|Hospital Course|8280,8287|false|false|false|||anxiety
Finding|Sign or Symptom|Hospital Course|8280,8287|false|false|false|C0860603|Anxiety symptoms|anxiety
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8288,8297|false|false|false|C1179435|Protein Component|component
Drug|Biologically Active Substance|Hospital Course|8288,8297|false|false|false|C1179435|Protein Component|component
Event|Event|Hospital Course|8288,8297|false|false|false|||component
Finding|Conceptual Entity|Hospital Course|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Idea or Concept|Hospital Course|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Finding|Intellectual Product|Hospital Course|8288,8297|false|false|false|C1524073;C1548799;C1705248|Component (part);Component, LOINC Axis 1;Specimen Child Role - Component|component
Event|Event|Hospital Course|8303,8310|false|false|false|||benefit
Event|Event|Hospital Course|8317,8325|false|false|false|||starting
Drug|Pharmacologic Substance|Hospital Course|8326,8330|false|false|false|C0360105;C2911696|Selective Serotonin Reuptake Inhibitors;Serotonin Reuptake Inhibitor [EPC]|SSRI
Event|Event|Hospital Course|8326,8330|false|false|false|||SSRI
Finding|Functional Concept|Hospital Course|8331,8345|false|false|false|C0332287|In addition to|in addition to
Event|Event|Hospital Course|8334,8342|false|false|false|||addition
Finding|Functional Concept|Hospital Course|8334,8342|false|false|false|C0332287;C1883712|Add - instruction imperative;In addition to|addition
Finding|Idea or Concept|Hospital Course|8346,8350|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|8346,8350|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|8346,8350|false|false|false|C1553498|home health encounter|home
Event|Event|Hospital Course|8351,8357|false|false|false|||benzos
Event|Event|Hospital Course|8366,8376|false|false|false|||prescribed
Event|Activity|Hospital Course|8380,8387|false|false|false|C3812666|Personal Contact|CONTACT
Event|Event|Hospital Course|8380,8387|false|false|false|||CONTACT
Finding|Functional Concept|Hospital Course|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Idea or Concept|Hospital Course|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Finding|Intellectual Product|Hospital Course|8380,8387|false|false|false|C0332158;C1705415;C3245509|Communication Contact;Contact - HL7 Attribution;Contact with|CONTACT
Phenomenon|Phenomenon or Process|Hospital Course|8380,8387|false|false|false|C0392367|Physical contact|CONTACT
Event|Event|Hospital Course|8394,8398|false|false|false|||Code
Event|Occupational Activity|Hospital Course|8394,8398|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|Hospital Course|8394,8398|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Event|Event|Hospital Course|8401,8405|false|false|false|||CODE
Event|Occupational Activity|Hospital Course|8401,8405|false|false|false|C0009219|Coding|CODE
Finding|Intellectual Product|Hospital Course|8401,8405|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|CODE
Procedure|Health Care Activity|Hospital Course|8401,8412|false|false|false|C0742531|CODE STATUS|CODE STATUS
Attribute|Clinical Attribute|Hospital Course|8406,8412|false|false|false|C5889824||STATUS
Event|Event|Hospital Course|8406,8412|false|false|false|||STATUS
Finding|Idea or Concept|Hospital Course|8406,8412|false|false|false|C1546481|What subject filter - Status|STATUS
Disorder|Disease or Syndrome|Hospital Course|8427,8430|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|Hospital Course|8427,8430|false|false|false|||HCP
Finding|Gene or Genome|Hospital Course|8427,8430|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Procedure|Health Care Activity|Hospital Course|8445,8454|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|8473,8483|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|8473,8483|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|8473,8488|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Hospital Course|8484,8488|false|false|false|||list
Finding|Intellectual Product|Hospital Course|8484,8488|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Hospital Course|8492,8500|false|false|false|||accurate
Drug|Organic Chemical|Hospital Course|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|8505,8513|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Hospital Course|8505,8513|false|false|false|||complete
Finding|Functional Concept|Hospital Course|8505,8513|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|8505,8513|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Hospital Course|8518,8531|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|8518,8531|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|8518,8531|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|8518,8531|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|8546,8549|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8550,8554|false|false|false|C2598155||Pain
Event|Event|Hospital Course|8550,8554|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|8550,8554|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|8550,8554|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|8559,8567|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|8559,8567|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8576,8579|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8576,8579|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8576,8579|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8576,8579|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8576,8579|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8584,8591|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|8584,8591|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|8611,8623|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|8611,8623|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|8641,8650|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|8641,8650|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|8651,8659|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8651,8659|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8660,8667|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8660,8667|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8660,8667|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8660,8667|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8678,8681|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8678,8681|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8678,8681|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8678,8681|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8678,8681|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8686,8694|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|8686,8694|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|8686,8694|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|8686,8701|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|8686,8701|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|8695,8701|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|8695,8701|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|8695,8701|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|8695,8701|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8712,8715|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8712,8715|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8712,8715|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8712,8715|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8712,8715|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|8720,8731|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|8720,8731|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|8735,8740|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|8750,8754|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|8750,8754|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|8750,8754|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8755,8764|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8760,8764|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|8760,8764|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|8765,8768|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8765,8768|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|8765,8768|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|8765,8768|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|8765,8768|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|8773,8780|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|8773,8788|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|8773,8788|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|8781,8788|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|8781,8788|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|8809,8820|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|8809,8820|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|8809,8820|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|8809,8831|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|8809,8831|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|8821,8831|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|Hospital Course|8821,8831|false|false|false|||Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8832,8837|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|8832,8837|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|8832,8837|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|8832,8837|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|8840,8844|false|false|false|||SPRY
Event|Event|Hospital Course|8848,8853|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|8854,8857|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|8858,8867|false|false|false|C1717415||allergies
Event|Event|Hospital Course|8858,8867|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|8858,8867|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|Hospital Course|8873,8892|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|8873,8892|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|8913,8923|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|8913,8923|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|8913,8935|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|8913,8935|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|8924,8935|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|8937,8945|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|8937,8945|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|8946,8953|false|false|false|||Release
Finding|Functional Concept|Hospital Course|8946,8953|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|8946,8953|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8946,8953|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|8976,8987|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|8976,8987|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|8995,9000|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|9010,9014|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|9010,9014|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|9010,9014|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9015,9024|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9020,9024|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|9020,9024|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|9034,9047|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|9034,9047|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|9050,9053|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|9050,9053|false|false|false|||TAB
Drug|Hormone|Hospital Course|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|9068,9078|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|9099,9109|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|9099,9109|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|9131,9143|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|9131,9143|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|9131,9143|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|9131,9143|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|9131,9146|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|9131,9146|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9157,9160|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9157,9160|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9157,9160|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9157,9160|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9157,9160|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9166,9176|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|9166,9176|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|9166,9176|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|9166,9184|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9166,9184|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|9177,9184|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9177,9184|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9177,9184|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|9187,9190|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|9187,9190|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|9187,9190|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|9187,9190|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9187,9190|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|9205,9216|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|9205,9216|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|9205,9216|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|9205,9224|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|9205,9224|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|9217,9224|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|9217,9224|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|9217,9224|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|9225,9228|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|9225,9228|false|false|false|||Neb
Finding|Cell Function|Hospital Course|9225,9228|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|9225,9228|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|9231,9234|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|9231,9234|false|false|false|||NEB
Finding|Cell Function|Hospital Course|9231,9234|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9231,9234|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|9242,9245|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|9246,9254|false|false|false|||Wheezing
Finding|Sign or Symptom|Hospital Course|9246,9254|false|false|false|C0043144|Wheezing|Wheezing
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|9260,9263|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Event|Event|Hospital Course|9260,9263|false|false|false|||cod
Finding|Finding|Hospital Course|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|9260,9263|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|9260,9273|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9264,9269|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|9264,9269|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|9264,9269|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|9264,9269|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|9264,9269|false|false|false|||liver
Finding|Finding|Hospital Course|9264,9269|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|9264,9269|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|9270,9273|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9276,9283|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|9276,9283|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|9276,9283|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|Hospital Course|9285,9289|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9285,9289|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9285,9289|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9285,9289|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9290,9293|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9290,9293|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9290,9293|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9290,9293|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9290,9293|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9299,9309|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|Hospital Course|9299,9309|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|Hospital Course|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|9310,9317|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|Hospital Course|9310,9317|false|false|false|||Vitamin
Drug|Hormone|Hospital Course|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|9310,9319|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|9310,9319|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|9318,9319|false|false|false|||D
Drug|Biologically Active Substance|Hospital Course|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|9321,9328|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|9321,9328|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|9321,9328|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|9321,9328|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|9321,9336|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|9321,9336|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|9329,9336|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|9329,9336|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|9329,9336|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|9329,9336|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|9337,9344|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|9337,9344|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|9337,9347|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|9370,9374|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|9370,9374|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|9370,9374|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|9370,9374|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|9375,9380|false|false|false|||DAILY
Drug|Organic Chemical|Hospital Course|9386,9395|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|9386,9395|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|9386,9395|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|9386,9403|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|9386,9403|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|9396,9403|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|9396,9403|false|false|false|||sulfate
Finding|Functional Concept|Hospital Course|9421,9431|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|9421,9431|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|9432,9435|false|false|false|||Q4H
Drug|Organic Chemical|Hospital Course|9441,9452|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9441,9452|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9441,9463|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|9441,9470|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|9441,9470|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|9453,9463|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|9453,9463|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|9464,9470|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|9483,9486|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|9483,9486|false|false|false|||INH
Finding|Functional Concept|Hospital Course|9483,9486|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9490,9493|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9490,9493|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9490,9493|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9490,9493|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9490,9493|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9499,9508|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|9499,9508|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|9523,9526|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9527,9534|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|9527,9534|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|9527,9534|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Organic Chemical|Hospital Course|9540,9551|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|9540,9551|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|Hospital Course|9566,9569|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|9570,9575|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|9570,9575|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|9570,9575|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|9570,9575|false|false|false|C0010200|Coughing|cough
Event|Event|Hospital Course|9580,9589|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|9580,9589|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|9580,9589|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|9580,9601|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|9590,9601|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|9590,9601|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Hospital Course|9590,9601|false|false|false|||Medications
Finding|Intellectual Product|Hospital Course|9590,9601|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|9606,9619|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|9606,9619|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Event|Event|Hospital Course|9606,9619|false|false|false|||Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|9606,9619|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|9634,9637|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|9638,9642|false|false|false|C2598155||Pain
Event|Event|Hospital Course|9638,9642|false|false|false|||Pain
Finding|Functional Concept|Hospital Course|9638,9642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|9638,9642|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|Hospital Course|9647,9656|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|Hospital Course|9647,9656|false|false|false|C0001927|albuterol|albuterol
Event|Event|Hospital Course|9647,9656|false|false|false|||albuterol
Drug|Organic Chemical|Hospital Course|9647,9664|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|Hospital Course|9647,9664|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|Hospital Course|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|Hospital Course|9657,9664|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|Hospital Course|9657,9664|false|false|false|||sulfate
Finding|Functional Concept|Hospital Course|9682,9692|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|Hospital Course|9682,9692|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|Hospital Course|9693,9696|false|false|false|||Q4H
Drug|Organic Chemical|Hospital Course|9701,9709|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Hospital Course|9701,9709|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9718,9721|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9718,9721|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9718,9721|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9718,9721|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9718,9721|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9726,9733|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|9726,9733|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|9753,9765|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|9753,9765|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|9783,9792|false|false|false|C0012373|diltiazem|Diltiazem
Drug|Pharmacologic Substance|Hospital Course|9783,9792|false|false|false|C0012373|diltiazem|Diltiazem
Finding|Finding|Hospital Course|9793,9801|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|9793,9801|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|9802,9809|false|false|false|||Release
Finding|Functional Concept|Hospital Course|9802,9809|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|9802,9809|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9802,9809|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9820,9823|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9820,9823|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9820,9823|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9820,9823|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9820,9823|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9828,9836|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|9828,9836|false|false|false|C1692318|docusate|Docusate
Event|Event|Hospital Course|9828,9836|false|false|false|||Docusate
Drug|Organic Chemical|Hospital Course|9828,9843|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|9828,9843|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|9837,9843|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Event|Event|Hospital Course|9837,9843|false|false|false|||Sodium
Finding|Physiologic Function|Hospital Course|9837,9843|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|9837,9843|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9854,9857|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9854,9857|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9854,9857|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9854,9857|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9854,9857|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|9862,9873|false|false|false|C0165590|dorzolamide|Dorzolamide
Drug|Pharmacologic Substance|Hospital Course|9862,9873|false|false|false|C0165590|dorzolamide|Dorzolamide
Finding|Functional Concept|Hospital Course|9877,9882|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|9892,9896|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|9892,9896|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|9892,9896|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9897,9906|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9902,9906|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|9902,9906|false|false|false|C5848506||EYES
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9907,9910|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9907,9910|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9907,9910|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|9907,9910|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|9907,9910|false|false|false|C1332410|BID gene|BID
Drug|Element, Ion, or Isotope|Hospital Course|9915,9922|false|false|false|C2346592|Ferrous|Ferrous
Drug|Inorganic Chemical|Hospital Course|9915,9930|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Pharmacologic Substance|Hospital Course|9915,9930|false|false|false|C0060282|ferrous sulfate|Ferrous Sulfate
Drug|Element, Ion, or Isotope|Hospital Course|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Inorganic Chemical|Hospital Course|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Drug|Pharmacologic Substance|Hospital Course|9923,9930|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|Sulfate
Event|Event|Hospital Course|9923,9930|false|false|false|||Sulfate
Drug|Organic Chemical|Hospital Course|9952,9963|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|9952,9963|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|Hospital Course|9952,9963|false|false|false|||Fluticasone
Drug|Organic Chemical|Hospital Course|9952,9974|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|Hospital Course|9952,9974|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|Hospital Course|9964,9974|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9975,9980|false|false|false|C0028429||NASAL
Drug|Biomedical or Dental Material|Hospital Course|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Organic Chemical|Hospital Course|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Drug|Pharmacologic Substance|Hospital Course|9975,9980|false|false|false|C0721966;C1272939|Nasal brand of oxymetazoline;Nasal dosage form|NASAL
Finding|Finding|Hospital Course|9975,9980|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Finding|Functional Concept|Hospital Course|9975,9980|false|false|false|C1522019;C4520890|Nasal (intended site);Nasal Route of Administration|NASAL
Event|Event|Hospital Course|9983,9987|false|false|false|||SPRY
Event|Event|Hospital Course|9991,9996|false|false|false|||DAILY
Finding|Gene or Genome|Hospital Course|9997,10000|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|10001,10010|false|false|false|C1717415||allergies
Event|Event|Hospital Course|10001,10010|false|false|false|||allergies
Finding|Pathologic Function|Hospital Course|10001,10010|false|false|false|C0020517|Hypersensitivity|allergies
Drug|Organic Chemical|Hospital Course|10016,10027|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10016,10027|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|Hospital Course|10016,10038|false|false|false|C0939232|fluticasone / salmeterol|Fluticasone-Salmeterol
Drug|Organic Chemical|Hospital Course|10016,10045|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Pharmacologic Substance|Hospital Course|10016,10045|false|false|false|C4762496|Fluticasone-Salmeterol Diskus|Fluticasone-Salmeterol Diskus
Drug|Organic Chemical|Hospital Course|10028,10038|false|false|false|C0073992|salmeterol|Salmeterol
Drug|Pharmacologic Substance|Hospital Course|10028,10038|false|false|false|C0073992|salmeterol|Salmeterol
Event|Event|Hospital Course|10039,10045|false|false|false|||Diskus
Drug|Biomedical or Dental Material|Hospital Course|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Organic Chemical|Hospital Course|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Drug|Pharmacologic Substance|Hospital Course|10058,10061|false|false|false|C0022209;C0598322|Inhalant dose form;isoniazid|INH
Event|Event|Hospital Course|10058,10061|false|false|false|||INH
Finding|Functional Concept|Hospital Course|10058,10061|false|false|false|C0205535|Inhalation Route of Administration|INH
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10065,10068|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10065,10068|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10065,10068|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10065,10068|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10065,10068|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10074,10085|false|false|false|C0018305|guaifenesin|Guaifenesin
Drug|Pharmacologic Substance|Hospital Course|10074,10085|false|false|false|C0018305|guaifenesin|Guaifenesin
Finding|Gene or Genome|Hospital Course|10100,10103|false|false|false|C1422467|CIAO3 gene|PRN
Drug|Organic Chemical|Hospital Course|10104,10109|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|Hospital Course|10104,10109|false|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|Hospital Course|10104,10109|false|false|false|||cough
Finding|Sign or Symptom|Hospital Course|10104,10109|false|false|false|C0010200|Coughing|cough
Drug|Organic Chemical|Hospital Course|10115,10134|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Pharmacologic Substance|Hospital Course|10115,10134|false|false|false|C0020261|hydrochlorothiazide|Hydrochlorothiazide
Drug|Organic Chemical|Hospital Course|10155,10165|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Pharmacologic Substance|Hospital Course|10155,10165|false|false|false|C0022251|isosorbide|Isosorbide
Drug|Organic Chemical|Hospital Course|10155,10177|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Drug|Pharmacologic Substance|Hospital Course|10155,10177|false|false|false|C0064079|isosorbide mononitrate|Isosorbide Mononitrate
Event|Event|Hospital Course|10166,10177|false|false|false|||Mononitrate
Finding|Finding|Hospital Course|10179,10187|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10179,10187|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Event|Event|Hospital Course|10188,10195|false|false|false|||Release
Finding|Functional Concept|Hospital Course|10188,10195|false|false|false|C0391871;C1283071|Release - action (qualifier value);Released (action)|Release
Procedure|Health Care Activity|Hospital Course|10188,10195|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10188,10195|false|false|false|C0030685;C0680255;C1963578|Discharge (release);Patient Discharge;Release (procedure)|Release
Drug|Organic Chemical|Hospital Course|10218,10229|false|false|false|C0090306|latanoprost|Latanoprost
Drug|Pharmacologic Substance|Hospital Course|10218,10229|false|false|false|C0090306|latanoprost|Latanoprost
Finding|Functional Concept|Hospital Course|10237,10242|false|false|false|C1522230|Ophthalmic Route of Administration|Ophth
Drug|Biomedical or Dental Material|Hospital Course|10252,10256|false|false|false|C0991568|Drops - Drug Form|DROP
Event|Activity|Hospital Course|10252,10256|false|false|false|C1705648|Dropping|DROP
Event|Event|Hospital Course|10252,10256|false|false|false|||DROP
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10257,10266|false|false|false|C0229118|Structure of both eyes|BOTH EYES
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10262,10266|false|false|false|C0015392|Eye|EYES
Attribute|Clinical Attribute|Hospital Course|10262,10266|false|false|false|C5848506||EYES
Drug|Organic Chemical|Hospital Course|10276,10285|false|false|false|C0024002|lorazepam|Lorazepam
Drug|Pharmacologic Substance|Hospital Course|10276,10285|false|false|false|C0024002|lorazepam|Lorazepam
Finding|Gene or Genome|Hospital Course|10300,10303|false|false|false|C1422467|CIAO3 gene|PRN
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10304,10311|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|10304,10311|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|10304,10311|false|false|false|C0860603|Anxiety symptoms|Anxiety
Drug|Organic Chemical|Hospital Course|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|10317,10330|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Event|Event|Hospital Course|10317,10330|false|false|false|||Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|10333,10336|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|Hospital Course|10333,10336|false|false|false|||TAB
Drug|Organic Chemical|Hospital Course|10351,10361|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|10351,10361|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Organic Chemical|Hospital Course|10383,10395|false|false|false|C0039771|theophylline|Theophylline
Drug|Pharmacologic Substance|Hospital Course|10383,10395|false|false|false|C0039771|theophylline|Theophylline
Event|Event|Hospital Course|10383,10395|false|false|false|||Theophylline
Procedure|Laboratory Procedure|Hospital Course|10383,10395|false|false|false|C0039773|Assay of theophylline|Theophylline
Drug|Organic Chemical|Hospital Course|10383,10398|false|false|false|C0939729|Theophylline SR|Theophylline SR
Drug|Pharmacologic Substance|Hospital Course|10383,10398|false|false|false|C0939729|Theophylline SR|Theophylline SR
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10409,10412|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10409,10412|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10409,10412|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10409,10412|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10409,10412|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10418,10428|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|Hospital Course|10418,10428|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|Hospital Course|10418,10428|false|false|false|||Tiotropium
Drug|Organic Chemical|Hospital Course|10418,10436|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|Hospital Course|10418,10436|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|Hospital Course|10429,10436|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|10429,10436|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|10429,10436|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|Hospital Course|10439,10442|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|Hospital Course|10439,10442|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|Hospital Course|10439,10442|false|false|false|||CAP
Finding|Gene or Genome|Hospital Course|10439,10442|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10439,10442|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Organic Chemical|Hospital Course|10457,10467|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Pharmacologic Substance|Hospital Course|10457,10467|false|false|false|C3464797|Calcitrate|Calcitrate
Drug|Organic Chemical|Hospital Course|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|10468,10475|false|false|false|C0042890|Vitamins|Vitamin
Event|Event|Hospital Course|10468,10475|false|false|false|||Vitamin
Drug|Hormone|Hospital Course|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|10468,10477|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|10468,10477|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Event|Event|Hospital Course|10476,10477|false|false|false|||D
Drug|Biologically Active Substance|Hospital Course|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|Hospital Course|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|Hospital Course|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|Hospital Course|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|Hospital Course|10479,10486|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|Hospital Course|10479,10486|false|false|false|||calcium
Finding|Physiologic Function|Hospital Course|10479,10486|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|Hospital Course|10479,10486|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|Hospital Course|10479,10494|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Pharmacologic Substance|Hospital Course|10479,10494|false|false|false|C0108101|calcium citrate|calcium citrate
Drug|Organic Chemical|Hospital Course|10487,10494|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Drug|Pharmacologic Substance|Hospital Course|10487,10494|false|false|false|C0008857;C0376259|Citrates;citrate|citrate
Event|Event|Hospital Course|10487,10494|false|false|false|||citrate
Procedure|Laboratory Procedure|Hospital Course|10487,10494|false|false|false|C0201956|Citrate measurement|citrate
Drug|Organic Chemical|Hospital Course|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Hospital Course|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Hospital Course|10495,10502|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Hospital Course|10495,10502|false|false|false|||vitamin
Drug|Organic Chemical|Hospital Course|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Pharmacologic Substance|Hospital Course|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Drug|Vitamin|Hospital Course|10495,10505|false|false|false|C0008318;C3265062|cholecalciferol;vitamin D3|vitamin D3
Anatomy|Body Space or Junction|Hospital Course|10528,10532|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|10528,10532|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|10528,10532|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|10528,10532|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Hospital Course|10533,10538|false|false|false|||DAILY
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Food|Hospital Course|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Immunologic Factor|Hospital Course|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Drug|Pharmacologic Substance|Hospital Course|10544,10547|false|false|false|C0056632;C0459207;C2702357;C3488428|Cyclophosphamide/Dacarbazine/Vincristine;cod, unspecified preparation;codfish allergenic extract|cod
Event|Event|Hospital Course|10544,10547|false|false|false|||cod
Finding|Finding|Hospital Course|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Gene or Genome|Hospital Course|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Finding|Pathologic Function|Hospital Course|10544,10547|false|false|false|C0007465;C0457523;C1420285;C5444130|Cancerization of Pancreatic Ducts;Cause of Death;Cemento-osseous dysplasia;SNRPB gene|cod
Drug|Food|Hospital Course|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Organic Chemical|Hospital Course|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Drug|Pharmacologic Substance|Hospital Course|10544,10557|false|false|false|C0009213|cod liver oil|cod liver oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10548,10553|false|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Hospital Course|10548,10553|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Hospital Course|10548,10553|false|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Hospital Course|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Hospital Course|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Hospital Course|10548,10553|false|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Hospital Course|10548,10553|false|false|false|||liver
Finding|Finding|Hospital Course|10548,10553|false|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Hospital Course|10548,10553|false|false|false|C0872387|Procedures on liver|liver
Drug|Biomedical or Dental Material|Hospital Course|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Food|Hospital Course|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Organic Chemical|Hospital Course|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Drug|Pharmacologic Substance|Hospital Course|10554,10557|false|false|false|C0028908;C1517288;C1947940;C3541397|Food Oil;Oil Dosage Form;Oils;oil ingredients|oil
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10560,10567|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Anatomy|Cell Component|Hospital Course|10560,10567|false|false|false|C0524463;C1325531|Microbial anatomical capsule structure;Structure of organ capsule|capsule
Drug|Biomedical or Dental Material|Hospital Course|10560,10567|false|false|false|C0006935|capsule (pharmacologic)|capsule
Anatomy|Body Space or Junction|Hospital Course|10569,10573|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Hospital Course|10569,10573|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Hospital Course|10569,10573|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Hospital Course|10569,10573|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10574,10577|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10574,10577|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10574,10577|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10574,10577|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10574,10577|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|10583,10594|false|false|false|C0027235|ipratropium|Ipratropium
Drug|Pharmacologic Substance|Hospital Course|10583,10594|false|false|false|C0027235|ipratropium|Ipratropium
Event|Event|Hospital Course|10583,10594|false|false|false|||Ipratropium
Drug|Organic Chemical|Hospital Course|10583,10602|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Pharmacologic Substance|Hospital Course|10583,10602|false|false|false|C0700580|ipratropium bromide|Ipratropium Bromide
Drug|Inorganic Chemical|Hospital Course|10595,10602|false|false|false|C0006222|Bromides|Bromide
Event|Event|Hospital Course|10595,10602|false|false|false|||Bromide
Procedure|Laboratory Procedure|Hospital Course|10595,10602|false|false|false|C0202341|Bromides measurement|Bromide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biologically Active Substance|Hospital Course|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Drug|Biomedical or Dental Material|Hospital Course|10603,10606|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|Neb
Event|Event|Hospital Course|10603,10606|false|false|false|||Neb
Finding|Cell Function|Hospital Course|10603,10606|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Finding|Gene or Genome|Hospital Course|10603,10606|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|Neb
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biologically Active Substance|Hospital Course|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Drug|Biomedical or Dental Material|Hospital Course|10609,10612|false|false|false|C1300458;C1610937|NEB protein, human;Nebulizer solution|NEB
Event|Event|Hospital Course|10609,10612|false|false|false|||NEB
Finding|Cell Function|Hospital Course|10609,10612|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|10609,10612|false|false|false|C1155733;C1417656|NEB gene;mitotic nuclear membrane disassembly|NEB
Finding|Gene or Genome|Hospital Course|10620,10623|false|false|false|C1422467|CIAO3 gene|PRN
Event|Event|Hospital Course|10624,10632|false|false|false|||Wheezing
Finding|Sign or Symptom|Hospital Course|10624,10632|false|false|false|C0043144|Wheezing|Wheezing
Drug|Hazardous or Poisonous Substance|Hospital Course|10638,10646|false|false|false|C0028040|nicotine|Nicotine
Drug|Organic Chemical|Hospital Course|10638,10646|false|false|false|C0028040|nicotine|Nicotine
Drug|Clinical Drug|Hospital Course|10638,10652|false|false|false|C0358855|Nicotine Transdermal Patch|Nicotine Patch
Drug|Biomedical or Dental Material|Hospital Course|10647,10652|false|false|false|C0445403;C1533128;C1707974|Body tissue patch material;Human patch material;Patch - Extended Release Film|Patch
Event|Event|Hospital Course|10647,10652|false|false|false|||Patch
Finding|Finding|Hospital Course|10647,10652|false|false|false|C0332461|Plaque (lesion)|Patch
Drug|Antibiotic|Hospital Course|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Clinical Drug|Hospital Course|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Organic Chemical|Hospital Course|10672,10684|false|false|false|C0052796;C0812732|INJECTION, AZITHROMYCIN, 500 MG ADMINISTERED;azithromycin|Azithromycin
Drug|Pharmacologic Substance|Hospital Course|10700,10708|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Event|Event|Hospital Course|10700,10708|false|false|false|||Duration
Event|Event|Hospital Course|10726,10730|false|false|false|||take
Drug|Hormone|Hospital Course|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Organic Chemical|Hospital Course|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|10742,10752|false|false|false|C0032952|prednisone|PredniSONE
Drug|Pharmacologic Substance|Hospital Course|10768,10776|false|false|false|C0720099|Duration brand of oxymetazoline|Duration
Procedure|Health Care Activity|Hospital Course|10802,10809|false|false|false|C0441640||Tapered
Event|Event|Hospital Course|10817,10821|false|false|false|||DOWN
Event|Event|Hospital Course|10826,10835|false|false|false|||Discharge
Finding|Body Substance|Hospital Course|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|10826,10835|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|10826,10835|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|10826,10847|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|10826,10847|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|10836,10847|false|false|false|C2926604||Disposition
Event|Event|Hospital Course|10836,10847|false|false|false|||Disposition
Procedure|Health Care Activity|Hospital Course|10836,10847|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|10849,10857|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|10849,10862|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|10858,10862|false|false|false|C1947933|care activity|Care
Event|Event|Hospital Course|10858,10862|false|false|false|||Care
Finding|Finding|Hospital Course|10858,10862|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|10858,10862|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Hospital Course|10865,10873|false|false|false|||Facility
Finding|Intellectual Product|Hospital Course|10865,10873|false|false|false|C4695111|ADMIN.FACILITY|Facility
Attribute|Clinical Attribute|Hospital Course|10885,10894|false|false|false|C0945731||Diagnosis
Event|Event|Hospital Course|10885,10894|false|false|false|||Diagnosis
Finding|Classification|Hospital Course|10885,10894|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|10885,10894|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|10885,10894|false|false|false|C0011900|Diagnosis|Diagnosis
Disorder|Disease or Syndrome|Hospital Course|10905,10909|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Hospital Course|10905,10909|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Hospital Course|10905,10909|false|false|false|||COPD
Finding|Gene or Genome|Hospital Course|10905,10909|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Hospital Course|10905,10922|false|false|false|C0740304|COPD exacerbation|COPD Exacerbation
Event|Event|Hospital Course|10910,10922|false|false|false|||Exacerbation
Finding|Finding|Hospital Course|10910,10922|false|false|false|C4086268|Exacerbation|Exacerbation
Disorder|Neoplastic Process|Hospital Course|10924,10933|false|false|false|C0027627|Neoplasm Metastasis|SECONDARY
Event|Event|Hospital Course|10924,10933|false|false|false|||SECONDARY
Finding|Functional Concept|Hospital Course|10924,10933|false|false|false|C1522484|metastatic qualifier|SECONDARY
Disorder|Disease or Syndrome|Hospital Course|10935,10939|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|Hospital Course|10935,10939|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10940,10947|false|false|false|C0003467;C0003469|Anxiety;Anxiety Disorders|Anxiety
Event|Event|Hospital Course|10940,10947|false|false|false|||Anxiety
Finding|Sign or Symptom|Hospital Course|10940,10947|false|false|false|C0860603|Anxiety symptoms|Anxiety
Disorder|Disease or Syndrome|Hospital Course|10948,10951|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|10948,10951|false|false|false|||HTN
Disorder|Disease or Syndrome|Hospital Course|10952,10955|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10952,10955|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|10952,10955|false|false|false|C1504769|DFFB protein, human|CAD
Event|Event|Hospital Course|10952,10955|false|false|false|||CAD
Finding|Gene or Genome|Hospital Course|10952,10955|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10952,10955|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Mental Process|Discharge Condition|10980,10986|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|10980,10993|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|10980,10993|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|10987,10993|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|10987,10993|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|10995,11000|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|10995,11000|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|11005,11013|false|false|false|||coherent
Finding|Finding|Discharge Condition|11005,11013|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|11015,11020|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|11015,11037|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|11015,11037|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|11024,11037|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|11024,11037|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|11024,11037|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|11039,11044|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|11039,11044|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|11039,11044|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|11039,11044|false|false|false|||Alert
Finding|Finding|Discharge Condition|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|11039,11044|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|11049,11060|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|11049,11060|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|11062,11070|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|11062,11070|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|11062,11070|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|11071,11077|false|false|false|C5889824||Status
Event|Event|Discharge Condition|11071,11077|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|11071,11077|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|11079,11089|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|11079,11089|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|11092,11100|false|false|false|||requires
Event|Event|Discharge Condition|11101,11111|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|11101,11111|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|11115,11118|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|11115,11118|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|11115,11118|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|11115,11118|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|11115,11118|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|11120,11126|false|false|false|||walker
Finding|Gene or Genome|Discharge Instructions|11165,11169|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|11189,11197|false|false|false|||admitted
Event|Event|Discharge Instructions|11215,11224|false|false|false|||developed
Event|Event|Discharge Instructions|11226,11235|false|false|false|||shortness
Attribute|Clinical Attribute|Discharge Instructions|11226,11245|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|Discharge Instructions|11226,11245|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|Discharge Instructions|11239,11245|false|false|false|C0225386|Breath|breath
Event|Event|Discharge Instructions|11250,11258|false|false|false|||wheezing
Finding|Sign or Symptom|Discharge Instructions|11250,11258|false|false|false|C0043144|Wheezing|wheezing
Finding|Finding|Discharge Instructions|11259,11266|false|false|false|C4534363|At home|at home
Event|Event|Discharge Instructions|11262,11266|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|11262,11266|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|11262,11266|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|11262,11266|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|11286,11290|false|false|false|||last
Event|Event|Discharge Instructions|11292,11301|false|false|false|||discharge
Finding|Body Substance|Discharge Instructions|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Discharge Instructions|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Discharge Instructions|11292,11301|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Discharge Instructions|11292,11301|false|false|false|C0030685|Patient Discharge|discharge
Event|Event|Discharge Instructions|11312,11319|false|false|false|||treated
Disorder|Disease or Syndrome|Discharge Instructions|11326,11330|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Discharge Instructions|11326,11330|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Discharge Instructions|11326,11330|false|false|false|||COPD
Finding|Gene or Genome|Discharge Instructions|11326,11330|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|Discharge Instructions|11326,11343|false|false|false|C0740304|COPD exacerbation|COPD exacerbation
Event|Event|Discharge Instructions|11331,11343|false|false|false|||exacerbation
Finding|Finding|Discharge Instructions|11331,11343|false|false|false|C4086268|Exacerbation|exacerbation
Event|Event|Discharge Instructions|11354,11363|false|false|false|||breathing
Event|Event|Discharge Instructions|11376,11382|false|false|false|||better
Finding|Idea or Concept|Discharge Instructions|11376,11382|false|false|false|C1550462|Observation Interpretation - better|better
Event|Event|Discharge Instructions|11388,11396|false|false|false|||physical
Finding|Finding|Discharge Instructions|11388,11396|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Finding|Functional Concept|Discharge Instructions|11388,11396|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|physical
Procedure|Health Care Activity|Discharge Instructions|11388,11396|false|false|false|C0031809|Physical Examination|physical
Event|Event|Discharge Instructions|11408,11417|false|false|false|||evaluated
Event|Event|Discharge Instructions|11427,11438|false|false|false|||recommended
Procedure|Health Care Activity|Discharge Instructions|11455,11465|false|false|false|C1698490|short stay encounter|short stay
Event|Event|Discharge Instructions|11461,11465|false|false|false|||stay
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|11469,11478|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|Discharge Instructions|11469,11478|false|false|false|C2707265||Pulmonary
Finding|Finding|Discharge Instructions|11469,11478|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|Discharge Instructions|11497,11501|false|false|false|||home
Finding|Idea or Concept|Discharge Instructions|11497,11501|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|11497,11501|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|11497,11501|false|false|false|C1553498|home health encounter|home
Event|Event|Discharge Instructions|11505,11512|false|false|false|||improve
Attribute|Clinical Attribute|Discharge Instructions|11518,11527|false|false|false|C5885990||breathing
Event|Event|Discharge Instructions|11518,11527|false|false|false|||breathing
Finding|Finding|Discharge Instructions|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|Discharge Instructions|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|Discharge Instructions|11518,11527|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|Discharge Instructions|11518,11527|false|false|false|C1160636|respiratory system process|breathing
Disorder|Disease or Syndrome|Discharge Instructions|11551,11555|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|11551,11555|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|11551,11555|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Event|Discharge Instructions|11559,11564|false|false|false|||rehab
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|11559,11564|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Discharge Instructions|11569,11573|false|false|false|||send
Event|Event|Discharge Instructions|11578,11589|false|false|false|||condolences
Finding|Classification|Discharge Instructions|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Discharge Instructions|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Discharge Instructions|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Discharge Instructions|11599,11605|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|Discharge Instructions|11621,11625|false|false|false|||loss
Finding|Finding|Discharge Instructions|11621,11625|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|Discharge Instructions|11643,11651|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|11643,11651|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|11643,11651|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|11659,11663|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|11659,11663|false|false|false|||care
Finding|Finding|Discharge Instructions|11659,11663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11659,11663|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|11659,11666|false|false|false|C1555558|care of - AddressPartType|care of
Procedure|Health Care Activity|Discharge Instructions|11689,11697|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|11698,11710|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|11698,11710|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|11698,11710|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

