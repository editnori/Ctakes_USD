CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|true|false||Unit
null|Unit device|Device|true|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|true|false||Unit
null|Unit of Measure|LabModifier|true|false||Unit
null|Unit|LabModifier|true|false||Unit
null|Enzyme Unit|LabModifier|true|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|Augmentin|Drug|false|false||Augmentin
null|Augmentin|Drug|false|false||Augmentinnull|Topamax|Drug|false|false||Topamax
null|Topamax|Drug|false|false||Topamaxnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Ultrasonography guided steroid injection|Procedure|false|false||Ultrasound guided steroid injectionnull|Ultrasonic|Finding|false|false||Ultrasoundnull|Urological ultrasound|Procedure|false|false||Ultrasound
null|Ultrasonography|Procedure|false|false||Ultrasoundnull|ultrasound device|Device|false|false||Ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||Ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||Ultrasoundnull|Injection of steroid|Procedure|false|false||steroid injectionnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|Right hip region structure|Anatomy|false|false||right hipnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Woman|Subject|false|false||woman
null|Human, Female adult|Subject|false|false||womannull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Malignant neoplasm of breast|Disorder|false|false||breast cancer
null|Breast Carcinoma|Disorder|false|false||breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|BRCA1 gene mutation|Disorder|false|false||BRCA1 gene mutationnull|BRCA1 gene|Finding|false|false||BRCA1 genenull|BRCA1 gene (lab test)|Procedure|false|false||BRCA1 genenull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Gene Mutation|Finding|false|false||gene mutation
null|Gene Mutant|Finding|false|false||gene mutationnull|Gross Extranodal Extension|Finding|false|false||gene
null|Genes|Finding|false|false||genenull|Mutation Abnormality|Disorder|false|false||mutationnull|Mutation|Finding|false|false||mutationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|Sleep Apnea Syndromes|Disorder|false|false||sleep apneanull|SLEEP APNEA (device)|Device|false|false||sleep apneanull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Apnea|Finding|false|false||apneanull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Hyperlipidemia|Disorder|false|false||hyperlipidemia
null|Hyperlipoproteinemias|Disorder|false|false||hyperlipidemianull|Serum lipids high (finding)|Finding|false|false||hyperlipidemianull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Syndrome|Disorder|false|false||syndromenull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|FBXW7 wt Allele|Finding|false|false||ago
null|FBXW7 gene|Finding|false|false||agonull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain of lower extremities|Finding|false|false||lower extremity painnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Extremity Pain question|Finding|false|false||extremity pain
null|Pain in limb|Finding|false|false||extremity painnull|Limb structure|Anatomy|false|false||extremitynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Ductal Breast Carcinoma|Disorder|false|false||ductal carcinoma
null|Ductal Carcinoma|Disorder|false|false||ductal carcinomanull|Ductal|Modifier|false|false||ductalnull|Carcinoma|Disorder|false|false||carcinomanull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|sentinel|Drug|false|false||sentinel
null|sentinel|Drug|false|false||sentinelnull|Lymph|Finding|false|false||lymphnull|biopsy characteristics|Finding|false|false||biopsy
null|null|Finding|false|false||biopsynull|Biopsy Procedures on the Pharynx, Adenoids, and Tonsils|Procedure|false|false||biopsy
null|Biopsy|Procedure|false|false||biopsy
null|Consent Type - biopsy|Procedure|false|false||biopsynull|Hematoma|Finding|false|false||hematomanull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Evacuation procedure|Procedure|false|false||evacuationnull|null|Time|false|false||Prior tonull|null|Time|false|false||Priornull|Procedure (set of actions)|Finding|false|false||procedures
null|Methods aspects|Finding|false|false||proceduresnull|Interventional procedure|Procedure|false|false||proceduresnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Pain of lower extremities|Finding|false|false||lower extremity painnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Extremity Pain question|Finding|false|false||extremity pain
null|Pain in limb|Finding|false|false||extremity painnull|Limb structure|Anatomy|false|false||extremitynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Similarity|Modifier|false|false||similarnull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Hematoma|Finding|false|false||hematomanull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Prophylactic treatment|Procedure|false|false||prophylaxisnull|prevention & control|Modifier|false|false||prophylaxisnull|Postoperative hematoma|Finding|false|false||postoperative hematomanull|Postoperative Period|Time|false|false||postoperativenull|Hematoma|Finding|false|false||hematomanull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Extremity Pain question|Finding|true|false||extremity pain
null|Pain in limb|Finding|true|false||extremity painnull|Limb structure|Anatomy|true|false||extremitynull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Instructions for Use of the CPT Codebook - Time|Finding|true|false||time
null|Time (foundation metadata concept)|Finding|true|false||time
null|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|true|false||time
null|Value type - Time|Finding|true|false||time
null|Data types - Time|Finding|true|false||time
null|null|Finding|true|false||timenull|Time|Time|true|false||timenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Severe Extremity Pain|Finding|false|false||severe pain
null|Severe pain|Finding|false|false||severe pain
null|Neck Pain Score 6|Finding|false|false||severe painnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Muscle Cramp|Finding|false|false||crampsnull|Middle|Modifier|false|false||midnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Structure of right thigh|Anatomy|false|false||right thighnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Spasm|Finding|false|false||spasmsnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Paresthesia|Disorder|true|false||tinglingnull|Has tingling sensation|Finding|true|false||tinglingnull|Weakness|Finding|false|false||weakness
null|Asthenia|Finding|false|false||weaknessnull|Side|Modifier|false|false||sidenull|Seen in breast clinic|Finding|false|false||seen in breast clinicnull|Breast clinic|Device|false|false||breast clinicnull|Breast clinic|Entity|false|false||breast clinicnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Further|Modifier|false|false||furthernull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Initially|Time|false|false||initiallynull|Absent pulse|Finding|false|false||pulselessnull|Limb structure|Anatomy|false|false||extremitynull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Structure of right foot|Anatomy|false|false||right footnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Minimal|Modifier|false|false||minimal
null|Mild (qualifier value)|Modifier|false|false||minimal
null|Minimum|Modifier|false|false||minimalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarin
null|warfarin|Drug|true|false||warfarinnull|enoxaparin|Drug|true|false||enoxaparin
null|enoxaparin|Drug|true|false||enoxaparinnull|Fixation of dental bridge|Procedure|true|false||bridgenull|Type of bridge device|Device|true|false||bridgenull|Compression Stockings|Device|false|false||compression stockings
null|Support stockings - garment|Device|false|false||compression stockingsnull|null|Finding|false|false||compression
null|Compressed structure|Finding|false|false||compressionnull|Compression Therapy|Procedure|false|false||compression
null|Data Compression|Procedure|false|false||compressionnull|Compression|Phenomenon|false|false||compressionnull|Stocking (hosiery)|Device|false|false||stockings
null|Socks|Device|false|false||stockingsnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Attempt|Event|false|false||attemptnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Right lower extremity|Anatomy|false|false||Right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Palpable|Modifier|false|false||palpablenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Left lower extremity|Anatomy|false|false||left lower extremitynull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Emotional tenderness|Finding|false|false||tenderness
null|Sore to touch|Finding|false|false||tendernessnull|Palpation|Procedure|false|false||palpationnull|Posterior part of right leg|Anatomy|false|false||right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Emotional tenderness|Finding|false|false||Tenderness
null|Sore to touch|Finding|false|false||Tendernessnull|Palpation|Procedure|false|false||palpationnull|Structure of right thigh|Anatomy|false|false||right thighnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Laboratory test finding|Lab|false|false||Labsnull|chemical aspects|Finding|false|false||Chemnull|Chemical procedure|Procedure|false|false||Chemnull|Science of Chemistry|Subject|false|false||Chemnull|Groups|Finding|false|false||panelnull|Panel Device|Device|false|false||panelnull|null|Modifier|false|false||Unremarkablenull|Complete Blood Count|Procedure|false|false||CBCnull|Nuclear cap binding complex location|Anatomy|false|false||CBCnull|Leukocytes|Anatomy|false|false||WBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Modnull|bacteria aspects|Finding|false|false||bacterianull|Bacteria <walking sticks>|Entity|false|false||bacteria
null|Bacteria|Entity|false|false||bacterianull|Imaging problem|Finding|false|false||Imagingnull|Diagnostic Imaging|Procedure|false|false||Imaging
null|Imaging Techniques|Procedure|false|false||Imagingnull|Imaging Technology|Title|false|false||Imagingnull|Ultrasonic|Finding|false|false||Ultrasoundnull|Urological ultrasound|Procedure|false|false||Ultrasound
null|Ultrasonography|Procedure|false|false||Ultrasoundnull|ultrasound device|Device|false|false||Ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||Ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||Ultrasoundnull|Posterior part of right leg|Anatomy|true|false||Right calfnull|Table Cell Horizontal Align - right|Finding|true|false||Rightnull|Right sided|Modifier|true|false||Right
null|Right|Modifier|true|false||Rightnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|true|false||deepnull|Veins|Anatomy|true|false||venousnull|Venous|Modifier|true|false||venousnull|Thrombosis|Finding|true|false||thrombosisnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower extremity>Lower extremity veins|Anatomy|false|false||lower extremity veins
null|Structure of vein of lower extremity|Anatomy|false|false||lower extremity veinsnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Venous structure of limb|Anatomy|false|false||extremity veinsnull|Limb structure|Anatomy|false|false||extremitynull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|null|Attribute|false|false||CT Lower Extremitynull|Lower Extremity|Anatomy|false|false||Lower Extremitynull|Body Site Modifier - Lower|Anatomy|false|false||Lowernull|Lower (action)|Event|false|false||Lowernull|Lower - spatial qualifier|Modifier|false|false||Lowernull|Extremity Right|Anatomy|false|false||Extremity Rightnull|Limb structure|Anatomy|false|false||Extremitynull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|null|Modifier|false|false||Unremarkablenull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Posterior part of right leg|Anatomy|false|false||right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Runoff|Modifier|false|false||runoffnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Procedure on vein|Procedure|true|false||veinsnull|Veins|Anatomy|true|false||veinsnull|Lower Extremity|Anatomy|true|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Limb structure|Anatomy|true|false||extremitynull|Views for patency|Modifier|true|false||patency
null|Open|Modifier|true|false||patencynull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|More|LabModifier|false|false||morenull|Focal|Modifier|true|false||focalnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Obvious|Modifier|true|false||obviousnull|Abnormality of the musculature|Disorder|true|false||muscular abnormalitynull|Muscle (organ)|Anatomy|true|false||muscularnull|Muscular|Modifier|true|false||muscularnull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|morphine|Drug|false|false||Morphine
null|morphine|Drug|false|false||Morphinenull|acetaminophen|Drug|false|false||APAP
null|acetaminophen|Drug|false|false||APAPnull|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED|Disorder|false|false||APAPnull|Dilaudid|Drug|false|false||Dilaudid
null|Dilaudid|Drug|false|false||Dilaudidnull|Total|Modifier|false|false||totalnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|Level of Care - Surgery|Finding|false|false||Surgery
null|Surgical procedure finding|Finding|false|false||Surgery
null|Surgical aspects|Finding|false|false||Surgerynull|Operative Surgical Procedures|Procedure|false|false||Surgerynull|General surgery specialty|Title|false|false||Surgery
null|Surgery specialty|Title|false|false||Surgerynull|Vascular Surgical Procedures|Procedure|false|false||vascular surgerynull|Vascular surgery specialty|Title|false|false||vascular surgerynull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Consultation|Procedure|false|false||consultnull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Deep Vein Thrombosis|Disorder|false|false||dvt
null|Deep thrombophlebitis|Disorder|false|false||dvtnull|area DVT|Anatomy|false|false||dvtnull|null|Attribute|false|false||dvtnull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Numerous|LabModifier|false|false||multiplenull|Stripping of vein|Procedure|false|false||vein strippingnull|Veins|Anatomy|false|false||veinnull|Stripping (procedure)|Procedure|false|false||strippingnull|Procedure (set of actions)|Finding|false|false||procedures
null|Methods aspects|Finding|false|false||proceduresnull|Interventional procedure|Procedure|false|false||proceduresnull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Pharmaceutical Preparations|Drug|false|false||medicinenull|Medicine|Title|false|false||medicinenull|Demonstrates adequate pain control|Finding|false|false||pain controlnull|Pain control|Procedure|false|false||pain control
null|Pain management (procedure)|Procedure|false|false||pain controlnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Control brand of phenylpropanolamine|Drug|false|false||control
null|CONTROL veterinary product|Drug|false|false||control
null|control substance|Drug|false|false||control
null|Control brand of phenylpropanolamine|Drug|false|false||controlnull|Control - Relationship modifier|Finding|false|false||control
null|Control function|Finding|false|false||control
null|Scientific Control|Finding|false|false||controlnull|Control Groups|Subject|false|false||controlnull|True Control Status|Modifier|false|false||control
null|control aspects|Modifier|false|false||controlnull|Vascular Surgical Procedures|Procedure|false|false||Vascular surgerynull|Vascular surgery specialty|Title|false|false||Vascular surgerynull|Blood Vessel|Anatomy|false|false||Vascularnull|Vascular|Modifier|false|false||Vascularnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Remote control command - Clear|Finding|true|false||clearnull|Clear|Modifier|true|false||clear
null|Transparent (qualitative concept)|Modifier|true|false||clearnull|Blood Vessel|Anatomy|true|false||vascularnull|Vascular|Modifier|true|false||vascularnull|Science of Etiology|Finding|true|false||etiology
null|Etiology aspects|Finding|true|false||etiology
null|Etiology|Finding|true|false||etiologynull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Similarity|Modifier|false|false||similarnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Then - dosing instruction fragment|Finding|true|false||thennull|Then|Time|true|false||thennull|Ultrasonic|Finding|true|false||ultrasoundnull|Urological ultrasound|Procedure|true|false||ultrasound
null|Ultrasonography|Procedure|true|false||ultrasoundnull|ultrasound device|Device|true|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|true|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|true|false||ultrasoundnull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Lower extremity>Toes|Anatomy|false|false||toes
null|Toes|Anatomy|false|false||toesnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Never - AcknowledgementCondition|Time|false|false||never
null|Never (frequency)|Time|false|false||nevernull|Terminology Kind|Finding|true|false||kindnull|null|Modifier|true|false||kindnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Stripping of vein|Procedure|false|false||vein strippingnull|Veins|Anatomy|false|false||veinnull|Stripping (procedure)|Procedure|false|false||strippingnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Chest Pain|Finding|true|false||chest painnull|null|Attribute|true|false||chest painnull|Chest problem|Finding|true|false||chestnull|Chest|Anatomy|true|false||chest
null|Anterior thoracic region|Anatomy|true|false||chestnull|Administration Method - Pain|Finding|true|false||pain
null|Pain|Finding|true|false||painnull|null|Attribute|true|false||painnull|Breath|Finding|true|false||breathnull|Recent|Time|true|false||recentnull|travel|Finding|true|false||travelnull|travel charge|Procedure|true|false||travelnull|Physical trauma|Disorder|true|false||trauma
null|Traumatic injury|Disorder|true|false||trauma
null|Trauma|Disorder|true|false||traumanull|Trauma assessment and care|Procedure|true|false||traumanull|Trauma, nursing specialty|Title|true|false||traumanull|trauma qualifier|Modifier|true|false||traumanull|Leg|Anatomy|true|false||leg
null|Lower Extremity|Anatomy|true|false||legnull|Dyslipidemias|Disorder|false|false||Dyslipidemianull|Varicosity|Disorder|false|false||Varicose veinsnull|Varicose|Modifier|false|false||Varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Ligation|Procedure|false|false||ligationnull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|CENPJ gene|Finding|false|false||CPapnull|Continuous Positive Airway Pressure|Procedure|false|false||CPapnull|recent upper respiratory infection|Finding|false|false||recent URInull|Recent|Time|false|false||recentnull|Upper Respiratory Infections|Disorder|false|false||URInull|Uniform Resource Identifier|Finding|false|false||URI
null|URI1 gene|Finding|false|false||URI
null|URI1 wt Allele|Finding|false|false||URInull|Course|Time|false|false||coursenull|Zithromax|Drug|false|false||Zithromax
null|Zithromax|Drug|false|false||Zithromaxnull|Bilateral|Modifier|false|false||bilateralnull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|ANTICOAGULATION (finding)|Finding|false|false||anticoagulation
null|Anticoagulation function|Finding|false|false||anticoagulation
null|Decreased Coagulation Activity [PE]|Finding|false|false||anticoagulationnull|Anticoagulation Therapy|Procedure|false|false||anticoagulationnull|Last|Modifier|false|false||lastnull|United States Military enlisted E3 (qualifier value)|Finding|false|false||A1Cnull|Hemoglobin A1c measurement|Procedure|false|false||A1Cnull|Cerebral Aneurysm|Disorder|false|false||cerebral aneurysmnull|Cerebral hemisphere structure (body structure)|Anatomy|false|false||cerebral
null|Brain|Anatomy|false|false||cerebralnull|Aneurysm|Finding|false|false||aneurysmnull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Diverticulosis|Disorder|false|false||diverticulosisnull|Colonic Polyps|Disorder|false|false||colon polypsnull|Neoplasm of uncertain or unknown behavior of colon|Disorder|false|false||colon
null|Colonic Diseases|Disorder|false|false||colon
null|Carcinoma in situ of colon|Disorder|false|false||colonnull|COLON PROBLEM|Finding|false|false||colonnull|Colon structure (body structure)|Anatomy|false|false||colon
null|Abdomen+Pelvis>Colon|Anatomy|false|false||colonnull|TUBE,COLON,22FR,RADIOPAQUE RUBBER B#7370|Device|false|false||colonnull|Colon <Coloninae>|Entity|false|false||colonnull|polyps|Disorder|false|false||polypsnull|null|Finding|false|false||polypsnull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Candidiasis, Chronic Mucocutaneous|Disorder|false|false||CMC
null|Capillary malformation (disorder)|Disorder|false|false||CMCnull|MCC protocol|Procedure|false|false||CMCnull|Circulating Melanoma Cell|Anatomy|false|false||CMCnull|Cleveland Multiport Catheter|Device|false|false||CMCnull|Chamic Languages|Entity|false|false||CMCnull|Arthroplasty|Procedure|false|false||joint arthroplastynull|Joint problem|Finding|false|false||jointnull|null|Anatomy|false|false||joint
null|Joints|Anatomy|false|false||joint
null|Articular system|Anatomy|false|false||jointnull|Joint Device|Device|false|false||jointnull|Temporomandibular joint arthroplasty by dentist|Procedure|false|false||arthroplasty
null|Arthroplasty|Procedure|false|false||arthroplasty
null|Reconstruction of joint|Procedure|false|false||arthroplastynull|Repair of musculotendinous cuff of shoulder|Procedure|false|false||rotator cuff repairnull|Rotator Cuff|Anatomy|false|false||rotator cuffnull|null|Device|false|false||rotatornull|Cuffing (morphologic abnormality)|Finding|false|false||cuffnull|Cuff - body part|Anatomy|false|false||cuffnull|Cuff Device|Device|false|false||cuffnull|Repair|Finding|false|false||repair
null|Wound Healing|Finding|false|false||repairnull|Repair - Remedial Action|Procedure|false|false||repair
null|Surgical repair|Procedure|false|false||repairnull|Excision|Procedure|false|false||excision
null|removal technique|Procedure|false|false||excisionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GSC-DT gene|Finding|false|false||digitnull|Digit structure|Anatomy|false|false||digitnull|Digit - number character|LabModifier|false|false||digitnull|Mass of body structure|Finding|false|false||mass
null|Morphology, Attenuation, Size, and Structure Criteria|Finding|false|false||mass
null|null|Finding|false|false||mass
null|FBN1 wt Allele|Finding|false|false||mass
null|FBN1 gene|Finding|false|false||mass
null|Mass of body region|Finding|false|false||massnull|Mass, a measure of quantity of matter|LabModifier|false|false||mass
null|Molecular Mass|LabModifier|false|false||massnull|Calculi|Finding|false|false||stonenull|Malignant neoplasm of pancreatic duct|Disorder|false|false||pancreatic ductnull|Abdomen>Pancreatic duct|Anatomy|false|false||pancreatic duct
null|Pancreatic duct|Anatomy|false|false||pancreatic ductnull|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreatic
null|Pancreatic Hormones|Drug|false|false||pancreaticnull|Pancreas|Anatomy|false|false||pancreaticnull|Duct (organ) structure|Anatomy|false|false||duct
null|canal [body parts]|Anatomy|false|false||ductnull|Duct Device|Device|false|false||ductnull|Exploration procedure|Procedure|false|false||explorationnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Tonsillectomy|Procedure|false|false||tonsillectomynull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Malignant neoplasm of brain|Disorder|false|false||BRAIN CANCER
null|Brain Neoplasms|Disorder|false|false||BRAIN CANCERnull|Brain Diseases|Disorder|false|false||BRAINnull|Head>Brain|Anatomy|false|false||BRAIN
null|Brain|Anatomy|false|false||BRAINnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Platinum-Group Metal|Drug|false|false||PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false||PGM
null|PHOSPHOGLUCOMUTASE|Drug|false|false||PGMnull|phosphoglycerate mutase activity|Finding|false|false||PGMnull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Aunt|Subject|false|false||Auntnull|ovarian neoplasm|Disorder|false|true||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|true||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|Malignant Neoplasms|Disorder|false|true||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|true||CANCERnull|Paternal aunt|Subject|false|false||paternal auntnull|Paternal Relative|Subject|false|false||paternalnull|Paternal (qualifier value)|Modifier|false|false||paternalnull|Aunt|Subject|false|false||auntnull|Endometrial Carcinoma|Disorder|false|false||ENDOMETRIAL CANCER
null|Malignant neoplasm of endometrium|Disorder|false|false||ENDOMETRIAL CANCERnull|Endometrial|Modifier|false|false||ENDOMETRIALnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|STAT5A protein, human|Drug|false|false||MGF
null|IGF1 protein, human|Drug|false|false||MGF
null|IGF1 protein, human|Drug|false|false||MGF
null|STAT5A protein, human|Drug|false|false||MGF
null|Kit Ligand, human|Drug|false|false||MGF
null|Kit Ligand, human|Drug|false|false||MGFnull|STAT5A wt Allele|Finding|false|false||MGF
null|KITLG gene|Finding|false|false||MGF
null|STAT5A gene|Finding|false|false||MGF
null|KITLG wt Allele|Finding|false|false||MGFnull|Malignant neoplasm of prostate|Disorder|false|false||PROSTATE CANCER
null|Prostate carcinoma|Disorder|false|false||PROSTATE CANCERnull|Neoplasm of uncertain or unknown behavior of prostate|Disorder|false|false||PROSTATE
null|Prostatic Diseases|Disorder|false|false||PROSTATE
null|Carcinoma in situ of prostate|Disorder|false|false||PROSTATE
null|Benign neoplasm of prostate|Disorder|false|false||PROSTATEnull|Structure of prostate (body structure)|Anatomy|false|false||PROSTATE
null|Prostate|Anatomy|false|false||PROSTATEnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Malignant neoplasm of kidney|Disorder|false|false||KIDNEY CANCER
null|Renal carcinoma|Disorder|false|false||KIDNEY CANCERnull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false||KIDNEY
null|Benign neoplasm of kidney|Disorder|false|false||KIDNEYnull|Kidney problem|Finding|false|false||KIDNEYnull|examination of kidney|Procedure|false|false||KIDNEY
null|Procedures on Kidney|Procedure|false|false||KIDNEYnull|Kidney|Anatomy|false|false||KIDNEY
null|Both kidneys|Anatomy|false|false||KIDNEYnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Kidney Failure|Disorder|false|false||RENAL FAILUREnull|Urologic Diseases|Disorder|false|false||RENALnull|Kidney|Anatomy|false|false||RENALnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Congestive|Modifier|false|false||CONGESTIVEnull|Malignant neoplasm of heart|Disorder|false|false||HEART
null|benign neoplasm of heart|Disorder|false|false||HEARTnull|HEART PROBLEM|Finding|false|false||HEARTnull|Chest>Heart|Anatomy|false|false||HEART
null|Heart|Anatomy|false|false||HEARTnull|Failure (biologic function)|Finding|false|false||FAILURE
null|Failure|Finding|false|false||FAILURE
null|Personal failure|Finding|false|false||FAILUREnull|Diabetes Mellitus|Disorder|false|false||DIABETES MELLITUSnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||DIABETES
null|Diabetes|Disorder|false|false||DIABETES
null|Diabetes Mellitus|Disorder|false|false||DIABETESnull|Tobacco Use Disorder|Disorder|false|false||TOBACCO ABUSEnull|tobacco leaf allergenic extract|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|Tobacco|Drug|false|false||TOBACCO
null|tobacco leaf allergenic extract|Drug|false|false||TOBACCOnull|Nicotiana tabacum|Entity|false|false||TOBACCOnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Sister - courtesy title|Finding|false|false||Sister
null|Relationship - Sister|Finding|false|false||Sisternull|Sister|Subject|false|false||Sisternull|ovarian neoplasm|Disorder|false|false||OVARIAN CANCER
null|Malignant neoplasm of ovary|Disorder|false|false||OVARIAN CANCERnull|Ovarian|Anatomy|false|false||OVARIANnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|true||age
null|Glycation End Products, Advanced|Drug|false|true||agenull|null|Attribute|false|true||agenull|Age|Subject|false|false||agenull|Brother - courtesy title|Finding|false|false||Brother
null|Relationship - Brother|Finding|false|false||Brothernull|Brothers|Subject|false|false||Brothernull|Throat cancer|Disorder|false|false||THROAT CANCERnull|Throat Homeopathic Medication|Drug|false|false||THROATnull|Specimen Type - Throat|Finding|false|false||THROAT
null|null|Finding|false|false||THROATnull|Throat|Anatomy|false|false||THROAT
null|Anterior portion of neck|Anatomy|false|false||THROAT
null|Pharyngeal structure|Anatomy|false|false||THROATnull|null|Attribute|false|false||CANCER dxnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Glycation End Products, Advanced|Drug|false|false||age
null|Glycation End Products, Advanced|Drug|false|false||agenull|null|Attribute|false|false||agenull|Age|Subject|false|false||agenull|Sister - courtesy title|Finding|false|false||Sister
null|Relationship - Sister|Finding|false|false||Sisternull|Sister|Subject|false|false||Sisternull|BRCA1 gene mutation|Disorder|false|false||BRCA1 MUTATIONnull|BRCA1 protein, human|Drug|false|false||BRCA1
null|BRCA1 protein, human|Drug|false|false||BRCA1null|BRCA1 gene|Finding|false|false||BRCA1null|Mutation Abnormality|Disorder|false|false||MUTATIONnull|Mutation|Finding|false|false||MUTATIONnull|Malignant neoplasm of breast|Disorder|false|true||BREAST CANCER
null|Breast Carcinoma|Disorder|false|true||BREAST CANCERnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||BREASTnull|Breast problem|Finding|false|false||BREASTnull|Procedures on breast|Procedure|false|false||BREASTnull|Breast|Anatomy|false|false||BREASTnull|Malignant Neoplasms|Disorder|false|false||CANCERnull|Specialty Type - cancer|Title|false|false||CANCERnull|Cancer <Cancridae>|Entity|false|false||CANCERnull|Daughter|Subject|false|false||Daughternull|Abnormal cervical smear|Finding|false|false||ABNORMAL PAP SMEARnull|Observation Interpretation - Abnormal|Finding|false|false||ABNORMAL
null|Abnormal|Finding|false|false||ABNORMALnull|Pap smear|Procedure|false|false||PAP SMEAR
null|Papanicolaou Test|Procedure|false|false||PAP SMEARnull|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false||PAP
null|alpha 2-plasmin inhibitor-plasmin complex|Drug|false|false||PAP
null|ACPP protein, human|Drug|false|false||PAP
null|ACPP protein, human|Drug|false|false||PAPnull|null|Finding|false|false||PAP
null|PAPOLA wt Allele|Finding|false|false||PAP
null|PDAP1 gene|Finding|false|false||PAP
null|TUSC2 wt Allele|Finding|false|false||PAP
null|ASAP1 wt Allele|Finding|false|false||PAP
null|ACP3 wt Allele|Finding|false|false||PAP
null|Pulmonary artery pressure|Finding|false|false||PAP
null|TUSC2 gene|Finding|false|false||PAP
null|ASAP2 gene|Finding|false|false||PAP
null|ASAP1 gene|Finding|false|false||PAP
null|REG3A gene|Finding|false|false||PAP
null|PITUITARY ADENOMA PREDISPOSITION|Finding|false|false||PAP
null|PAPOLA gene|Finding|false|false||PAP
null|ACP3 gene|Finding|false|false||PAP
null|REG3A wt Allele|Finding|false|false||PAP
null|MRPS30 gene|Finding|false|false||PAPnull|pars anterior of the paramedian lobule|Anatomy|false|false||PAPnull|Papiamento language|Entity|false|false||PAPnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|SON gene|Finding|false|false||Sonnull|Son (person)|Subject|false|false||Sonnull|Songhay Languages|Entity|false|false||Sonnull|Substance Abuse Problems|Disorder|false|false||SUBSTANCE ABUSE
null|Harmful pattern of substance use|Disorder|false|false||SUBSTANCE ABUSEnull|Substance|Drug|false|false||SUBSTANCEnull|administrative information regarding test substance|Finding|false|false||SUBSTANCEnull|null|Attribute|false|false||SUBSTANCEnull|Substance (attribute)|Modifier|false|false||SUBSTANCEnull|Drug abuse|Disorder|false|false||ABUSEnull|Victim of abuse (finding)|Finding|false|false||ABUSEnull|Abuse|Event|false|false||ABUSEnull|Heroin overdose|Disorder|false|false||heroin overdosenull|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroin
null|heroin|Drug|false|false||heroinnull|Poisoning by heroin|Disorder|false|false||heroinnull|Drug Overdose|Disorder|false|false||overdosenull|Event Qualification - Overdose|Finding|false|false||overdose
null|Overdose|Finding|false|false||overdosenull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|SAT1 protein, human|Drug|false|false||Sat
null|SAT1 protein, human|Drug|false|false||Satnull|College Entrance Examination Board Scholastic Aptitude Test|Finding|false|false||Sat
null|SAT1 wt Allele|Finding|false|false||Sat
null|SAT1 gene|Finding|false|false||Satnull|Santali language|Entity|false|false||Satnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|true|false||Alert
null|Alert brand of caffeine|Drug|true|false||Alertnull|Mentally alert|Finding|true|false||Alert
null|Consciousness clear|Finding|true|false||Alert
null|Alert note|Finding|true|false||Alert
null|Alert|Finding|true|false||Alertnull|null|Attribute|true|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|true|false||HEENTnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|true|false||PERRLnull|Supple neck|Finding|true|false||neck supplenull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|true|false||neck
null|Neck|Anatomy|true|false||necknull|Supple|Finding|true|false||supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Elevated|Modifier|true|false||elevated
null|High|Modifier|true|false||elevatednull|Chest problem|Finding|true|false||Chestnull|Chest|Anatomy|true|false||Chest
null|Anterior thoracic region|Anatomy|true|false||Chestnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Surgical incisions|Procedure|false|false||incisionsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Healed|Finding|false|false||healednull|Axilla|Anatomy|false|false||axillanull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|true|false||rhythm
null|rhythmic process (biological)|Finding|true|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|true|false||Lungsnull|Remote control command - Clear|Finding|true|false||Clearnull|Clear|Modifier|true|false||Clear
null|Transparent (qualitative concept)|Modifier|true|false||Clearnull|Auscultation|Procedure|true|false||auscultationnull|Wheezing|Finding|true|false||wheezesnull|Basilar Rales|Finding|true|false||crackles
null|Rales|Finding|true|false||cracklesnull|Malignant neoplasm of abdomen|Disorder|true|false||Abdomennull|Abdomen problem|Finding|true|false||Abdomennull|Abdomen|Anatomy|true|false||Abdomen
null|Abdominal Cavity|Anatomy|true|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Movement|Finding|false|false||movementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Swelling|Finding|false|false||Swelling
null|Edema|Finding|false|false||Swellingnull|Palpable|Modifier|false|false||Palpablenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Symmetric Relationship|Finding|false|false||symmetric
null|Symmetrical|Finding|false|false||symmetricnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|C1orf210 gene|Finding|false|false||Tempnull|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Procedure|false|false||Tempnull|Temperature|LabModifier|false|false||Tempnull|delivery (history)|Finding|false|false||delivery
null|Transfer Technique|Finding|false|false||delivery
null|null|Finding|false|false||deliverynull|Obstetric Delivery|Procedure|false|false||deliverynull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|Alert brand of caffeine|Drug|true|false||Alert
null|Alert brand of caffeine|Drug|true|false||Alertnull|Mentally alert|Finding|true|false||Alert
null|Consciousness clear|Finding|true|false||Alert
null|Alert note|Finding|true|false||Alert
null|Alert|Finding|true|false||Alertnull|null|Attribute|true|false||Alertnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|true|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|true|false||HEENTnull|Myelofibrosis|Disorder|false|false||MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false||MMMnull|Oropharyngeal|Anatomy|false|false||oropharynxnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Pupil equal round and reacting to light|Finding|true|false||PERRLnull|Supple neck|Finding|true|false||neck supplenull|Passive joint movement of neck (finding)|Finding|true|false||neck
null|Neck problem|Finding|true|false||necknull|dendritic spine neck|Anatomy|true|false||neck
null|Neck|Anatomy|true|false||necknull|Supple|Finding|true|false||supplenull|Jugular venous pressure|Finding|true|false||JVPnull|Elevated|Modifier|true|false||elevated
null|High|Modifier|true|false||elevatednull|Chest problem|Finding|true|false||Chestnull|Chest|Anatomy|true|false||Chest
null|Anterior thoracic region|Anatomy|true|false||Chestnull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Surgical incisions|Procedure|false|false||incisionsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Healed|Finding|false|false||healednull|Axilla|Anatomy|false|false||axillanull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Removal of drain|Procedure|false|false||drain removalnull|Drain - SpecimenType|Drug|false|false||drainnull|Drain Specimen Code|Finding|false|false||drainnull|Drain device|Device|false|false||drainnull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|true|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Malignant neoplasm of abdomen|Disorder|false|false||Abdomennull|Abdomen problem|Finding|false|false||Abdomennull|Abdomen|Anatomy|false|false||Abdomen
null|Abdominal Cavity|Anatomy|false|false||Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false||bowel soundsnull|Intestines|Anatomy|false|false||bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Present|Finding|false|false||present
null|Presentation|Finding|false|false||presentnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Asymmetry (qualifier value)|Modifier|true|false||asymmetricnull|Swelling|Finding|true|false||swelling
null|Edema|Finding|true|false||swellingnull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of trochanteric bursa|Anatomy|false|false||trochanteric bursanull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|Tender|Modifier|false|false||tendernull|Palpation|Procedure|false|false||palpationnull|Right tibia|Anatomy|false|false||right tibianull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Bone structure of tibia|Anatomy|false|false||tibianull|Tibia <Rostellariidae>|Entity|false|false||tibianull|Rupture of Membranes|Finding|false|false||ROM
null|ROM1 gene|Finding|false|false||ROMnull|Range of motion technique (procedure)|Procedure|false|false||ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Knee flexion|Finding|false|false||knee flexionnull|Examination of knee joint|Procedure|false|false||kneenull|Knee region structure|Anatomy|false|false||knee
null|Knee|Anatomy|false|false||knee
null|Lower extremity>Knee|Anatomy|false|false||knee
null|Knee joint|Anatomy|false|false||kneenull|null|Finding|false|false||flexionnull|W flexion|Attribute|false|false||flexionnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Telephone Extension Number|Finding|false|false||extension
null|Extension|Finding|false|false||extensionnull|Palpable|Modifier|false|false||Palpablenull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false||Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false||Skinnull|Skin Specimen Source Code|Finding|false|false||Skin
null|Skin Specimen|Finding|false|false||Skinnull|Skin, Human|Anatomy|false|false||Skin
null|Skin|Anatomy|false|false||Skinnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Lower Extremity|Anatomy|false|false||lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Relational Operator - Equal|Finding|false|false||equalnull|Equal|Modifier|false|false||equalnull|Bilateral|Modifier|false|false||both sidesnull|TNFSF14 protein, human|Drug|false|false||light
null|TNFSF14 protein, human|Drug|false|false||lightnull|Light - subjective measurement|Finding|false|false||light
null|TNFSF14 wt Allele|Finding|false|false||light
null|TNFSF14 gene|Finding|false|false||light
null|Light color|Finding|false|false||lightnull|Phototherapy|Procedure|false|false||lightnull|Light|Phenomenon|false|false||lightnull|Light (qualifier)|Modifier|false|false||lightnull|Touch Perception|Finding|false|false||touch
null|Touch sensation|Finding|false|false||touchnull|Therapeutic Touch|Procedure|false|false||touchnull|Tactile|Modifier|false|false||touchnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Rh Negative Blood Group|Finding|false|false||Negative
null|Negative|Finding|false|false||Negative
null|Negative Finding|Finding|false|false||Negativenull|Expression Negative|Lab|false|false||Negativenull|Negative - qualifier|Modifier|false|false||Negative
null|Negative Charge|Modifier|false|false||Negativenull|Negative Number|LabModifier|false|false||Negativenull|Hallway|Device|false|false||hallwaynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Bone structure of tibia|Anatomy|false|false||tibialnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|IL5 protein, human|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|thyrotropin-releasing hormone|Drug|false|false||TRF
null|Tocotrienol-rich Fraction|Drug|false|false||TRF
null|Thyrotropin-Releasing Hormone, human|Drug|false|false||TRFnull|TERF1 wt Allele|Finding|false|false||TRF
null|TERF1 gene|Finding|false|false||TRF
null|IL5 gene|Finding|false|false||TRFnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Mandibular right central incisor mesial prosthesis|Device|false|false||25PMnull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Leukocytes|Anatomy|false|false||WBCnull|Erythrocytes|Drug|false|false||RBCnull|Erythrocytes|Anatomy|false|false||RBCnull|null|Attribute|false|false||RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Structure of vein of lower extremity|Anatomy|false|false||lower extremity vein
null|Lower extremity>Lower extremity veins|Anatomy|false|false||lower extremity veinnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Venous structure of limb|Anatomy|false|false||extremity veinnull|Limb structure|Anatomy|false|false||extremitynull|Veins|Anatomy|false|false||veinnull|Posterior part of right leg|Anatomy|true|false||Right calfnull|Table Cell Horizontal Align - right|Finding|true|false||Rightnull|Right sided|Modifier|true|false||Right
null|Right|Modifier|true|false||Rightnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Deep Resection Margin|Attribute|true|false||deepnull|Deep (qualifier value)|Modifier|true|false||deepnull|Venous thrombosis after immobility|Finding|true|false||venous thrombosis
null|Venous Thrombosis|Finding|true|false||venous thrombosisnull|Veins|Anatomy|true|false||venousnull|Venous|Modifier|true|false||venousnull|Thrombosis|Finding|true|false||thrombosisnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower extremity>Lower extremity veins|Anatomy|false|false||lower extremity veins
null|Structure of vein of lower extremity|Anatomy|false|false||lower extremity veinsnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Venous structure of limb|Anatomy|false|false||extremity veinsnull|Limb structure|Anatomy|false|false||extremitynull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|null|Modifier|false|false||Unremarkablenull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Posterior part of right leg|Anatomy|false|false||right calfnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Vessel Positions|Anatomy|false|false||vessel
null|Blood Vessel|Anatomy|false|false||vesselnull|Vessel (unit of presentation)|LabModifier|false|false||vesselnull|Runoff|Modifier|false|false||runoffnull|Foot problem|Finding|false|false||footnull|Lower extremity>Foot|Anatomy|false|false||foot
null|Foot|Anatomy|false|false||footnull|Foot Unit of Length|LabModifier|false|false||footnull|Procedure on vein|Procedure|true|false||veinsnull|Veins|Anatomy|true|false||veinsnull|Lower Extremity|Anatomy|true|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|true|false||lowernull|Lower (action)|Event|true|false||lowernull|Lower - spatial qualifier|Modifier|true|false||lowernull|Limb structure|Anatomy|true|false||extremitynull|Views for patency|Modifier|true|false||patency
null|Open|Modifier|true|false||patencynull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|More|LabModifier|false|false||morenull|Focal|Modifier|true|false||focalnull|Collection Object - UML Entity|Finding|true|false||collection
null|Item Collection|Finding|true|false||collection
null|Collections (publication)|Finding|true|false||collection
null|Collection (action)|Finding|true|false||collectionnull|Obvious|Modifier|true|false||obviousnull|Abnormality of the musculature|Disorder|true|false||muscular abnormalitynull|Muscle (organ)|Anatomy|true|false||muscularnull|Muscular|Modifier|true|false||muscularnull|Congenital Abnormality|Disorder|true|false||abnormalitynull|Abnormality|Finding|true|false||abnormalitynull|Uneventful|Finding|false|false||Uneventfulnull|Ultrasonic|Finding|false|false||ultrasoundnull|Urological ultrasound|Procedure|false|false||ultrasound
null|Ultrasonography|Procedure|false|false||ultrasoundnull|ultrasound device|Device|false|false||ultrasoundnull|Ultrasonic Shockwave|Phenomenon|false|false||ultrasound
null|Ultrasonics (sound)|Phenomenon|false|false||ultrasoundnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Long Variable|Modifier|false|false||long
null|Long|Modifier|false|false||longnull|Anesthetic [APC]|Drug|false|false||anesthetic
null|Anesthetics|Drug|false|false||anestheticnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Greater|LabModifier|false|false||greaternull|Structure of trochanteric bursa|Anatomy|false|false||trochanteric bursanull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|null|Time|false|false||Priornull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Small amount|LabModifier|false|false||small amountnull|Small|LabModifier|false|false||smallnull|Amount class - Amount|Finding|false|false||amountnull|Quantity|LabModifier|false|false||amountnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Greater|LabModifier|false|false||greaternull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|Dystrophic calcification|Finding|false|false||dystrophic calcificationnull|dystrophic|Finding|false|false||dystrophicnull|Physiologic calcification|Finding|false|false||calcification
null|Calcification|Finding|false|false||calcification
null|Calcinosis|Finding|false|false||calcificationnull|Calcified (qualifier value)|Modifier|false|false||calcificationnull|bursal|Modifier|false|false||bursalnull|Space (Astronomy)|Phenomenon|false|false||spacenull|Space - property|Modifier|false|false||spacenull|Suspicion|Finding|false|false||suspicionnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|PMH - past medical history|Finding|false|false||PMH
null|Medical History|Finding|false|false||PMHnull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid syndromenull|Syndrome|Disorder|false|false||syndromenull|Deep thrombophlebitis|Disorder|false|false||DVTsnull|Personal Experience Scales|Finding|false|false||PEs
null|PES1 gene|Finding|false|false||PEsnull|Structure of ankle and/or foot (body structure)|Anatomy|false|false||PEs
null|Hindfoot of quadruped|Anatomy|false|false||PEs
null|Paw|Anatomy|false|false||PEs
null|Foot|Anatomy|false|false||PEsnull|Iranian Persian language|Entity|false|false||PEsnull|Coumadin|Drug|false|false||Coumadin
null|Coumadin|Drug|false|false||Coumadinnull|Recent|Time|false|false||recentnull|Malignant neoplasm of breast|Disorder|false|false||breast cancer
null|Breast Carcinoma|Disorder|false|false||breast cancernull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Malignant Neoplasms|Disorder|false|false||cancernull|Specialty Type - cancer|Title|false|false||cancernull|Cancer <Cancridae>|Entity|false|false||cancernull|Lumpectomy of breast|Procedure|false|false||lumpectomy
null|Excision of mass (procedure)|Procedure|false|false||lumpectomynull|Acute-on-chronic|Time|false|false||acute on chronicnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Right lower extremity|Anatomy|false|false||right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Pain of right hip joint|Finding|false|false||right hip painnull|Right hip region structure|Anatomy|false|false||right hipnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Hip joint pain|Finding|false|false||hip pain
null|Hip pain|Finding|false|false||hip painnull|null|Attribute|false|false||hip painnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Right lower extremity|Anatomy|false|false||Right lower extremitynull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Lower Extremity|Anatomy|false|false||lower extremitynull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Limb structure|Anatomy|false|false||extremitynull|Deep thrombophlebitis|Disorder|true|false||DVT
null|Deep Vein Thrombosis|Disorder|true|false||DVTnull|area DVT|Anatomy|true|false||DVTnull|null|Attribute|true|false||DVTnull|Structure of calf of leg|Anatomy|true|false||calf
null|null|Anatomy|true|false||calfnull|Cattle calf (organism)|Entity|true|false||calfnull|Procedure on vein|Procedure|true|false||veinsnull|Veins|Anatomy|true|false||veinsnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|true|false||well
null|Good|Modifier|true|false||well
null|Healthy|Modifier|true|false||wellnull|right trochanteric bursitis|Disorder|false|false||Right trochanteric bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Right anterior|Modifier|false|false||Right anteriornull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Lower anterior|Modifier|false|false||anterior lowernull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Pain in limb, lower leg|Finding|false|false||lower leg pain
null|Pain in lower limb|Finding|false|false||lower leg painnull|Lower extremity>Lower leg|Anatomy|false|false||lower leg
null|Leg|Anatomy|false|false||lower legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Pain in lower limb|Finding|false|false||leg painnull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Right sided|Modifier|false|false||Right sided
null|Right|Modifier|false|false||Right sidednull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Observation Interpretation - worse|Finding|false|false||worse
null|Worse|Finding|false|false||worsenull|Worsening (qualifier value)|Modifier|false|false||worsenull|Last|Modifier|false|false||lastnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Focal|Modifier|false|false||focalnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Right tibia|Anatomy|false|false||right tibianull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Bone structure of tibia|Anatomy|false|false||tibianull|Tibia <Rostellariidae>|Entity|false|false||tibianull|Consistent with|Finding|false|false||consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false||consistentnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|X-RAY SENSITIVITY|Finding|false|false||XRsnull|Bone structure of tibia|Anatomy|true|false||tibianull|Tibia <Rostellariidae>|Entity|true|false||tibianull|Fibula|Anatomy|true|false||fibulanull|Right hip region structure|Anatomy|true|false||right hipnull|Table Cell Horizontal Align - right|Finding|true|false||rightnull|Right sided|Modifier|true|false||right
null|Right|Modifier|true|false||rightnull|heme iron polypeptide|Drug|true|false||hip
null|ST13 protein, human|Drug|true|false||hip
null|ST13 protein, human|Drug|true|false||hip
null|RPL29 protein, human|Drug|true|false||hip
null|RPL29 protein, human|Drug|true|false||hip
null|HHIP protein, human|Drug|true|false||hip
null|HHIP protein, human|Drug|true|false||hip
null|heme iron polypeptide|Drug|true|false||hipnull|RPL29 wt Allele|Finding|true|false||hip
null|REG3A gene|Finding|true|false||hip
null|RPL29 gene|Finding|true|false||hip
null|ST13 wt Allele|Finding|true|false||hip
null|ST13 gene|Finding|true|false||hip
null|HHIP gene|Finding|true|false||hip
null|HHIP wt Allele|Finding|true|false||hip
null|REG3A wt Allele|Finding|true|false||hipnull|Procedure on hip|Procedure|true|false||hipnull|Lower extremity>Hip|Anatomy|true|false||hip
null|Hip structure|Anatomy|true|false||hip
null|Structure of habenulopeduncular tract|Anatomy|true|false||hip
null|Bone structure of ischium|Anatomy|true|false||hipnull|Obvious|Modifier|true|false||obviousnull|Pathology processes|Finding|true|false||pathology
null|Pathological aspects|Finding|true|false||pathologynull|Pathology procedure|Procedure|true|false||pathologynull|Pathology|Title|true|false||pathologynull|Neurologic Symptoms|Finding|true|false||neurologic symptomsnull|Neurologic (qualifier value)|Modifier|true|false||neurologicnull|Symptoms aspect|Finding|true|false||symptoms
null|Symptoms|Finding|true|false||symptomsnull|Radiculopathy|Disorder|true|false||radiculopathynull|Weakness|Finding|true|false||weakness
null|Asthenia|Finding|true|false||weaknessnull|Numbness|Finding|true|false||numbness
null|Hypesthesia|Finding|true|false||numbnessnull|Academic degree|Finding|false|false||degreenull|Levels (qualifier value)|Modifier|false|false||degreenull|Degree Unit of Plane Angle|LabModifier|false|false||degree
null|Degree or extent|LabModifier|false|false||degreenull|Chronic sciatica|Disorder|false|false||chronic sciaticanull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Sciatica|Finding|false|false||sciaticanull|Mildly decreased|Finding|false|false||Mildly decreasednull|MILDLY|Modifier|false|false||Mildly
null|Mild (qualifier value)|Modifier|false|false||Mildlynull|Decreased patellar reflex|Finding|false|false||decreased patellar reflexnull|Knee reflex|Finding|false|false||patellar reflexnull|Patella|Anatomy|false|false||patellarnull|Reflex motion descriptor|Finding|false|false||reflex
null|Reflex action|Finding|false|false||reflex
null|Observation of reflex|Finding|false|false||reflexnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Protective muscle spasm|Finding|false|false||guardingnull|Strength (attribute)|Finding|false|false||strengthnull|Pharmaceutical Strength|LabModifier|false|false||strength
null|Physical Strength|LabModifier|false|false||strengthnull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Injection of steroid|Procedure|false|false||steroid injectionnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|Improvement|Finding|false|false||improvementnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|fluid - substance|Drug|false|false||fluid
null|Liquid substance|Drug|false|false||fluidnull|Fluid Specimen Code|Finding|false|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Synovial bursa|Anatomy|false|false||bursanull|Bursa <Bursidae>|Entity|false|false||bursanull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|shin pain|Finding|false|false||shin painnull|Shin|Anatomy|false|false||shinnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Transcription Initiation|Finding|false|false||initiation
null|Initiation|Finding|false|false||initiation
null|null|Finding|false|false||initiationnull|AOD use initiation|Time|false|false||initiationnull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|Lidocaine Patch|Drug|false|false||lidocaine patchnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Patch - Extended Release Film|Drug|false|false||patch
null|Human patch material|Drug|false|false||patch
null|Body tissue patch material|Drug|false|false||patchnull|Plaque (lesion)|Finding|false|false||patchnull|Patch Dosage Form|Device|false|false||patch
null|Surgical patch|Device|false|false||patchnull|Patch (unit of presentation)|LabModifier|false|false||patch
null|Patch Dosing Unit|LabModifier|false|false||patchnull|In addition to|Finding|false|false||in addition tonull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Tylenol|Drug|false|false||tylenol
null|Tylenol|Drug|false|false||tylenolnull|Increase|Finding|false|false||increasenull|Frequency|Finding|false|false||frequency
null|How Often|Finding|false|false||frequencynull|With frequency|Time|false|false||frequency
null|Frequencies (time pattern)|Time|false|false||frequencynull|Kind of quantity - Frequency|LabModifier|false|false||frequency
null|Statistical Frequency|LabModifier|false|false||frequency
null|Spatial Frequency|LabModifier|false|false||frequencynull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Every eight hours|Time|false|false||q8hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Every four hours|Time|false|false||q4hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Visit User Code - Home|Finding|true|false||home
null|Address type - Home|Finding|true|false||homenull|home health encounter|Procedure|true|false||homenull|Organization unit type - Home|Entity|true|false||homenull|Person location type - Home|Modifier|true|false||home
null|Home environment|Modifier|true|false||homenull|hydromorphone|Drug|true|false||hydromorphone
null|hydromorphone|Drug|true|false||hydromorphonenull|CIAO3 gene|Finding|true|false||PRNnull|As required|Time|true|false||PRN
null|Pro Re Nata|Time|true|false||PRNnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|hydromorphone|Drug|false|false||hydromorphone
null|hydromorphone|Drug|false|false||hydromorphonenull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Episode of|Time|false|false||episodenull|tramadol|Drug|false|false||Tramadol
null|tramadol|Drug|false|false||Tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||Tramadolnull|Tablet Dosage Form|Drug|false|false||tabletsnull|Increased metabolic requirement|Finding|false|false||increased requirementnull|Requirement|Finding|false|false||requirementnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|Ambulate|Finding|false|false||ambulatenull|SAFE-Biopharma Standard|Finding|false|false||safenull|Discharge to home|Procedure|false|false||discharge homenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|Processing type - Evaluation|Finding|false|false||evaluationnull|Evaluation procedure|Procedure|false|false||evaluation
null|Evaluation|Procedure|false|false||evaluationnull|Enthusiastic|Finding|false|false||eagernull|Vascular surgeon|Subject|false|false||vascular surgeonnull|Blood Vessel|Anatomy|false|false||vascularnull|Vascular|Modifier|false|false||vascularnull|null|Attribute|false|false||surgeonnull|Surgeon|Subject|false|false||surgeonnull|Appointments|Event|false|false||appointmentnull|Early|Time|false|false||earlynull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Transaction counts and value totals - year|Finding|false|false||year
null|Precision - year|Finding|false|false||yearnull|year|Time|false|false||yearnull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Pain|Finding|false|false||painfulnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Iron deficiency anemia|Disorder|false|false||Iron deficiency anemianull|Iron deficiency anemia|Disorder|false|false||Iron deficiency
null|Iron deficiency|Disorder|false|false||Iron deficiencynull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Deficiency anemias|Disorder|false|false||deficiency anemianull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Anemia|Disorder|false|false||Anemianull|Anemia <Anemiaceae>|Entity|false|false||Anemianull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Overnight|Time|false|false||overnightnull|Concern|Finding|true|false||concernnull|Hemorrhage|Finding|true|false||bleedingnull|iron studies|Procedure|false|false||iron studiesnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Scientific Study|Procedure|false|false||studiesnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Deficiency|Finding|false|false||deficientnull|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritin
null|Ferritin|Drug|false|false||ferritinnull|Ferritin measurement|Procedure|false|false||ferritinnull|Fatigue|Finding|false|false||fatiguenull|Restless Legs Syndrome|Disorder|false|false||restless leg syndromenull|Restless Legs Syndrome|Disorder|false|false||restless legnull|Restlessness|Finding|false|false||restless
null|Agitation|Finding|false|false||restlessnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Syndrome|Disorder|false|false||syndromenull|Science of Etiology|Finding|false|false||Etiology
null|Etiology aspects|Finding|false|false||Etiology
null|Etiology|Finding|false|false||Etiologynull|Recent|Time|false|false||recentnull|Left breast|Anatomy|false|false||left breastnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Breast hematoma|Finding|false|false||breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Hematoma|Finding|false|false||hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Unlikely|Finding|false|false||unlikelynull|Unlikely Related to Intervention|Modifier|false|false||unlikelynull|Timing, LOINC Axis 3|Finding|false|false||timingnull|Timing|Time|false|false||timingnull|Seizures|Finding|false|false||fitsnull|null|Time|false|false||Priornull|Esophagogastroduodenoscopy|Procedure|false|false||EGDnull|Gastritis|Disorder|false|false||gastritisnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Proton Pump Inhibitors|Drug|false|false||PPInull|Prepulse Inhibition|Finding|false|false||PPInull|null|Time|false|false||priornull|Consent Type - Colonoscopy|Procedure|false|false||colonoscopy
null|colonoscopy|Procedure|false|false||colonoscopynull|findings aspects|Finding|false|false||findingsnull|null|Attribute|false|false||findingsnull|Suggestive of|Finding|false|false||suggestive ofnull|Suggestive of|Finding|false|false||suggestivenull|Celiac Disease|Disorder|false|false||celiac diseasenull|CTLA4 gene|Finding|false|false||celiac diseasenull|Celiac Disease|Disorder|false|false||celiacnull|Disease|Disorder|false|false||diseasenull|TGM2 protein, human|Drug|false|false||ttg
null|TGM2 protein, human|Drug|false|false||ttg
null|TGM2 protein, human|Drug|false|false||ttgnull|TGM2 wt Allele|Finding|false|false||ttgnull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|immunoglobulin A, human|Drug|false|false||IgA
null|immunoglobulin A|Drug|false|false||IgA
null|immunoglobulin A|Drug|false|false||IgA
null|immunoglobulin A, human|Drug|false|false||IgAnull|CD79A wt Allele|Finding|false|false||IgA
null|CD79A gene|Finding|false|false||IgAnull|Immunoglobulin A measurement|Procedure|false|false||IgAnull|polyps|Disorder|false|false||polypsnull|null|Finding|false|false||polypsnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Vitamins A and D preparation|Drug|false|false||a vitamin Dnull|vitamin A|Drug|false|false||a vitamin
null|vitamin A|Drug|false|false||a vitamin
null|vitamin A|Drug|false|false||a vitaminnull|Vitamin D Drug Class|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|D Vitamin|Drug|false|false||vitamin D
null|Vitamin D [EPC]|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|Vitamin D Drug Class|Drug|false|false||vitamin Dnull|Vitamin D measurement|Procedure|false|false||vitamin Dnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Evidence|Finding|false|false||evidencenull|Malabsorption Syndrome|Disorder|false|false||malabsorptionnull|Malabsorption|Finding|false|false||malabsorptionnull|Iso|Entity|false|false||isonull|Daily|Time|false|false||dailynull|Dietary Supplementation|Procedure|false|false||supplementationnull|ferric gluconate|Drug|false|false||ferric gluconate
null|ferric gluconate|Drug|false|false||ferric gluconatenull|ferric cation|Drug|false|false||ferric
null|ferric cation|Drug|false|false||ferricnull|gluconate|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|Gluconates|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconate
null|gluconate|Drug|false|false||gluconatenull|TGM2 protein, human|Drug|false|false||TTG
null|TGM2 protein, human|Drug|false|false||TTG
null|TGM2 protein, human|Drug|false|false||TTGnull|TGM2 wt Allele|Finding|false|false||TTGnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|Anticoagulation drug level below therapeutic|Finding|false|false||Subtherapeutic INRnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Lupus anticoagulant positive|Lab|false|false||Lupus anticoagulant positivenull|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulant
null|Lupus Coagulation Inhibitor|Drug|false|false||Lupus anticoagulantnull|Lupus anticoagulant disorder|Disorder|false|false||Lupus anticoagulantnull|null|Finding|false|false||Lupus anticoagulantnull|Lupus anticoagulant assay|Procedure|false|false||Lupus anticoagulantnull|Chronic discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus|Disorder|false|false||Lupus
null|Lupus Vulgaris|Disorder|false|false||Lupus
null|Discoid lupus erythematosus|Disorder|false|false||Lupus
null|Lupus Erythematosus, Systemic|Disorder|false|false||Lupusnull|Anti-coagulant [EPC]|Drug|false|false||anticoagulant
null|Anticoagulants|Drug|false|false||anticoagulantnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|day|Time|false|false||daysnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Last|Modifier|false|false||lastnull|Hematoma|Finding|false|false||hematomanull|Lovenox|Drug|true|false||Lovenox
null|Lovenox|Drug|true|false||Lovenoxnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Hospitalization|Procedure|false|false||hospitalizationnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Daily|Time|false|false||dailynull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Continuous|Finding|false|false||continuenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Vitamin D Deficiency|Disorder|false|false||Vitamin D deficiencynull|Decreased circulating vitamin D concentration|Finding|false|false||Vitamin D deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Vitamin D Drug Class|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|vitamin D|Drug|false|false||vitamin D
null|D Vitamin|Drug|false|false||vitamin D
null|Vitamin D [EPC]|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|ergocalciferol|Drug|false|false||vitamin D
null|Vitamin D Drug Class|Drug|false|false||vitamin Dnull|Vitamin D measurement|Procedure|false|false||vitamin Dnull|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Daily|Time|false|false||dailynull|Repeat Object|Finding|false|false||Repeat
null|Repeat|Finding|false|false||Repeatnull|Repeat Pattern|Time|false|false||Repeatnull|Malabsorption Syndrome|Disorder|false|false||malabsorptionnull|Malabsorption|Finding|false|false||malabsorptionnull|Iron deficiency anemia|Disorder|false|false||iron deficiency
null|Iron deficiency|Disorder|false|false||iron deficiencynull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|CODE STATUS|Procedure|false|false||Code statusnull|MDF Attribute Type - Code|Finding|false|false||Code
null|A Codes|Finding|false|false||Code
null|Code|Finding|false|false||Codenull|Coding|Event|false|false||Codenull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|Full|Modifier|false|false||Fullnull|Hereditary Coproporphyria|Disorder|false|false||HCPnull|PTPN6 wt Allele|Finding|false|false||HCP
null|CPOX gene|Finding|false|false||HCP
null|AMBP wt Allele|Finding|false|false||HCP
null|PTPN6 gene|Finding|false|false||HCP
null|AMBP gene|Finding|false|false||HCPnull|Granddaughter|Subject|false|false||granddaughternull|right trochanteric bursitis|Disorder|false|false||Right trochanteric bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Diagnostic Service Section ID - Physical Therapy|Finding|false|false||physical therapynull|Physical therapy|Procedure|false|false||physical therapynull|Physical therapy (field)|Title|false|false||physical therapynull|physical examination (physical finding)|Finding|false|false||physical
null|Physical|Finding|false|false||physicalnull|Physical Examination|Procedure|false|false||physicalnull|Therapy Object (animal model)|Finding|false|false||therapy
null|therapeutic aspects|Finding|false|false||therapynull|Therapeutic procedure|Procedure|false|false||therapynull|Right anterior|Modifier|false|false||Right anteriornull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|Three times daily|Time|false|false||three times dailynull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|during hospitalization|Time|false|false||during hospitalizationnull|Hospitalization|Procedure|false|false||hospitalizationnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Supply (process)|Finding|false|false||supply
null|Supply (system)|Finding|false|false||supply
null|supply aspects|Finding|false|false||supplynull|Healthcare supplies|Device|false|false||supplynull|Providing (action)|Event|false|false||supplynull|supply & distribution|LabModifier|false|false||supply
null|Economic supply|LabModifier|false|false||supplynull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||Plannull|Treatment Plan|Finding|false|false||Plan
null|Planned|Finding|false|false||Plan
null|null|Finding|false|false||Plannull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|next - HtmlLinkType|Finding|false|false||nextnull|Following|Time|false|false||next
null|Then|Time|false|false||nextnull|Adjacent|Modifier|false|false||nextnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Bone structure of lumbar vertebra|Anatomy|false|false||lumbar spine
null|Lumbar spine structure|Anatomy|false|false||lumbar spinenull|Lumbar Region|Anatomy|false|false||lumbarnull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|chronic pain (diagnosis)|Disorder|false|false||chronic painnull|Chronic pain|Finding|false|false||chronic painnull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Electromyogram of eye|Procedure|false|false||EMG
null|Electromyography|Procedure|false|false||EMGnull|Electromyographs|Device|false|false||EMGnull|Vascular Surgical Procedures|Procedure|false|false||Vascular surgerynull|Vascular surgery specialty|Title|false|false||Vascular surgerynull|Blood Vessel|Anatomy|false|false||Vascularnull|Vascular|Modifier|false|false||Vascularnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Biomaterial Treatment|Finding|false|false||treatment
null|Treating|Finding|false|false||treatment
null|therapeutic aspects|Finding|false|false||treatmentnull|treatment - ActInformationManagementReason|Procedure|false|false||treatment
null|Administration (procedure)|Procedure|false|false||treatment
null|Therapeutic procedure|Procedure|false|false||treatmentnull|Pain|Finding|false|false||painfulnull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Iron deficiency anemia|Disorder|false|false||Iron deficiency anemianull|Iron deficiency anemia|Disorder|false|false||Iron deficiency
null|Iron deficiency|Disorder|false|false||Iron deficiencynull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Deficiency anemias|Disorder|false|false||deficiency anemianull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|ferryl iron|Drug|false|false||IV ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|Pending - Allergy Clinical Status|Finding|false|false||pending
null|Pending - referral status|Finding|false|false||pendingnull|Pending - status|Time|false|false||pendingnull|pending - ManagedParticipationStatus|Modifier|false|false||pending
null|pending - RoleStatus|Modifier|false|false||pending
null|Pending - Day type|Modifier|false|false||pendingnull|TGM2 protein, human|Drug|false|false||TTG
null|TGM2 protein, human|Drug|false|false||TTG
null|TGM2 protein, human|Drug|false|false||TTGnull|TGM2 wt Allele|Finding|false|false||TTGnull|Further|Modifier|false|false||furthernull|Relate - vinyl resin|Drug|false|false||relatednull|Role Link Type - related|Finding|false|false||related
null|Related (finding)|Finding|false|false||relatednull|Definitely Related to Intervention|Modifier|false|false||related
null|Relationships|Modifier|false|false||relatednull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Breast hematoma|Finding|false|false||breast hematomanull|Neoplasm of uncertain or unknown behavior of breast|Disorder|false|false||breastnull|Breast problem|Finding|false|false||breastnull|Procedures on breast|Procedure|false|false||breastnull|Breast|Anatomy|false|false||breastnull|Hematoma|Finding|false|false||hematomanull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|Antiphospholipid Syndrome|Disorder|false|false||antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|Anticoagulation drug level below therapeutic|Finding|false|false||subtherapeutic INRnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Clinic|Device|false|false||clinic
null|Ambulatory Care Facilities|Device|false|false||clinicnull|Clinic|Entity|false|false||clinic
null|Ambulatory Care Facilities|Entity|false|false||clinicnull|Patient location type - Clinic|Modifier|false|false||clinic
null|Person location type - Clinic|Modifier|false|false||clinicnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|Indication of (contextual qualifier)|Finding|false|false||Reason fornull|Indication of (contextual qualifier)|Finding|false|false||Reasonnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Duplicate component (foundation metadata concept)|Finding|false|false||duplicate
null|Double (qualifier value)|Finding|false|false||duplicatenull|Replicate|Event|false|false||duplicatenull|Duplicate|Modifier|false|false||duplicatenull|Override|Finding|false|false||overridenull|Similarity|Modifier|false|false||similarnull|With intensity|Modifier|false|false||severity
null|Severities|Modifier|false|false||severitynull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|erythromycin|Drug|false|false||Erythromycin
null|erythromycin|Drug|false|false||Erythromycinnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Ointments|Drug|false|false||Ointnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|Four times daily|Time|false|false||QIDnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false||Leg swellingnull|Leg|Anatomy|false|false||Leg
null|Lower Extremity|Anatomy|false|false||Legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|hydromorphone|Drug|false|false||HYDROmorphone
null|hydromorphone|Drug|false|false||HYDROmorphonenull|Dilaudid|Drug|false|false||Dilaudid
null|Dilaudid|Drug|false|false||Dilaudidnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Three times daily|Time|false|false||three times dailynull|Thrice|LabModifier|false|false||three timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false||PTCH
null|PTCH1 wt Allele|Finding|false|false||PTCH
null|PTCH1 gene|Finding|false|false||PTCH
null|PTCH1 protein, human|Finding|false|false||PTCHnull|Every morning|Time|false|false||QAMnull|Right hip region structure|Anatomy|false|false||right hipnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|heme iron polypeptide|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|ST13 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|RPL29 protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|HHIP protein, human|Drug|false|false||hip
null|heme iron polypeptide|Drug|false|false||hipnull|RPL29 wt Allele|Finding|false|false||hip
null|REG3A gene|Finding|false|false||hip
null|RPL29 gene|Finding|false|false||hip
null|ST13 wt Allele|Finding|false|false||hip
null|ST13 gene|Finding|false|false||hip
null|HHIP gene|Finding|false|false||hip
null|HHIP wt Allele|Finding|false|false||hip
null|REG3A wt Allele|Finding|false|false||hipnull|Procedure on hip|Procedure|false|false||hipnull|Lower extremity>Hip|Anatomy|false|false||hip
null|Hip structure|Anatomy|false|false||hip
null|Structure of habenulopeduncular tract|Anatomy|false|false||hip
null|Bone structure of ischium|Anatomy|false|false||hipnull|lidocaine|Drug|false|false||lidocaine
null|lidocaine|Drug|false|false||lidocainenull|Lidocaine measurement|Procedure|false|false||lidocainenull|Apply (administration method)|Finding|false|false||Apply
null|Apply (instruction)|Finding|false|false||Apply
null|null|Finding|false|false||Apply
null|Apply|Finding|false|false||Applynull|Patch Dosage Form|Device|false|false||patchesnull|Daily|Time|false|false||dailynull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|refill|Finding|false|false||Refillsnull|tramadol|Drug|false|false||TraMADol
null|tramadol|Drug|false|false||TraMADolnull|Tramadol measurement (procedure)|Procedure|false|false||TraMADolnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|tramadol|Drug|false|false||tramadol
null|tramadol|Drug|false|false||tramadolnull|Tramadol measurement (procedure)|Procedure|false|false||tramadolnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false||by mouthnull|Oral cavity|Anatomy|false|false||mouth
null|Oral region|Anatomy|false|false||mouthnull|Every six hours|Time|false|false||Every six hoursnull|Every - dosing instruction fragment|Finding|false|false||Everynull|Every (qualifier)|Modifier|false|false||Everynull|Hour|Time|false|false||hoursnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Fever symptoms (finding)|Finding|false|false||Fever
null|Fever|Finding|false|false||Fevernull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|NEB protein, human|Drug|false|false||NEB
null|NEB protein, human|Drug|false|false||NEB
null|Nebulizer solution|Drug|false|false||NEBnull|NEB gene|Finding|false|false||NEB
null|mitotic nuclear membrane disassembly|Finding|false|false||NEBnull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Wheezing|Finding|false|false||wheezenull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|erythromycin|Drug|false|false||Erythromycin
null|erythromycin|Drug|false|false||Erythromycinnull|Ophthalmic Route of Administration|Finding|false|false||Ophthnull|Ointments|Drug|false|false||Ointnull|Structure of both eyes|Anatomy|false|false||BOTH EYESnull|Eye|Anatomy|false|false||EYESnull|null|Attribute|false|false||EYESnull|Four times daily|Time|false|false||QIDnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Swelling of lower limb|Finding|false|false||Leg swellingnull|Leg|Anatomy|false|false||Leg
null|Lower Extremity|Anatomy|false|false||Legnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|omeprazole|Drug|false|false||Omeprazole
null|omeprazole|Drug|false|false||Omeprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|polyethylene glycols|Drug|false|false||Polyethylene Glycol
null|polyethylene glycols|Drug|false|false||Polyethylene Glycolnull|high-density polyethylene|Drug|false|false||Polyethylene
null|high-density polyethylene|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|polyethylenes|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylene
null|Polyethylene|Drug|false|false||Polyethylenenull|ethylene glycol|Drug|false|false||Glycol
null|Glycol|Drug|false|false||Glycol
null|ethylene glycol|Drug|false|false||Glycol
null|Glycols|Drug|false|false||Glycolnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|sertraline|Drug|false|false||Sertraline
null|sertraline|Drug|false|false||Sertralinenull|Daily|Time|false|false||DAILYnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleep
null|Sleep brand of diphenhydramine hydrochloride|Drug|false|false||sleepnull|Sleep|Finding|false|false||sleepnull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Storage Unit|Device|false|false||UNIT
null|Unit device|Device|false|false||UNITnull|Unit - NCI Thesaurus Property|LabModifier|false|false||UNIT
null|Unit of Measure|LabModifier|false|false||UNIT
null|Unit|LabModifier|false|false||UNIT
null|Enzyme Unit|LabModifier|false|false||UNITnull|Daily|Time|false|false||DAILYnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarin
null|warfarin|Drug|false|false||Warfarinnull|Weekly|Time|false|false||/WEEKnull|Transaction counts and value totals - week|Finding|false|false||WEEKnull|week|Time|false|false||WEEKnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|True primary (qualifier value)|Time|false|false||PRIMARYnull|Primary|Modifier|false|false||PRIMARYnull|right trochanteric bursitis|Disorder|false|false||Right trochanteric bursitisnull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Greater trochanteric pain syndrome|Disorder|false|false||trochanteric bursitisnull|Bursitis|Disorder|false|false||bursitisnull|Right anterior|Modifier|false|false||Right anteriornull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Adenohypophyseal Diseases|Disorder|false|false||anteriornull|Anterior|Modifier|false|false||anteriornull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Right sided|Modifier|false|false||Right sided
null|Right|Modifier|false|false||Right sidednull|Table Cell Horizontal Align - right|Finding|false|false||Rightnull|Right sided|Modifier|false|false||Right
null|Right|Modifier|false|false||Rightnull|Varicosity|Disorder|false|false||varicose veinsnull|Varicose|Modifier|false|false||varicosenull|Procedure on vein|Procedure|false|false||veinsnull|Veins|Anatomy|false|false||veinsnull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Iron deficiency anemia|Disorder|false|false||Iron deficiency anemianull|Iron deficiency anemia|Disorder|false|false||Iron deficiency
null|Iron deficiency|Disorder|false|false||Iron deficiencynull|Iron Drug Class|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|iron|Drug|false|false||Iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||Ironnull|Iron measurement|Procedure|false|false||Ironnull|Deficiency anemias|Disorder|false|false||deficiency anemianull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Anemia|Disorder|false|false||anemianull|Anemia <Anemiaceae>|Entity|false|false||anemianull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Deep thrombophlebitis|Disorder|false|false||DVT
null|Deep Vein Thrombosis|Disorder|false|false||DVTnull|area DVT|Anatomy|false|false||DVTnull|null|Attribute|false|false||DVTnull|on warfarin|Procedure|false|false||on warfarinnull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Antiphospholipid Syndrome|Disorder|false|false||Antiphospholipid antibody syndromenull|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibody
null|Antiphospholipid Antibodies|Drug|false|false||Antiphospholipid antibodynull|Antiphospholipid antibody positivity|Finding|false|false||Antiphospholipid antibodynull|Immunoglobulins|Drug|false|false||antibody
null|Immunoglobulins|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibody
null|Antibodies|Drug|false|false||antibodynull|Antibody (immunoassay)|Procedure|false|false||antibodynull|Immunoglobulin complex location, circulating|Anatomy|false|false||antibody
null|immunoglobulin complex location|Anatomy|false|false||antibodynull|Syndrome|Disorder|false|false||syndromenull|Anticoagulation drug level below therapeutic|Finding|false|false||Subtherapeutic INRnull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|Vitamin D Deficiency|Disorder|false|false||Vitamin D deficiencynull|Decreased circulating vitamin D concentration|Finding|false|false||Vitamin D deficiencynull|Vitamin D Drug Class|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|vitamin D|Drug|false|false||Vitamin D
null|D Vitamin|Drug|false|false||Vitamin D
null|Vitamin D [EPC]|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|ergocalciferol|Drug|false|false||Vitamin D
null|Vitamin D Drug Class|Drug|false|false||Vitamin Dnull|Vitamin D measurement|Procedure|false|false||Vitamin Dnull|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitamin
null|Vitamins|Drug|false|false||Vitaminnull|Malnutrition|Disorder|false|false||deficiencynull|Deficiency|Finding|false|false||deficiencynull|deficiency aspects|Modifier|false|false||deficiencynull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Helping Behavior|Finding|false|false||assistancenull|Assisted (qualifier value)|Modifier|false|false||assistancenull|AICDA protein, human|Drug|false|false||aid
null|AICDA protein, human|Drug|false|false||aidnull|AICDA wt Allele|Finding|false|false||aid
null|AICDA gene|Finding|false|false||aidnull|AID - Artificial insemination by donor|Procedure|false|false||aid
null|dacarbazine/doxorubicin/ifosfamide protocol|Procedure|false|false||aidnull|Aid (attribute)|Modifier|false|false||aid
null|Assisted (qualifier value)|Modifier|false|false||aidnull|Walkers|Device|false|false||walkernull|CANE, INCLUDES CANES OF ALL MATERIALS, ADJUSTABLE OR FIXED, WITH TIP|Device|false|false||canenull|Cane - plant part|Entity|false|false||canenull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Very Much|Finding|false|false||a lotnull|Stock (in-store merchandise)|Finding|false|false||lotnull|nucleus of the lateral olfactory tract|Anatomy|false|false||lot
null|Olfactory tract|Anatomy|false|false||lotnull|Lot (entire collection)|Modifier|false|false||lotnull|Pain in lower limb|Finding|false|false||leg painnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Difficult (qualifier value)|Finding|false|false||difficultnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Injection of steroid|Procedure|false|false||steroid injectionnull|Steroid [EPC]|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroid
null|Steroids|Drug|false|false||steroidnull|Injection|Drug|false|false||injectionnull|Injection Route of Administration|Finding|false|false||injectionnull|Injection of therapeutic agent|Procedure|false|false||injection
null|Injection procedure|Procedure|false|false||injectionnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Lower extremity>Thigh|Anatomy|false|false||thigh
null|Thigh structure|Anatomy|false|false||thighnull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Greater trochanteric pain syndrome|Disorder|false|false||Trochanteric Bursitisnull|Bursitis|Disorder|false|false||Bursitisnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Lovenox|Drug|false|false||Lovenox
null|Lovenox|Drug|false|false||Lovenoxnull|What subject filter - Order|Finding|false|false||order
null|Medical Order|Finding|false|false||order
null|Order (taxonomic)|Finding|false|false||order
null|Order (record artifact)|Finding|false|false||order
null|Order (document)|Finding|false|false||ordernull|Order [PK]|Phenomenon|false|false||ordernull|Order (action)|Event|false|false||ordernull|Order (arrangement)|Modifier|false|false||order
null|Permutation|Modifier|false|false||ordernull|Fixation of dental bridge|Procedure|false|false||bridgenull|Type of bridge device|Device|false|false||bridgenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Current (present time)|Time|false|false||currentlynull|warfarin dose|Procedure|false|false||warfarin dosenull|null|Attribute|false|false||warfarin dosenull|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarin
null|warfarin|Drug|false|false||warfarinnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Daily|Time|false|false||dailynull|Integrated Neuromusculoskeletal Release|Procedure|false|false||INR
null|International Normalized Ratio|Procedure|false|false||INRnull|Coagulation tissue factor induced.INR|Attribute|false|false||INRnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|objective (goal)|Finding|false|false||goal
null|Act Mood - Goal|Finding|false|false||goalnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Intravenous Route of Administration|Finding|false|false||intravenousnull|Intravenous|Modifier|false|false||intravenousnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Deficiency|Finding|false|false||deficientnull|More|LabModifier|false|false||morenull|Fatigue|Finding|false|false||fatiguednull|Usual|Modifier|false|false||usualnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Appointments|Event|false|false||appointmentnull|Primary care provider|Subject|false|false||primary care doctornull|Location Service Code - Primary Care|Finding|false|false||primary carenull|Primary Health Care|Procedure|false|false||primary carenull|True primary (qualifier value)|Time|false|false||primarynull|Primary|Modifier|false|false||primarynull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Pain in limb, lower leg|Finding|false|false||lower leg pain
null|Pain in lower limb|Finding|false|false||lower leg painnull|Lower extremity>Lower leg|Anatomy|false|false||lower leg
null|Leg|Anatomy|false|false||lower legnull|Body Site Modifier - Lower|Anatomy|false|false||lowernull|Lower (action)|Event|false|false||lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Pain in lower limb|Finding|false|false||leg painnull|Lower Extremity|Anatomy|false|false||leg
null|Leg|Anatomy|false|false||legnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Talking With Your Doctor|Finding|false|false||talk to your doctornull|Does talk|Finding|false|false||talk
null|Speech|Finding|false|false||talk
null|Speaking (function)|Finding|false|false||talknull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Spine Problem|Finding|false|false||spinenull|Neuron spine|Anatomy|false|false||spine
null|Vertebral column|Anatomy|false|false||spinenull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|diclofenac|Drug|false|false||DICLOFENAC
null|diclofenac|Drug|false|false||DICLOFENACnull|Gel - ContainerSeparator|Drug|false|false||GEL
null|Electrophoresis Gel|Drug|false|false||GEL
null|Gel|Drug|false|false||GEL
null|Gel physical state|Drug|false|false||GELnull|Blood group antibody screen.GEL|Procedure|false|false||GELnull|Voltaren|Drug|false|false||VOLTAREN
null|Voltaren|Drug|false|false||VOLTARENnull|Motrin|Drug|false|false||Motrin
null|Motrin|Drug|false|false||Motrinnull|Advil|Drug|false|false||Advil
null|Advil|Drug|false|false||Advilnull|AVIL gene|Finding|false|false||Advilnull|Topical Dosage Form|Drug|false|false||topicalnull|Topical Route of Administration|Finding|false|false||topicalnull|Topical surface|Modifier|false|false||topicalnull|Formation|Finding|false|false||formnull|null|Attribute|false|false||formnull|Manufactured form|Device|false|false||formnull|Qualitative form|Modifier|false|false||formnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Iron Drug Class|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|iron|Drug|false|false||iron
null|Ferrum metallicum, Homeopathic preparation|Drug|false|false||ironnull|Iron measurement|Procedure|false|false||ironnull|Deficiency|Finding|false|false||deficientnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|Role Class - part|Finding|false|false||partnull|Part|Modifier|false|false||partnull|Part Dosing Unit|LabModifier|false|false||partnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Vitelliform Macular Dystrophy|Disorder|false|false||bestnull|BEST1 wt Allele|Finding|false|false||best
null|BEST1 gene|Finding|false|false||bestnull|best (quality)|Modifier|false|false||bestnull|Health|Finding|false|false||healthnull|Team|Subject|false|false||teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions