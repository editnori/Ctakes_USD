 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|30,34
No|35,37
:|37,38
_|41,42
_|42,43
_|43,44
<EOL>|44,45
<EOL>|46,47
Admission|47,56
Date|57,61
:|61,62
_|64,65
_|65,66
_|66,67
Discharge|81,90
Date|91,95
:|95,96
_|99,100
_|100,101
_|101,102
<EOL>|102,103
<EOL>|104,105
Date|105,109
of|110,112
Birth|113,118
:|118,119
_|121,122
_|122,123
_|123,124
Sex|137,140
:|140,141
M|144,145
<EOL>|145,146
<EOL>|147,148
Service|148,155
:|155,156
MEDICINE|157,165
<EOL>|165,166
<EOL>|167,168
No|180,182
Known|183,188
Allergies|189,198
/|199,200
Adverse|201,208
Drug|209,213
Reactions|214,223
<EOL>|223,224
<EOL>|225,226
Attending|226,235
:|235,236
_|237,238
_|238,239
_|239,240
.|240,241
<EOL>|241,242
<EOL>|243,244
cardiogenic|261,272
_|273,274
_|274,275
_|275,276
,|276,277
NSTEMI|278,284
<EOL>|284,285
<EOL>|286,287
Major|287,292
Surgical|293,301
or|302,304
Invasive|305,313
Procedure|314,323
:|323,324
<EOL>|324,325
-|325,326
cardiac|327,334
catheterization|335,350
with|351,355
DES|356,359
to|360,362
mid-LAD|363,370
occlusion|371,380
via|381,384
R|385,386
<EOL>|387,388
radial|388,394
access|395,401
<EOL>|401,402
-|402,403
IABP|404,408
placement|409,418
and|419,422
removal|423,430
<EOL>|430,431
<EOL>|432,433
Mr.|461,464
_|465,466
_|466,467
_|467,468
is|469,471
a|472,473
_|474,475
_|475,476
_|476,477
M|478,479
with|480,484
HTN|485,488
,|488,489
HLD|490,493
,|493,494
DMII|495,499
,|499,500
and|501,504
prior|505,510
MI|511,513
with|514,518
<EOL>|519,520
medical|520,527
management|528,538
w|539,540
/|540,541
o|541,542
cath|543,547
presented|548,557
to|558,560
_|561,562
_|562,563
_|563,564
with|565,569
_|570,571
_|571,572
_|572,573
<EOL>|574,575
transferred|575,586
to|587,589
_|590,591
_|591,592
_|592,593
for|594,597
catheterization|598,613
for|614,617
concern|618,625
for|626,629
STEMI|630,635
.|635,636
<EOL>|637,638
<EOL>|638,639
Patient|639,646
has|647,650
long|651,655
standing|656,664
angina|665,671
pain|672,676
w|677,678
/|678,679
exertion|680,688
.|688,689
On|690,692
_|693,694
_|694,695
_|695,696
night|697,702
<EOL>|703,704
had|704,707
acute|708,713
onset|714,719
b|720,721
/|721,722
l|722,723
non-radiating|724,737
_|738,739
_|739,740
_|740,741
CP|742,744
not|745,748
resolved|749,757
with|758,762
SL|763,765
<EOL>|766,767
NTG|767,770
that|771,775
persisted|776,785
on|786,788
_|789,790
_|790,791
_|791,792
morning|793,800
.|800,801
In|802,804
addition|805,813
had|814,817
3|818,819
episodes|820,828
<EOL>|829,830
of|830,832
diarrhea|833,841
and|842,845
weakness|846,854
/|854,855
malaise|855,862
so|863,865
he|866,868
went|869,873
to|874,876
_|877,878
_|878,879
_|879,880
.|880,881
No|882,884
<EOL>|885,886
orthopnea|886,895
,|895,896
PND|897,900
,|900,901
_|902,903
_|903,904
_|904,905
edema|906,911
,|911,912
palpitations|913,925
,|925,926
or|927,929
SOB|930,933
.|933,934
<EOL>|935,936
<EOL>|936,937
In|937,939
the|940,943
ED|944,946
,|946,947
initial|948,955
vitals|956,962
were|963,967
:|967,968
<EOL>|970,971
Exam|971,975
:|975,976
Chest|977,982
pain|983,987
_|988,989
_|989,990
_|990,991
nonradiating|992,1004
<EOL>|1004,1005
Labs|1005,1009
:|1009,1010
Trop|1011,1015
I|1016,1017
1.14|1018,1022
,|1022,1023
WBC|1024,1027
29.6|1028,1032
,|1032,1033
Hct|1034,1037
38.7|1038,1042
,|1042,1043
Plt|1044,1047
148|1048,1051
,|1051,1052
INR|1053,1056
1.25|1057,1061
,|1061,1062
Na|1063,1065
<EOL>|1066,1067
127|1067,1070
,|1070,1071
K|1072,1073
+|1073,1074
4.6|1075,1078
,|1078,1079
BUN|1080,1083
30|1084,1086
/|1086,1087
Cr1|1087,1090
.|1090,1091
86|1091,1093
<EOL>|1093,1094
Imaging|1094,1101
:|1101,1102
EKG|1103,1106
showed|1107,1113
ST|1114,1116
elevations|1117,1127
in|1128,1130
AVR|1131,1134
(|1135,1136
2mm|1136,1139
)|1139,1140
,|1140,1141
borderline|1142,1152
<EOL>|1153,1154
elevation|1154,1163
in|1164,1166
V1|1167,1169
,|1169,1170
and|1171,1174
otherwise|1175,1184
diffuse|1185,1192
ST|1193,1195
depressions|1196,1207
.|1207,1208
Bedside|1209,1216
<EOL>|1217,1218
ECHO|1218,1222
w|1223,1224
/|1224,1225
septal|1226,1232
wall|1233,1237
motion|1238,1244
abnormalities|1245,1258
.|1258,1259
CXR|1260,1263
w|1264,1265
/|1265,1266
o|1266,1267
any|1268,1271
acute|1272,1277
<EOL>|1278,1279
abnormalities|1279,1292
.|1292,1293
<EOL>|1294,1295
Patient|1295,1302
was|1303,1306
given|1307,1312
:|1312,1313
Heparin|1314,1321
gtt|1322,1325
,|1325,1326
Nitro|1327,1332
gtt|1333,1336
,|1336,1337
ASA|1338,1341
324mg|1342,1347
,|1347,1348
Ticagrelor|1349,1359
<EOL>|1360,1361
180mg|1361,1366
@|1367,1368
1500|1369,1373
,|1373,1374
Vanco|1375,1380
125mg|1381,1386
PO|1387,1389
,|1389,1390
_|1391,1392
_|1392,1393
_|1393,1394
<EOL>|1394,1395
<EOL>|1395,1396
Transferred|1396,1407
to|1408,1410
_|1411,1412
_|1412,1413
_|1413,1414
for|1415,1418
cardiac|1419,1426
cath|1427,1431
.|1431,1432
Vitals|1433,1439
on|1440,1442
transfer|1443,1451
were|1452,1456
:|1456,1457
<EOL>|1458,1459
106|1459,1462
/|1462,1463
64|1463,1465
,|1465,1466
86|1467,1469
,|1469,1470
100|1471,1474
%|1474,1475
on|1476,1478
2L|1479,1481
,|1481,1482
afebrile|1483,1491
<EOL>|1491,1492
Cath|1492,1496
lab|1497,1500
where|1501,1506
he|1507,1509
still|1510,1515
had|1516,1519
_|1520,1521
_|1521,1522
_|1522,1523
pain|1524,1528
on|1529,1531
heparin|1532,1539
and|1540,1543
nitro|1544,1549
gtt|1550,1553
.|1553,1554
<EOL>|1555,1556
Catheterization|1556,1571
showed|1572,1578
mid-LAD|1579,1586
septal|1587,1593
occlusion|1594,1603
,|1603,1604
diffuse|1605,1612
disease|1613,1620
<EOL>|1621,1622
throughout|1622,1632
RCA|1633,1636
,|1636,1637
complete|1638,1646
occlusion|1647,1656
of|1657,1659
circumflex|1660,1670
w|1671,1672
/|1672,1673
collaterals|1674,1685
,|1685,1686
<EOL>|1687,1688
and|1688,1691
20|1692,1694
%|1694,1695
stenosis|1696,1704
of|1705,1707
L|1708,1709
main|1710,1714
.|1714,1715
DES|1716,1719
to|1720,1722
mid-LAD|1723,1730
occlusion|1731,1740
via|1741,1744
R|1745,1746
<EOL>|1747,1748
radial|1748,1754
access|1755,1761
.|1761,1762
Hypotensive|1763,1774
throughout|1775,1785
so|1786,1788
given|1789,1794
750cc|1795,1800
IVF|1801,1804
.|1804,1805
<EOL>|1806,1807
Coughing|1807,1815
post-procedure|1816,1830
with|1831,1835
LVEDP|1836,1841
25|1842,1844
so|1845,1847
given|1848,1853
Lasix|1854,1859
20mg|1860,1864
IV|1865,1867
.|1867,1868
<EOL>|1869,1870
Was|1870,1873
then|1874,1878
hypertensive|1879,1891
to|1892,1894
150|1895,1898
so|1899,1901
given|1902,1907
further|1908,1915
Lasix|1916,1921
40mg|1922,1926
IV|1927,1929
.|1929,1930
<EOL>|1930,1931
<EOL>|1931,1932
Admitted|1932,1940
to|1941,1943
CCU|1944,1947
for|1948,1951
hypotension|1952,1963
throughout|1964,1974
procedure|1975,1984
,|1984,1985
WBC|1986,1989
30|1990,1992
,|1992,1993
<EOL>|1994,1995
and|1995,1998
lack|1999,2003
of|2004,2006
_|2007,2008
_|2008,2009
_|2009,2010
beds|2011,2015
.|2015,2016
In|2017,2019
the|2020,2023
CCU|2024,2027
,|2027,2028
patient|2029,2036
reports|2037,2044
no|2045,2047
chest|2048,2053
pain|2054,2058
<EOL>|2059,2060
but|2060,2063
continues|2064,2073
to|2074,2076
have|2077,2081
productive|2082,2092
cough|2093,2098
and|2099,2102
diarrhea|2103,2111
.|2111,2112
<EOL>|2112,2113
<EOL>|2113,2114
Of|2114,2116
note|2117,2121
,|2121,2122
two|2123,2126
weeks|2127,2132
ago|2133,2136
had|2137,2140
endoscopy|2141,2150
and|2151,2154
diagnosed|2155,2164
with|2165,2169
H|2170,2171
<EOL>|2172,2173
Pylori|2173,2179
.|2179,2180
Currently|2181,2190
on|2191,2193
clarithromycin|2194,2208
and|2209,2212
amoxicillin|2213,2224
.|2224,2225
On|2226,2228
_|2229,2230
_|2230,2231
_|2231,2232
<EOL>|2233,2234
night|2234,2239
developed|2240,2249
diarrhea|2250,2258
.|2258,2259
Also|2260,2264
had|2265,2268
15lb|2269,2273
weight|2274,2280
loss|2281,2285
in|2286,2288
past|2289,2293
4|2294,2295
<EOL>|2296,2297
months|2297,2303
.|2303,2304
<EOL>|2304,2305
<EOL>|2305,2306
<EOL>|2307,2308
1|2330,2331
)|2331,2332
HTN|2333,2336
<EOL>|2336,2337
2|2337,2338
)|2338,2339
HLD|2340,2343
<EOL>|2343,2344
3|2344,2345
)|2345,2346
DMII|2347,2351
<EOL>|2351,2352
4|2352,2353
)|2353,2354
CAD|2355,2358
s|2359,2360
/|2360,2361
p|2361,2362
MI|2363,2365
-|2366,2367
medically|2368,2377
managed|2378,2385
<EOL>|2385,2386
5|2386,2387
)|2387,2388
H.|2389,2391
Pylori|2392,2398
<EOL>|2398,2399
6|2399,2400
)|2400,2401
Spinal|2402,2408
stenosis|2409,2417
<EOL>|2417,2418
<EOL>|2419,2420
:|2434,2435
<EOL>|2435,2436
_|2436,2437
_|2437,2438
_|2438,2439
<EOL>|2439,2440
:|2454,2455
<EOL>|2455,2456
Father|2456,2462
:|2462,2463
possible|2464,2472
dilated|2473,2480
cardiomyopathy|2481,2495
<EOL>|2495,2496
No|2496,2498
family|2499,2505
history|2506,2513
of|2514,2516
early|2517,2522
MI|2523,2525
,|2525,2526
arrhythmia|2527,2537
,|2537,2538
or|2539,2541
sudden|2542,2548
cardiac|2549,2556
<EOL>|2557,2558
death|2558,2563
;|2563,2564
otherwise|2565,2574
non-contributory|2575,2591
.|2591,2592
<EOL>|2594,2595
<EOL>|2596,2597
On|2612,2614
admission|2615,2624
:|2624,2625
<EOL>|2625,2626
-|2626,2627
-|2627,2628
-|2628,2629
-|2629,2630
-|2630,2631
-|2631,2632
-|2632,2633
-|2633,2634
-|2634,2635
-|2635,2636
-|2636,2637
-|2637,2638
-|2638,2639
-|2639,2640
-|2640,2641
<EOL>|2641,2642
VS|2642,2644
:|2644,2645
afebrile|2646,2654
,|2654,2655
160|2656,2659
/|2659,2660
80|2660,2662
,|2662,2663
114|2664,2667
,|2667,2668
94|2669,2671
%|2671,2672
on|2673,2675
15L|2676,2679
Non-rebreather|2680,2694
<EOL>|2694,2695
Weight|2695,2701
:|2701,2702
69kg|2703,2707
<EOL>|2707,2708
Tele|2708,2712
:|2712,2713
NSR|2714,2717
<EOL>|2717,2718
Gen|2718,2721
:|2721,2722
Slightly|2723,2731
tachypneic|2732,2742
older|2743,2748
man|2749,2752
audibly|2753,2760
wheezing|2761,2769
but|2770,2773
<EOL>|2774,2775
comfortably|2775,2786
finishing|2787,2796
sentences|2797,2806
<EOL>|2807,2808
HEENT|2808,2813
:|2813,2814
EOMI|2815,2819
,|2819,2820
PERRLA|2821,2827
,|2827,2828
<EOL>|2828,2829
NECK|2829,2833
:|2833,2834
No|2835,2837
JVD|2838,2841
<EOL>|2841,2842
CV|2842,2844
:|2844,2845
Tachycardic|2846,2857
,|2857,2858
difficult|2859,2868
to|2869,2871
appreciate|2872,2882
heart|2883,2888
sounds|2889,2895
due|2896,2899
to|2900,2902
<EOL>|2903,2904
significant|2904,2915
rhonchi|2916,2923
<EOL>|2924,2925
LUNGS|2925,2930
:|2930,2931
b|2932,2933
/|2933,2934
l|2934,2935
rhonchi|2936,2943
throughout|2944,2954
w|2955,2956
/|2956,2957
mild|2958,2962
end|2963,2966
expiratory|2967,2977
wheezing|2978,2986
<EOL>|2987,2988
and|2988,2991
R|2992,2993
base|2994,2998
crackles|2999,3007
<EOL>|3007,3008
ABD|3008,3011
:|3011,3012
Soft|3013,3017
,|3017,3018
Non-tender|3019,3029
,|3029,3030
non-distended|3031,3044
<EOL>|3044,3045
EXT|3045,3048
:|3048,3049
2|3050,3051
+|3051,3052
L|3053,3054
radial|3055,3061
pulses|3062,3068
,|3068,3069
R|3070,3071
arm|3072,3075
w|3076,3077
/|3077,3078
band|3079,3083
in|3084,3086
place|3087,3092
and|3093,3096
normal|3097,3103
<EOL>|3104,3105
motor|3105,3110
/|3110,3111
sensory|3111,3118
function|3119,3127
intact|3128,3134
distally|3135,3143
,|3143,3144
RLE|3145,3148
non-palpable|3149,3161
DP|3162,3164
but|3165,3168
<EOL>|3169,3170
dopplerable|3170,3181
,|3181,3182
1|3183,3184
+|3184,3185
LLE|3186,3189
DP.|3190,3193
b|3194,3195
/|3195,3196
l|3196,3197
_|3198,3199
_|3199,3200
_|3200,3201
slightly|3202,3210
cold|3211,3215
but|3216,3219
normal|3220,3226
<EOL>|3227,3228
sensation|3228,3237
w|3238,3239
/|3239,3240
full|3241,3245
motor|3246,3251
strength|3252,3260
and|3261,3264
ROM|3265,3268
<EOL>|3268,3269
SKIN|3269,3273
:|3273,3274
No|3275,3277
rashes|3278,3284
or|3285,3287
chronic|3288,3295
edematous|3296,3305
changes|3306,3313
<EOL>|3313,3314
NEURO|3314,3319
:|3319,3320
Alert|3321,3326
and|3327,3330
attentive|3331,3340
,|3340,3341
AOX3|3342,3346
,|3346,3347
Moving|3348,3354
all|3355,3358
extremities|3359,3370
<EOL>|3370,3371
<EOL>|3371,3372
At|3372,3374
discharge|3375,3384
:|3384,3385
<EOL>|3385,3386
-|3386,3387
-|3387,3388
-|3388,3389
-|3389,3390
-|3390,3391
-|3391,3392
-|3392,3393
-|3393,3394
-|3394,3395
-|3395,3396
-|3396,3397
-|3397,3398
-|3398,3399
-|3399,3400
<EOL>|3400,3401
Weight|3401,3407
:|3407,3408
63.7|3410,3414
kg|3414,3416
(|3417,3418
63.4|3418,3422
)|3422,3423
<EOL>|3424,3425
I|3425,3426
/|3426,3427
O|3427,3428
:|3428,3429
980|3430,3433
/|3433,3434
800|3434,3437
<EOL>|3437,3438
T|3438,3439
98.4|3440,3444
BP|3445,3447
123|3448,3451
/|3451,3452
68|3452,3454
(|3455,3456
102|3456,3459
-|3459,3460
133|3460,3463
/|3463,3464
62|3464,3466
-|3466,3467
87|3467,3469
)|3469,3470
P|3471,3472
86|3473,3475
(|3476,3477
71|3477,3479
-|3479,3480
100|3480,3483
)|3483,3484
RR|3485,3487
20|3488,3490
O2|3491,3493
99|3494,3496
%|3496,3497
RA|3498,3500
<EOL>|3503,3504
<EOL>|3505,3506
Gen|3506,3509
:|3509,3510
awake|3511,3516
,|3516,3517
alert|3518,3523
,|3523,3524
oriented|3525,3533
to|3534,3536
self|3537,3541
,|3541,3542
date|3543,3547
,|3547,3548
hospital|3549,3557
<EOL>|3557,3558
HEENT|3558,3563
:|3563,3564
EOMI|3565,3569
,|3569,3570
PERRLA|3571,3577
,|3577,3578
<EOL>|3578,3579
NECK|3579,3583
:|3583,3584
No|3585,3587
JVD|3588,3591
<EOL>|3591,3592
CV|3592,3594
:|3594,3595
Tachycardic|3596,3607
,|3607,3608
difficult|3609,3618
to|3619,3621
appreciate|3622,3632
heart|3633,3638
sounds|3639,3645
<EOL>|3646,3647
LUNGS|3647,3652
:|3652,3653
Bibasilar|3655,3664
crackles|3665,3673
<EOL>|3673,3674
ABD|3674,3677
:|3677,3678
Soft|3679,3683
,|3683,3684
Non-tender|3685,3695
,|3695,3696
non-distended|3697,3710
<EOL>|3710,3711
EXT|3711,3714
:|3714,3715
2|3716,3717
+|3717,3718
b|3719,3720
/|3720,3721
l|3721,3722
radial|3723,3729
pulses|3730,3736
,|3736,3737
R|3738,3739
arm|3740,3743
normal|3745,3751
motor|3752,3757
/|3757,3758
sensory|3758,3765
function|3766,3774
<EOL>|3775,3776
intact|3776,3782
distally|3783,3791
,|3791,3792
RLE|3793,3796
non-palpable|3797,3809
DP|3810,3812
but|3813,3816
dopplerable|3817,3828
,|3828,3829
trace|3830,3835
<EOL>|3836,3837
edema|3837,3842
b|3843,3844
/|3844,3845
l|3845,3846
.|3846,3847
b|3848,3849
/|3849,3850
l|3850,3851
_|3852,3853
_|3853,3854
_|3854,3855
slightly|3856,3864
cold|3865,3869
but|3870,3873
normal|3874,3880
sensation|3881,3890
w|3891,3892
/|3892,3893
full|3894,3898
<EOL>|3899,3900
motor|3900,3905
strength|3906,3914
and|3915,3918
ROM|3919,3922
<EOL>|3922,3923
SKIN|3923,3927
:|3927,3928
No|3929,3931
rashes|3932,3938
or|3939,3941
chronic|3942,3949
edematous|3950,3959
changes|3960,3967
<EOL>|3967,3968
NEURO|3968,3973
:|3973,3974
Alert|3975,3980
and|3981,3984
attentive|3985,3994
,|3994,3995
AOX3|3996,4000
,|4000,4001
Moving|4002,4008
all|4009,4012
extremities|4013,4024
<EOL>|4024,4025
<EOL>|4025,4026
<EOL>|4027,4028
Pertinent|4028,4037
Results|4038,4045
:|4045,4046
<EOL>|4046,4047
Labs|4047,4051
on|4052,4054
Admission|4055,4064
:|4064,4065
<EOL>|4065,4066
-|4066,4067
-|4067,4068
-|4068,4069
-|4069,4070
-|4070,4071
-|4071,4072
-|4072,4073
-|4073,4074
-|4074,4075
-|4075,4076
-|4076,4077
-|4077,4078
-|4078,4079
-|4079,4080
-|4080,4081
-|4081,4082
-|4082,4083
-|4083,4084
-|4084,4085
<EOL>|4085,4086
_|4086,4087
_|4087,4088
_|4088,4089
09|4090,4092
:|4092,4093
23PM|4093,4097
WBC|4100,4103
-|4103,4104
36|4104,4106
.|4106,4107
8|4107,4108
*|4108,4109
RBC|4110,4113
-|4113,4114
4|4114,4115
.|4115,4116
40|4116,4118
*|4118,4119
HGB|4120,4123
-|4123,4124
14.0|4124,4128
HCT|4129,4132
-|4132,4133
40.6|4133,4137
MCV|4138,4141
-|4141,4142
92|4142,4144
<EOL>|4145,4146
MCH|4146,4149
-|4149,4150
31.8|4150,4154
MCHC|4155,4159
-|4159,4160
34.5|4160,4164
RDW|4165,4168
-|4168,4169
12.5|4169,4173
RDWSD|4174,4179
-|4179,4180
41.8|4180,4184
<EOL>|4184,4185
_|4185,4186
_|4186,4187
_|4187,4188
09|4189,4191
:|4191,4192
23PM|4192,4196
PLT|4199,4202
SMR|4203,4206
-|4206,4207
NORMAL|4207,4213
PLT|4214,4217
COUNT|4218,4223
-|4223,4224
176|4224,4227
<EOL>|4227,4228
_|4228,4229
_|4229,4230
_|4230,4231
09|4232,4234
:|4234,4235
23PM|4235,4239
NEUTS|4242,4247
-|4247,4248
81|4248,4250
*|4250,4251
BANDS|4252,4257
-|4257,4258
10|4258,4260
*|4260,4261
LYMPHS|4262,4268
-|4268,4269
3|4269,4270
*|4270,4271
MONOS|4272,4277
-|4277,4278
6|4278,4279
EOS|4280,4283
-|4283,4284
0|4284,4285
<EOL>|4286,4287
BASOS|4287,4292
-|4292,4293
0|4293,4294
_|4295,4296
_|4296,4297
_|4297,4298
MYELOS|4299,4305
-|4305,4306
0|4306,4307
AbsNeut|4308,4315
-|4315,4316
33|4316,4318
.|4318,4319
49|4319,4321
*|4321,4322
AbsLymp|4323,4330
-|4330,4331
1|4331,4332
.|4332,4333
10|4333,4335
*|4335,4336
<EOL>|4337,4338
AbsMono|4338,4345
-|4345,4346
2|4346,4347
.|4347,4348
21|4348,4350
*|4350,4351
AbsEos|4352,4358
-|4358,4359
0|4359,4360
.|4360,4361
00|4361,4363
*|4363,4364
AbsBaso|4365,4372
-|4372,4373
0|4373,4374
.|4374,4375
00|4375,4377
*|4377,4378
<EOL>|4378,4379
_|4379,4380
_|4380,4381
_|4381,4382
09|4383,4385
:|4385,4386
23PM|4386,4390
_|4393,4394
_|4394,4395
_|4395,4396
PTT|4397,4400
-|4400,4401
49|4401,4403
.|4403,4404
6|4404,4405
*|4405,4406
_|4407,4408
_|4408,4409
_|4409,4410
<EOL>|4410,4411
_|4411,4412
_|4412,4413
_|4413,4414
09|4415,4417
:|4417,4418
23PM|4418,4422
GLUCOSE|4425,4432
-|4432,4433
264|4433,4436
*|4436,4437
UREA|4438,4442
N|4443,4444
-|4444,4445
30|4445,4447
*|4447,4448
CREAT|4449,4454
-|4454,4455
1|4455,4456
.|4456,4457
4|4457,4458
*|4458,4459
<EOL>|4460,4461
SODIUM|4461,4467
-|4467,4468
129|4468,4471
*|4471,4472
POTASSIUM|4473,4482
-|4482,4483
4.1|4483,4486
CHLORIDE|4487,4495
-|4495,4496
96|4496,4498
TOTAL|4499,4504
CO2|4505,4508
-|4508,4509
14|4509,4511
*|4511,4512
ANION|4513,4518
<EOL>|4519,4520
GAP|4520,4523
-|4523,4524
23|4524,4526
*|4526,4527
<EOL>|4527,4528
_|4528,4529
_|4529,4530
_|4530,4531
09|4532,4534
:|4534,4535
23PM|4535,4539
CALCIUM|4542,4549
-|4549,4550
8|4550,4551
.|4551,4552
2|4552,4553
*|4553,4554
PHOSPHATE|4555,4564
-|4564,4565
3.0|4565,4568
MAGNESIUM|4569,4578
-|4578,4579
1.7|4579,4582
<EOL>|4583,4584
CHOLEST|4584,4591
-|4591,4592
157|4592,4595
<EOL>|4595,4596
_|4596,4597
_|4597,4598
_|4598,4599
09|4600,4602
:|4602,4603
23PM|4603,4607
%|4610,4611
HbA1c|4611,4616
-|4616,4617
5.9|4617,4620
eAG|4621,4624
-|4624,4625
123|4625,4628
<EOL>|4628,4629
_|4629,4630
_|4630,4631
_|4631,4632
09|4633,4635
:|4635,4636
23PM|4636,4640
CK|4643,4645
-|4645,4646
MB|4646,4648
-|4648,4649
44|4649,4651
*|4651,4652
cTropnT|4653,4660
-|4660,4661
0|4661,4662
.|4662,4663
69|4663,4665
*|4665,4666
<EOL>|4666,4667
_|4667,4668
_|4668,4669
_|4669,4670
09|4671,4673
:|4673,4674
23PM|4674,4678
TRIGLYCER|4681,4690
-|4690,4691
90|4691,4693
HDL|4694,4697
CHOL|4698,4702
-|4702,4703
42|4703,4705
CHOL|4706,4710
/|4710,4711
HDL|4711,4714
-|4714,4715
3.7|4715,4718
<EOL>|4719,4720
LDL|4720,4723
(|4723,4724
CALC|4724,4728
)|4728,4729
-|4729,4730
97|4730,4732
<EOL>|4732,4733
_|4733,4734
_|4734,4735
_|4735,4736
09|4737,4739
:|4739,4740
23PM|4740,4744
HYPOCHROM|4747,4756
-|4756,4757
NORMAL|4757,4763
ANISOCYT|4764,4772
-|4772,4773
NORMAL|4773,4779
POIKILOCY|4780,4789
-|4789,4790
1|4790,4791
+|4791,4792
<EOL>|4793,4794
MACROCYT|4794,4802
-|4802,4803
NORMAL|4803,4809
MICROCYT|4810,4818
-|4818,4819
NORMAL|4819,4825
POLYCHROM|4826,4835
-|4835,4836
NORMAL|4836,4842
BURR|4843,4847
-|4847,4848
1|4848,4849
+|4849,4850
<EOL>|4850,4851
<EOL>|4851,4852
Labs|4852,4856
at|4857,4859
Discharge|4860,4869
:|4869,4870
<EOL>|4870,4871
-|4871,4872
-|4872,4873
-|4873,4874
-|4874,4875
-|4875,4876
-|4876,4877
-|4877,4878
-|4878,4879
-|4879,4880
-|4880,4881
-|4881,4882
-|4882,4883
-|4883,4884
-|4884,4885
-|4885,4886
-|4886,4887
-|4887,4888
-|4888,4889
-|4889,4890
<EOL>|4890,4891
_|4891,4892
_|4892,4893
_|4893,4894
05|4895,4897
:|4897,4898
50AM|4898,4902
BLOOD|4903,4908
WBC|4909,4912
-|4912,4913
11|4913,4915
.|4915,4916
2|4916,4917
*|4917,4918
RBC|4919,4922
-|4922,4923
3|4923,4924
.|4924,4925
59|4925,4927
*|4927,4928
Hgb|4929,4932
-|4932,4933
11|4933,4935
.|4935,4936
2|4936,4937
*|4937,4938
Hct|4939,4942
-|4942,4943
34|4943,4945
.|4945,4946
7|4946,4947
*|4947,4948
<EOL>|4949,4950
MCV|4950,4953
-|4953,4954
97|4954,4956
MCH|4957,4960
-|4960,4961
31.2|4961,4965
MCHC|4966,4970
-|4970,4971
32.3|4971,4975
RDW|4976,4979
-|4979,4980
13.2|4980,4984
RDWSD|4985,4990
-|4990,4991
46|4991,4993
.|4993,4994
7|4994,4995
*|4995,4996
Plt|4997,5000
_|5001,5002
_|5002,5003
_|5003,5004
<EOL>|5004,5005
_|5005,5006
_|5006,5007
_|5007,5008
05|5009,5011
:|5011,5012
50AM|5012,5016
BLOOD|5017,5022
Neuts|5023,5028
-|5028,5029
76|5029,5031
*|5031,5032
Bands|5033,5038
-|5038,5039
0|5039,5040
Lymphs|5041,5047
-|5047,5048
16|5048,5050
*|5050,5051
Monos|5052,5057
-|5057,5058
5|5058,5059
<EOL>|5060,5061
Eos|5061,5064
-|5064,5065
2|5065,5066
Baso|5067,5071
-|5071,5072
0|5072,5073
_|5074,5075
_|5075,5076
_|5076,5077
Metas|5078,5083
-|5083,5084
1|5084,5085
*|5085,5086
Myelos|5087,5093
-|5093,5094
0|5094,5095
AbsNeut|5096,5103
-|5103,5104
8|5104,5105
.|5105,5106
51|5106,5108
*|5108,5109
<EOL>|5110,5111
AbsLymp|5111,5118
-|5118,5119
1|5119,5120
.|5120,5121
79|5121,5123
AbsMono|5124,5131
-|5131,5132
0|5132,5133
.|5133,5134
56|5134,5136
AbsEos|5137,5143
-|5143,5144
0|5144,5145
.|5145,5146
22|5146,5148
AbsBaso|5149,5156
-|5156,5157
0|5157,5158
.|5158,5159
00|5159,5161
*|5161,5162
<EOL>|5162,5163
_|5163,5164
_|5164,5165
_|5165,5166
05|5167,5169
:|5169,5170
50AM|5170,5174
BLOOD|5175,5180
_|5181,5182
_|5182,5183
_|5183,5184
PTT|5185,5188
-|5188,5189
27.3|5189,5193
_|5194,5195
_|5195,5196
_|5196,5197
<EOL>|5197,5198
_|5198,5199
_|5199,5200
_|5200,5201
05|5202,5204
:|5204,5205
50AM|5205,5209
BLOOD|5210,5215
Glucose|5216,5223
-|5223,5224
165|5224,5227
*|5227,5228
UreaN|5229,5234
-|5234,5235
43|5235,5237
*|5237,5238
Creat|5239,5244
-|5244,5245
1.1|5245,5248
Na|5249,5251
-|5251,5252
136|5252,5255
<EOL>|5256,5257
K|5257,5258
-|5258,5259
4.3|5259,5262
Cl|5263,5265
-|5265,5266
103|5266,5269
HCO3|5270,5274
-|5274,5275
22|5275,5277
AnGap|5278,5283
-|5283,5284
15|5284,5286
<EOL>|5286,5287
_|5287,5288
_|5288,5289
_|5289,5290
05|5291,5293
:|5293,5294
50AM|5294,5298
BLOOD|5299,5304
ALT|5305,5308
-|5308,5309
38|5309,5311
AST|5312,5315
-|5315,5316
32|5316,5318
LD|5319,5321
(|5321,5322
LDH|5322,5325
)|5325,5326
-|5326,5327
481|5327,5330
*|5330,5331
AlkPhos|5332,5339
-|5339,5340
99|5340,5342
<EOL>|5343,5344
TotBili|5344,5351
-|5351,5352
0.4|5352,5355
<EOL>|5355,5356
_|5356,5357
_|5357,5358
_|5358,5359
05|5360,5362
:|5362,5363
50AM|5363,5367
BLOOD|5368,5373
Albumin|5374,5381
-|5381,5382
3|5382,5383
.|5383,5384
3|5384,5385
*|5385,5386
Calcium|5387,5394
-|5394,5395
8.4|5395,5398
Phos|5399,5403
-|5403,5404
3.6|5404,5407
Mg|5408,5410
-|5410,5411
2.4|5411,5414
<EOL>|5414,5415
<EOL>|5415,5416
Relevant|5416,5424
Imaging|5425,5432
:|5432,5433
<EOL>|5433,5434
-|5434,5435
-|5435,5436
-|5436,5437
-|5437,5438
-|5438,5439
-|5439,5440
-|5440,5441
-|5441,5442
-|5442,5443
-|5443,5444
-|5444,5445
-|5445,5446
-|5446,5447
-|5447,5448
-|5448,5449
-|5449,5450
-|5450,5451
<EOL>|5451,5452
TTE|5452,5455
_|5456,5457
_|5457,5458
_|5458,5459
:|5459,5460
<EOL>|5460,5461
The|5461,5464
left|5465,5469
atrium|5470,5476
is|5477,5479
mildly|5480,5486
dilated|5487,5494
.|5494,5495
The|5496,5499
estimated|5500,5509
right|5510,5515
atrial|5516,5522
<EOL>|5523,5524
pressure|5524,5532
is|5533,5535
_|5536,5537
_|5537,5538
_|5538,5539
mmHg|5540,5544
.|5544,5545
Left|5546,5550
ventricular|5551,5562
wall|5563,5567
thicknesses|5568,5579
and|5580,5583
<EOL>|5584,5585
cavity|5585,5591
size|5592,5596
are|5597,5600
normal|5601,5607
.|5607,5608
Overall|5609,5616
left|5617,5621
ventricular|5622,5633
systolic|5634,5642
<EOL>|5643,5644
function|5644,5652
is|5653,5655
moderately|5656,5666
depressed|5667,5676
(|5677,5678
LVEF|5678,5682
=|5682,5683
?|5684,5685
35|5686,5688
-|5688,5689
40|5689,5691
%|5691,5692
-|5693,5694
assessment|5695,5705
<EOL>|5706,5707
limited|5707,5714
by|5715,5717
suboptimal|5718,5728
image|5729,5734
quality|5735,5742
and|5743,5746
significant|5747,5758
beat|5759,5763
to|5764,5766
beat|5767,5771
<EOL>|5772,5773
variability|5773,5784
)|5784,5785
.|5785,5786
There|5787,5792
is|5793,5795
hypokinesis|5796,5807
of|5808,5810
the|5811,5814
mid-distal|5815,5825
LV|5826,5828
segments|5829,5837
<EOL>|5838,5839
and|5839,5842
apex|5843,5847
.|5847,5848
There|5849,5854
is|5855,5857
no|5858,5860
ventricular|5861,5872
septal|5873,5879
defect|5880,5886
.|5886,5887
Right|5888,5893
<EOL>|5894,5895
ventricular|5895,5906
chamber|5907,5914
size|5915,5919
and|5920,5923
free|5924,5928
wall|5929,5933
motion|5934,5940
are|5941,5944
normal|5945,5951
.|5951,5952
The|5953,5956
<EOL>|5957,5958
ascending|5958,5967
aorta|5968,5973
is|5974,5976
mildly|5977,5983
dilated|5984,5991
.|5991,5992
The|5993,5996
number|5997,6003
of|6004,6006
aortic|6007,6013
valve|6014,6019
<EOL>|6020,6021
leaflets|6021,6029
can|6030,6033
not|6033,6036
be|6037,6039
determined|6040,6050
.|6050,6051
There|6052,6057
is|6058,6060
mild|6061,6065
aortic|6066,6072
valve|6073,6078
<EOL>|6079,6080
stenosis|6080,6088
(|6089,6090
valve|6090,6095
area|6096,6100
1.2|6101,6104
-|6104,6105
1.9|6105,6108
cm2|6108,6111
)|6111,6112
.|6112,6113
No|6114,6116
aortic|6117,6123
regurgitation|6124,6137
is|6138,6140
<EOL>|6141,6142
seen|6142,6146
.|6146,6147
The|6148,6151
mitral|6152,6158
valve|6159,6164
appears|6165,6172
structurally|6173,6185
normal|6186,6192
with|6193,6197
trivial|6198,6205
<EOL>|6206,6207
mitral|6207,6213
regurgitation|6214,6227
.|6227,6228
The|6229,6232
pulmonary|6233,6242
artery|6243,6249
systolic|6250,6258
pressure|6259,6267
<EOL>|6268,6269
could|6269,6274
not|6275,6278
be|6279,6281
determined|6282,6292
.|6292,6293
There|6294,6299
is|6300,6302
a|6303,6304
trivial|6305,6312
/|6312,6313
physiologic|6313,6324
<EOL>|6325,6326
pericardial|6326,6337
effusion|6338,6346
.|6346,6347
<EOL>|6348,6349
<EOL>|6349,6350
Compared|6350,6358
with|6359,6363
the|6364,6367
prior|6368,6373
focused|6374,6381
study|6382,6387
(|6388,6389
images|6389,6395
reviewed|6396,6404
)|6404,6405
of|6406,6408
<EOL>|6409,6410
_|6410,6411
_|6411,6412
_|6412,6413
,|6413,6414
left|6415,6419
ventricular|6420,6431
systolic|6432,6440
function|6441,6449
is|6450,6452
probably|6453,6461
<EOL>|6462,6463
similar|6463,6470
,|6470,6471
although|6472,6480
suboptimal|6481,6491
image|6492,6497
quality|6498,6505
of|6506,6508
both|6509,6513
studies|6514,6521
<EOL>|6522,6523
precludes|6523,6532
definite|6533,6541
comparison|6542,6552
.|6552,6553
<EOL>|6555,6556
<EOL>|6556,6557
_|6557,6558
_|6558,6559
_|6559,6560
CXR|6561,6564
<EOL>|6564,6565
<EOL>|6566,6567
Generalized|6584,6595
improvement|6596,6607
in|6608,6610
both|6611,6615
lungs|6616,6621
is|6622,6624
probably|6625,6633
due|6634,6637
to|6638,6640
<EOL>|6641,6642
decrease|6642,6650
in|6651,6653
pulmonary|6654,6663
<EOL>|6664,6665
edema|6665,6670
,|6670,6671
now|6672,6675
mild|6676,6680
,|6680,6681
and|6682,6685
decrease|6686,6694
in|6695,6697
previous|6698,6706
moderate|6707,6715
right|6716,6721
pleural|6722,6729
<EOL>|6730,6731
effusion|6731,6739
.|6739,6740
<EOL>|6742,6743
There|6743,6748
is|6749,6751
still|6752,6757
substantial|6758,6769
consolidation|6770,6783
in|6784,6786
the|6787,6790
right|6791,6796
upper|6797,6802
lobe|6803,6807
<EOL>|6808,6809
probably|6809,6817
<EOL>|6818,6819
pneumonia|6819,6828
but|6829,6832
the|6833,6836
bilateral|6837,6846
lower|6847,6852
lobe|6853,6857
components|6858,6868
have|6869,6873
improved|6874,6882
.|6882,6883
<EOL>|6884,6885
Heart|6886,6891
size|6892,6896
<EOL>|6897,6898
top|6898,6901
-|6901,6902
normal|6902,6908
.|6908,6909
No|6911,6913
pneumothorax|6914,6926
.|6926,6927
<EOL>|6928,6929
<EOL>|6929,6930
MICRO|6930,6935
<EOL>|6935,6936
=|6936,6937
=|6937,6938
=|6938,6939
=|6939,6940
=|6940,6941
=|6941,6942
=|6942,6943
=|6943,6944
<EOL>|6944,6945
FINAL|6945,6950
REPORT|6951,6957
_|6958,6959
_|6959,6960
_|6960,6961
<EOL>|6961,6962
<EOL>|6962,6963
C.|6966,6968
difficile|6969,6978
DNA|6979,6982
amplification|6983,6996
assay|6997,7002
(|7003,7004
Final|7004,7009
_|7010,7011
_|7011,7012
_|7012,7013
:|7013,7014
<EOL>|7015,7016
CLOSTRIDIUM|7022,7033
DIFFICILE|7034,7043
.|7043,7044
<EOL>|7045,7046
Positive|7055,7063
for|7064,7067
toxigenic|7068,7077
C.|7078,7080
difficile|7081,7090
by|7091,7093
the|7094,7097
Illumigene|7098,7108
<EOL>|7109,7110
DNA|7110,7113
<EOL>|7113,7114
amplification|7123,7136
.|7136,7137
(|7149,7150
Reference|7150,7159
Range|7160,7165
-|7165,7166
Negative|7166,7174
)|7174,7175
.|7175,7176
<EOL>|7177,7178
<EOL>|7178,7179
_|7179,7180
_|7180,7181
_|7181,7182
12|7183,7185
:|7185,7186
53|7186,7188
pm|7189,7191
SPUTUM|7192,7198
Source|7204,7210
:|7210,7211
Expectorated|7212,7224
.|7224,7225
<EOL>|7226,7227
<EOL>|7227,7228
GRAM|7231,7235
STAIN|7236,7241
(|7242,7243
Final|7243,7248
_|7249,7250
_|7250,7251
_|7251,7252
:|7252,7253
<EOL>|7254,7255
<|7261,7262
10|7262,7264
PMNs|7265,7269
and|7270,7273
<|7274,7275
10|7275,7277
epithelial|7278,7288
cells|7289,7294
/|7294,7295
100X|7295,7299
field|7300,7305
.|7305,7306
<EOL>|7307,7308
2|7314,7315
+|7315,7316
_|7319,7320
_|7320,7321
_|7321,7322
per|7323,7326
1000X|7327,7332
FIELD|7333,7338
)|7338,7339
:|7339,7340
GRAM|7343,7347
NEGATIVE|7348,7356
ROD|7357,7360
(|7360,7361
S|7361,7362
)|7362,7363
.|7363,7364
<EOL>|7365,7366
2|7372,7373
+|7373,7374
_|7377,7378
_|7378,7379
_|7379,7380
per|7381,7384
1000X|7385,7390
FIELD|7391,7396
)|7396,7397
:|7397,7398
BUDDING|7401,7408
YEAST|7409,7414
.|7414,7415
<EOL>|7416,7417
QUALITY|7423,7430
OF|7431,7433
SPECIMEN|7434,7442
CAN|7443,7446
NOT|7446,7449
BE|7450,7452
ASSESSED|7453,7461
.|7461,7462
<EOL>|7463,7464
<EOL>|7464,7465
RESPIRATORY|7468,7479
CULTURE|7480,7487
(|7488,7489
Preliminary|7489,7500
)|7500,7501
:|7501,7502
<EOL>|7503,7504
Further|7510,7517
incubation|7518,7528
required|7529,7537
to|7538,7540
determine|7541,7550
the|7551,7554
presence|7555,7563
or|7564,7566
<EOL>|7567,7568
absence|7568,7575
of|7576,7578
<EOL>|7578,7579
commensal|7585,7594
respiratory|7595,7606
flora|7607,7612
.|7612,7613
<EOL>|7614,7615
KLEBSIELLA|7621,7631
PNEUMONIAE|7632,7642
.|7642,7643
SPARSE|7647,7653
GROWTH|7654,7660
.|7660,7661
<EOL>|7662,7663
Cefazolin|7672,7681
interpretative|7682,7696
criteria|7697,7705
are|7706,7709
based|7710,7715
on|7716,7718
a|7719,7720
dosage|7721,7727
<EOL>|7728,7729
regimen|7729,7736
of|7737,7739
<EOL>|7739,7740
2g|7749,7751
every|7752,7757
8h|7758,7760
.|7760,7761
<EOL>|7762,7763
GRAM|7769,7773
NEGATIVE|7774,7782
ROD|7783,7786
#|7787,7788
2.|7788,7790
SPARSE|7794,7800
GROWTH|7801,7807
.|7807,7808
<EOL>|7809,7810
<EOL>|7810,7811
SENSITIVITIES|7841,7854
:|7854,7855
MIC|7856,7859
expressed|7860,7869
in|7870,7872
<EOL>|7873,7874
MCG|7874,7877
/|7877,7878
ML|7878,7880
<EOL>|7880,7881
<EOL>|7903,7904
_|7904,7905
_|7905,7906
_|7906,7907
_|7907,7908
_|7908,7909
_|7909,7910
_|7910,7911
_|7911,7912
_|7912,7913
_|7913,7914
_|7914,7915
_|7915,7916
_|7916,7917
_|7917,7918
_|7918,7919
_|7919,7920
_|7920,7921
_|7921,7922
_|7922,7923
_|7923,7924
_|7924,7925
_|7925,7926
_|7926,7927
_|7927,7928
_|7928,7929
_|7929,7930
_|7930,7931
_|7931,7932
_|7932,7933
_|7933,7934
_|7934,7935
_|7935,7936
_|7936,7937
_|7937,7938
_|7938,7939
_|7939,7940
_|7940,7941
_|7941,7942
_|7942,7943
_|7943,7944
_|7944,7945
_|7945,7946
_|7946,7947
_|7947,7948
_|7948,7949
_|7949,7950
_|7950,7951
_|7951,7952
_|7952,7953
_|7953,7954
_|7954,7955
_|7955,7956
_|7956,7957
_|7957,7958
_|7958,7959
_|7959,7960
_|7960,7961
<EOL>|7961,7962
KLEBSIELLA|7991,8001
PNEUMONIAE|8002,8012
<EOL>|8012,8013
||8042,8043
<EOL>|8046,8047
AMPICILLIN|8047,8057
/|8057,8058
SULBACTAM|8058,8067
-|8067,8068
-|8068,8069
4|8074,8075
S|8076,8077
<EOL>|8077,8078
CEFAZOLIN|8078,8087
-|8087,8088
-|8088,8089
-|8089,8090
-|8090,8091
-|8091,8092
-|8092,8093
-|8093,8094
-|8094,8095
-|8095,8096
-|8096,8097
-|8097,8098
-|8098,8099
-|8099,8100
<|8103,8104
=|8104,8105
4|8105,8106
S|8107,8108
<EOL>|8108,8109
CEFEPIME|8109,8117
-|8117,8118
-|8118,8119
-|8119,8120
-|8120,8121
-|8121,8122
-|8122,8123
-|8123,8124
-|8124,8125
-|8125,8126
-|8126,8127
-|8127,8128
-|8128,8129
-|8129,8130
-|8130,8131
<|8134,8135
=|8135,8136
1|8136,8137
S|8138,8139
<EOL>|8139,8140
CEFTAZIDIME|8140,8151
-|8151,8152
-|8152,8153
-|8153,8154
-|8154,8155
-|8155,8156
-|8156,8157
-|8157,8158
-|8158,8159
-|8159,8160
-|8160,8161
-|8161,8162
<|8165,8166
=|8166,8167
1|8167,8168
S|8169,8170
<EOL>|8170,8171
CEFTRIAXONE|8171,8182
-|8182,8183
-|8183,8184
-|8184,8185
-|8185,8186
-|8186,8187
-|8187,8188
-|8188,8189
-|8189,8190
-|8190,8191
-|8191,8192
-|8192,8193
<|8196,8197
=|8197,8198
1|8198,8199
S|8200,8201
<EOL>|8201,8202
CIPROFLOXACIN|8202,8215
-|8215,8216
-|8216,8217
-|8217,8218
-|8218,8219
-|8219,8220
-|8220,8221
-|8221,8222
-|8222,8223
-|8223,8224
<|8224,8225
=|8225,8226
0.25|8226,8230
S|8231,8232
<EOL>|8232,8233
GENTAMICIN|8233,8243
-|8243,8244
-|8244,8245
-|8245,8246
-|8246,8247
-|8247,8248
-|8248,8249
-|8249,8250
-|8250,8251
-|8251,8252
-|8252,8253
-|8253,8254
-|8254,8255
<|8258,8259
=|8259,8260
1|8260,8261
S|8262,8263
<EOL>|8263,8264
MEROPENEM|8264,8273
-|8273,8274
-|8274,8275
-|8275,8276
-|8276,8277
-|8277,8278
-|8278,8279
-|8279,8280
-|8280,8281
-|8281,8282
-|8282,8283
-|8283,8284
-|8284,8285
-|8285,8286
<|8286,8287
=|8287,8288
0.25|8288,8292
S|8293,8294
<EOL>|8294,8295
PIPERACILLIN|8295,8307
/|8307,8308
TAZO|8308,8312
-|8312,8313
-|8313,8314
-|8314,8315
-|8315,8316
-|8316,8317
<|8320,8321
=|8321,8322
4|8322,8323
S|8324,8325
<EOL>|8325,8326
TOBRAMYCIN|8326,8336
-|8336,8337
-|8337,8338
-|8338,8339
-|8339,8340
-|8340,8341
-|8341,8342
-|8342,8343
-|8343,8344
-|8344,8345
-|8345,8346
-|8346,8347
-|8347,8348
<|8351,8352
=|8352,8353
1|8353,8354
S|8355,8356
<EOL>|8356,8357
TRIMETHOPRIM|8357,8369
/|8369,8370
SULFA|8370,8375
-|8375,8376
-|8376,8377
-|8377,8378
-|8378,8379
<|8382,8383
=|8383,8384
1|8384,8385
S|8386,8387
<EOL>|8387,8388
<EOL>|8388,8389
<EOL>|8390,8391
Mr.|8414,8417
_|8418,8419
_|8419,8420
_|8420,8421
is|8422,8424
a|8425,8426
_|8427,8428
_|8428,8429
_|8429,8430
M|8431,8432
w|8433,8434
/|8434,8435
HTN|8436,8439
,|8439,8440
HLD|8441,8444
,|8444,8445
DMII|8446,8450
,|8450,8451
and|8452,8455
old|8456,8459
MI|8460,8462
transferred|8463,8474
<EOL>|8475,8476
from|8476,8480
_|8481,8482
_|8482,8483
_|8483,8484
w|8485,8486
/|8486,8487
NSTEMI|8488,8494
w|8495,8496
/|8496,8497
diffuse|8498,8505
3|8506,8507
vessel|8508,8514
disease|8515,8522
s|8523,8524
/|8524,8525
p|8525,8526
DES|8527,8530
to|8531,8533
<EOL>|8534,8535
mid-LAD|8535,8542
occlusion|8543,8552
found|8553,8558
to|8559,8561
have|8562,8566
severe|8567,8573
Cdiff|8574,8579
.|8579,8580
<EOL>|8580,8581
<EOL>|8581,8582
ACTIVE|8582,8588
ISSUES|8589,8595
<EOL>|8595,8596
=|8596,8597
=|8597,8598
=|8598,8599
=|8599,8600
=|8600,8601
=|8601,8602
=|8602,8603
=|8603,8604
=|8604,8605
=|8605,8606
=|8606,8607
=|8607,8608
=|8608,8609
=|8609,8610
<EOL>|8610,8611
#|8611,8612
NSTEMI|8613,8619
<EOL>|8620,8621
NSTEMI|8621,8627
based|8628,8633
on|8634,8636
STE|8637,8640
aVR|8641,8644
and|8645,8648
V1|8649,8651
but|8652,8655
o|8656,8657
/|8657,8658
w|8658,8659
ST|8660,8662
depressions|8663,8674
w|8675,8676
/|8676,8677
<EOL>|8678,8679
significant|8679,8690
multi|8691,8696
vessel|8697,8703
disease|8704,8711
but|8712,8715
significant|8716,8727
stenosis|8728,8736
in|8737,8739
LAD|8740,8743
<EOL>|8744,8745
s|8745,8746
/|8746,8747
p|8747,8748
DES|8749,8752
that|8753,8757
occluded|8758,8766
diagnonal|8767,8776
.|8776,8777
Repeat|8778,8784
cath|8785,8789
unchanged|8790,8799
.|8799,8800
He|8801,8803
was|8804,8807
<EOL>|8808,8809
started|8809,8816
on|8817,8819
plavix|8820,8826
,|8826,8827
atorvastatin|8828,8840
,|8840,8841
ACE|8842,8845
-|8845,8846
I|8846,8847
,|8847,8848
and|8849,8852
metoprolol|8853,8863
.|8863,8864
Echo|8865,8869
<EOL>|8870,8871
showed|8871,8877
LVEF|8878,8882
35|8883,8885
-|8885,8886
40|8886,8888
%|8888,8889
with|8890,8894
hypokinesis|8895,8906
of|8907,8909
mid-distal|8910,8920
LV|8921,8923
segments|8924,8932
<EOL>|8933,8934
and|8934,8937
apex|8938,8942
.|8942,8943
He|8944,8946
was|8947,8950
started|8951,8958
on|8959,8961
warfarin|8962,8970
for|8971,8974
his|8975,8978
hypokinetic|8979,8990
LV|8991,8993
as|8994,8996
<EOL>|8997,8998
well|8998,9002
as|9003,9005
his|9006,9009
atrial|9010,9016
fibrillation|9017,9029
as|9030,9032
discussed|9033,9042
below|9043,9048
.|9048,9049
<EOL>|9049,9050
<EOL>|9050,9051
#|9051,9052
_|9053,9054
_|9054,9055
_|9055,9056
<EOL>|9056,9057
Possibly|9057,9065
mixed|9066,9071
cardiogenic|9072,9083
/|9083,9084
distributive|9084,9096
given|9097,9102
mixed|9103,9108
venous|9109,9115
O2|9116,9118
<EOL>|9119,9120
65|9120,9122
%|9122,9123
,|9123,9124
CI|9125,9127
2.1|9128,9131
,|9131,9132
PCWP|9133,9137
25|9138,9140
.|9140,9141
He|9142,9144
initially|9145,9154
required|9155,9163
pressors|9164,9172
and|9173,9176
balloon|9177,9184
<EOL>|9185,9186
pump|9186,9190
and|9191,9194
was|9195,9198
then|9199,9203
successfully|9204,9216
weaned|9217,9223
off|9224,9227
both|9228,9232
.|9232,9233
He|9234,9236
remained|9237,9245
<EOL>|9246,9247
hemodynamically|9247,9262
stable|9263,9269
during|9270,9276
rest|9277,9281
of|9282,9284
hospital|9285,9293
course|9294,9300
.|9300,9301
<EOL>|9302,9303
<EOL>|9303,9304
#|9304,9305
Atrial|9306,9312
Fibrillation|9313,9325
<EOL>|9325,9326
Patient|9326,9333
with|9334,9338
a|9339,9340
reported|9341,9349
history|9350,9357
of|9358,9360
paroxysmal|9361,9371
afib|9372,9376
per|9377,9380
his|9381,9384
PCP|9385,9388
<EOL>|9389,9390
for|9390,9393
which|9394,9399
he|9400,9402
was|9403,9406
maintained|9407,9417
on|9418,9420
digoxin|9421,9428
as|9429,9431
well|9432,9436
as|9437,9439
aspirin|9440,9447
325mg|9448,9453
<EOL>|9454,9455
PO|9455,9457
daily|9458,9463
prior|9464,9469
to|9470,9472
admission|9473,9482
.|9482,9483
He|9485,9487
was|9488,9491
found|9492,9497
to|9498,9500
be|9501,9503
in|9504,9506
atrial|9507,9513
<EOL>|9514,9515
fibrillation|9515,9527
during|9528,9534
admission|9535,9544
and|9545,9548
the|9549,9552
decision|9553,9561
was|9562,9565
made|9566,9570
to|9571,9573
<EOL>|9574,9575
anticoagulate|9575,9588
with|9589,9593
Coumadin|9594,9602
.|9602,9603
He|9605,9607
was|9608,9611
continued|9612,9621
on|9622,9624
home|9625,9629
dose|9630,9634
<EOL>|9635,9636
digoxin|9636,9643
.|9643,9644
His|9646,9649
home|9650,9654
dose|9655,9659
aspirin|9660,9667
was|9668,9671
decreased|9672,9681
as|9682,9684
discussed|9685,9694
above|9695,9700
<EOL>|9701,9702
with|9702,9706
initiation|9707,9717
of|9718,9720
Coumadin|9721,9729
.|9729,9730
<EOL>|9730,9731
<EOL>|9731,9732
#|9732,9733
Hematuria|9734,9743
:|9743,9744
<EOL>|9745,9746
Likely|9746,9752
traumatic|9753,9762
in|9763,9765
setting|9766,9773
of|9774,9776
systemic|9777,9785
anticoagulation|9786,9801
,|9801,9802
as|9803,9805
<EOL>|9806,9807
patient|9807,9814
pulled|9815,9821
at|9822,9824
_|9825,9826
_|9826,9827
_|9827,9828
.|9828,9829
Cytology|9830,9838
was|9839,9842
negative|9843,9851
.|9851,9852
He|9853,9855
will|9856,9860
followup|9861,9869
<EOL>|9870,9871
outpatient|9871,9881
with|9882,9886
urology|9887,9894
.|9894,9895
<EOL>|9895,9896
<EOL>|9896,9897
#|9897,9898
Dyspnea|9899,9906
:|9906,9907
<EOL>|9908,9909
Patient|9909,9916
had|9917,9920
acute|9921,9926
episodes|9927,9935
of|9936,9938
dyspnea|9939,9946
.|9946,9947
This|9949,9953
was|9954,9957
mainly|9958,9964
<EOL>|9965,9966
attributed|9966,9976
to|9977,9979
pulmonary|9980,9989
edema|9990,9995
and|9996,9999
improved|10000,10008
with|10009,10013
diruesis|10014,10022
.|10022,10023
<EOL>|10025,10026
Additionally|10026,10038
,|10038,10039
CXR|10040,10043
showed|10044,10050
possible|10051,10059
consolidation|10060,10073
of|10074,10076
RUL|10077,10080
,|10080,10081
<EOL>|10082,10083
concerning|10083,10093
for|10094,10097
aspiration|10098,10108
pneumonia|10109,10118
.|10118,10119
However|10120,10127
,|10127,10128
treatment|10129,10138
was|10139,10142
<EOL>|10143,10144
deferred|10144,10152
as|10153,10155
he|10156,10158
had|10159,10162
no|10163,10165
other|10166,10171
focal|10172,10177
signs|10178,10183
of|10184,10186
infectious|10187,10197
pna|10198,10201
.|10201,10202
He|10204,10206
<EOL>|10207,10208
did|10208,10211
have|10212,10216
sputum|10217,10223
cultures|10224,10232
which|10233,10238
grew|10239,10243
Klebsiella|10244,10254
pneumonia|10255,10264
but|10265,10268
on|10269,10271
<EOL>|10272,10273
discussion|10273,10283
with|10284,10288
ID|10289,10291
,|10291,10292
felt|10293,10297
this|10298,10302
did|10303,10306
not|10307,10310
warrant|10311,10318
any|10319,10322
treatment|10323,10332
as|10333,10335
<EOL>|10336,10337
he|10337,10339
was|10340,10343
asymptomatic|10344,10356
.|10356,10357
He|10359,10361
was|10362,10365
discharged|10366,10376
on|10377,10379
po|10380,10382
lasix|10383,10388
20|10389,10391
mg|10392,10394
daily|10395,10400
<EOL>|10401,10402
with|10402,10406
next|10407,10411
electrolytes|10412,10424
to|10425,10427
be|10428,10430
checked|10431,10438
_|10439,10440
_|10440,10441
_|10441,10442
.|10442,10443
<EOL>|10444,10445
<EOL>|10446,10447
#|10447,10448
C|10449,10450
diff|10451,10455
,|10455,10456
severe|10457,10463
:|10463,10464
<EOL>|10465,10466
Had|10466,10469
loose|10470,10475
stool|10476,10481
in|10482,10484
setting|10485,10492
of|10493,10495
antibiotic|10496,10506
tx|10507,10509
for|10510,10513
Hpylori|10514,10521
<EOL>|10522,10523
(|10523,10524
initiated|10524,10533
outpatient|10534,10544
)|10544,10545
.|10545,10546
Given|10547,10552
WBC|10553,10556
>|10557,10558
15|10558,10560
,|10560,10561
_|10562,10563
_|10563,10564
_|10564,10565
,|10565,10566
age|10567,10570
>|10571,10572
_|10572,10573
_|10573,10574
_|10574,10575
treated|10576,10583
as|10584,10586
<EOL>|10587,10588
severe|10588,10594
.|10594,10595
Patient|10596,10603
was|10604,10607
started|10608,10615
on|10616,10618
vancomycin|10619,10629
125mg|10630,10635
PO|10636,10638
qid|10639,10642
for|10643,10646
14|10647,10649
<EOL>|10650,10651
day|10651,10654
course|10655,10661
(|10662,10663
day|10663,10666
_|10667,10668
_|10668,10669
_|10669,10670
,|10670,10671
last|10672,10676
day|10677,10680
_|10681,10682
_|10682,10683
_|10683,10684
.|10684,10685
<EOL>|10686,10687
<EOL>|10688,10689
#|10689,10690
GASTROESOPHAGEAL|10691,10707
REFLUX|10708,10714
DISEASE|10715,10722
(|10723,10724
GERD|10724,10728
)|10728,10729
:|10729,10730
<EOL>|10731,10732
Endoscopy|10732,10741
confirmed|10742,10751
H|10752,10753
Pylori|10754,10760
treated|10761,10768
with|10769,10773
PPI|10774,10777
+|10778,10779
<EOL>|10780,10781
clarithromycin|10781,10795
/|10795,10796
amoxicillin|10796,10807
since|10808,10813
_|10814,10815
_|10815,10816
_|10816,10817
for|10818,10821
14|10822,10824
days|10825,10829
.|10829,10830
Omeprazole|10831,10841
<EOL>|10842,10843
was|10843,10846
continued|10847,10856
.|10856,10857
Antibiotics|10858,10869
held|10870,10874
in|10875,10877
setting|10878,10885
of|10886,10888
c|10889,10890
.|10890,10891
diff|10891,10895
infection|10896,10905
.|10905,10906
<EOL>|10907,10908
<EOL>|10908,10909
#|10909,10910
Delirium|10911,10919
:|10919,10920
<EOL>|10921,10922
Patient|10922,10929
with|10930,10934
frequent|10935,10943
sundowning|10944,10954
during|10955,10961
hospitalization|10962,10977
<EOL>|10978,10979
requiring|10979,10988
Seroquel|10989,10997
po|10998,11000
.|11000,11001
<EOL>|11001,11002
<EOL>|11002,11003
CHRONIC|11003,11010
ISSUES|11011,11017
<EOL>|11017,11018
=|11018,11019
=|11019,11020
=|11020,11021
=|11021,11022
=|11022,11023
=|11023,11024
=|11024,11025
=|11025,11026
=|11026,11027
=|11027,11028
=|11028,11029
=|11029,11030
=|11030,11031
=|11031,11032
=|11032,11033
<EOL>|11033,11034
#|11034,11035
Spinal|11036,11042
Stenosis|11043,11051
:|11051,11052
Continued|11053,11062
gabapentin|11063,11073
,|11073,11074
d|11075,11076
/|11076,11077
ced|11077,11080
naproxen|11081,11089
.|11089,11090
Did|11092,11095
<EOL>|11096,11097
not|11097,11100
complain|11101,11109
of|11110,11112
pain|11113,11117
throughout|11118,11128
hospital|11129,11137
course|11138,11144
.|11144,11145
Explained|11147,11156
he|11157,11159
<EOL>|11160,11161
should|11161,11167
not|11168,11171
take|11172,11176
any|11177,11180
more|11181,11185
NSAIDS|11186,11192
in|11193,11195
setting|11196,11203
of|11204,11206
recent|11207,11213
ACS|11214,11217
and|11218,11221
now|11222,11225
<EOL>|11226,11227
on|11227,11229
Coumadin|11230,11238
,|11238,11239
Plavix|11240,11246
and|11247,11250
asa|11251,11254
.|11254,11255
<EOL>|11256,11257
#|11257,11258
DM|11259,11261
:|11261,11262
maintained|11263,11273
on|11274,11276
ISS|11277,11280
during|11281,11287
admission|11288,11297
and|11298,11301
discharged|11302,11312
on|11313,11315
home|11316,11320
<EOL>|11321,11322
glipizide|11322,11331
and|11332,11335
metformin|11336,11345
<EOL>|11345,11346
#|11346,11347
HTN|11348,11351
:|11351,11352
Home|11353,11357
dose|11358,11362
metoprolol|11363,11373
uptitrated|11374,11384
.|11384,11385
Home|11387,11391
dose|11392,11396
lisinopril|11397,11407
<EOL>|11408,11409
decreased|11409,11418
.|11418,11419
Home|11421,11425
dose|11426,11430
imdur|11431,11436
discontinued|11437,11449
.|11449,11450
<EOL>|11450,11451
#|11451,11452
HLD|11453,11456
:|11456,11457
Transitioned|11458,11470
home|11471,11475
dose|11476,11480
simvastatin|11481,11492
to|11493,11495
atorvastatin|11496,11508
<EOL>|11508,11509
<EOL>|11509,11510
TRANSITIONAL|11510,11522
ISSUES|11523,11529
<EOL>|11529,11530
=|11530,11531
=|11531,11532
=|11532,11533
=|11533,11534
=|11534,11535
=|11535,11536
=|11536,11537
=|11537,11538
=|11538,11539
=|11539,11540
=|11540,11541
=|11541,11542
=|11542,11543
=|11543,11544
=|11544,11545
=|11545,11546
=|11546,11547
=|11547,11548
=|11548,11549
=|11549,11550
=|11550,11551
<EOL>|11551,11552
-|11552,11553
Discharge|11554,11563
weight|11564,11570
:|11570,11571
63.7|11572,11576
kg|11576,11578
<EOL>|11579,11580
-|11580,11581
patient|11582,11589
will|11590,11594
require|11595,11602
urology|11603,11610
followup|11611,11619
given|11620,11625
hematuria|11626,11635
during|11636,11642
<EOL>|11643,11644
admission|11644,11653
.|11653,11654
Urine|11656,11661
cytology|11662,11670
negative|11671,11679
.|11679,11680
<EOL>|11680,11681
-|11681,11682
patient|11683,11690
will|11691,11695
need|11696,11700
to|11701,11703
be|11704,11706
treated|11707,11714
for|11715,11718
hpylori|11719,11726
once|11727,11731
he|11732,11734
completes|11735,11744
<EOL>|11745,11746
a|11746,11747
course|11748,11754
of|11755,11757
PO|11758,11760
Vancomycin|11761,11771
for|11772,11775
Severe|11776,11782
CDiff|11783,11788
<EOL>|11788,11789
-|11789,11790
Please|11791,11797
check|11798,11803
electrolytes|11804,11816
on|11817,11819
_|11820,11821
_|11821,11822
_|11822,11823
on|11824,11826
lasix|11827,11832
<EOL>|11832,11833
-|11833,11834
Coumadin|11835,11843
initiated|11844,11853
given|11854,11859
atrial|11860,11866
fibrillation|11867,11879
,|11879,11880
ASA|11881,11884
decreased|11885,11894
<EOL>|11895,11896
from|11896,11900
325|11901,11904
mg|11905,11907
to|11908,11910
81|11911,11913
mg|11914,11916
daily|11917,11922
<EOL>|11922,11923
-|11923,11924
Started|11925,11932
on|11933,11935
Plavix|11936,11942
given|11943,11948
recent|11949,11955
stent|11956,11961
placement|11962,11971
,|11971,11972
atorvastatin|11973,11985
<EOL>|11986,11987
80|11987,11989
mg|11990,11992
(|11993,11994
stopped|11994,12001
simvastatin|12002,12013
)|12013,12014
,|12014,12015
and|12016,12019
Lasix|12020,12025
20|12026,12028
mg|12029,12031
po|12032,12034
daily|12035,12040
<EOL>|12040,12041
-|12041,12042
Home|12043,12047
metoprolol|12048,12058
was|12059,12062
increased|12063,12072
from|12073,12077
25|12078,12080
mg|12081,12083
XL|12084,12086
to|12087,12089
50|12090,12092
mg|12093,12095
XL|12096,12098
daily|12099,12104
,|12104,12105
<EOL>|12106,12107
lisinopril|12107,12117
decreased|12118,12127
to|12128,12130
2.5|12131,12134
mg|12135,12137
po|12138,12140
daily|12141,12146
and|12147,12150
home|12151,12155
imdur|12156,12161
was|12162,12165
<EOL>|12166,12167
discontinued|12167,12179
<EOL>|12179,12180
-|12180,12181
patient|12182,12189
will|12190,12194
need|12195,12199
to|12200,12202
continue|12203,12211
a|12212,12213
14|12214,12216
day|12217,12220
course|12221,12227
of|12228,12230
PO|12231,12233
Vanc|12234,12238
(|12239,12240
day|12240,12243
<EOL>|12244,12245
_|12245,12246
_|12246,12247
_|12247,12248
-|12248,12249
_|12250,12251
_|12251,12252
_|12252,12253
last|12254,12258
day|12259,12262
_|12263,12264
_|12264,12265
_|12265,12266
for|12267,12270
cdiff|12271,12276
infection|12277,12286
<EOL>|12286,12287
-|12287,12288
Patient|12289,12296
instructed|12297,12307
to|12308,12310
not|12311,12314
take|12315,12319
any|12320,12323
NSAIDS|12324,12330
<EOL>|12330,12331
-|12331,12332
SLP|12333,12336
treatment|12337,12346
at|12347,12349
rehab|12350,12355
for|12356,12359
pharyngeal|12360,12370
strengthening|12371,12384
exercises|12385,12394
<EOL>|12394,12395
<EOL>|12396,12397
Medications|12397,12408
on|12409,12411
Admission|12412,12421
:|12421,12422
<EOL>|12422,12423
The|12423,12426
Preadmission|12427,12439
Medication|12440,12450
list|12451,12455
is|12456,12458
accurate|12459,12467
and|12468,12471
complete|12472,12480
.|12480,12481
<EOL>|12481,12482
1.|12482,12484
Gabapentin|12485,12495
600|12496,12499
mg|12500,12502
PO|12503,12505
TID|12506,12509
<EOL>|12510,12511
2.|12511,12513
Naproxen|12514,12522
500|12523,12526
mg|12527,12529
PO|12530,12532
DAILY|12533,12538
<EOL>|12539,12540
3.|12540,12542
MetFORMIN|12543,12552
(|12553,12554
Glucophage|12554,12564
)|12564,12565
500|12566,12569
mg|12570,12572
PO|12573,12575
BID|12576,12579
<EOL>|12580,12581
4.|12581,12583
Metoprolol|12584,12594
Succinate|12595,12604
XL|12605,12607
25|12608,12610
mg|12611,12613
PO|12614,12616
DAILY|12617,12622
<EOL>|12623,12624
5.|12624,12626
GlipiZIDE|12627,12636
2.5|12637,12640
mg|12641,12643
PO|12644,12646
BID|12647,12650
<EOL>|12651,12652
6.|12652,12654
Simvastatin|12655,12666
40|12667,12669
mg|12670,12672
PO|12673,12675
QPM|12676,12679
<EOL>|12680,12681
7.|12681,12683
Isosorbide|12684,12694
Mononitrate|12695,12706
(|12707,12708
Extended|12708,12716
Release|12717,12724
)|12724,12725
60|12726,12728
mg|12729,12731
PO|12732,12734
DAILY|12735,12740
<EOL>|12741,12742
8.|12742,12744
Lisinopril|12745,12755
10|12756,12758
mg|12759,12761
PO|12762,12764
DAILY|12765,12770
<EOL>|12771,12772
9.|12772,12774
Digoxin|12775,12782
0.125|12783,12788
mg|12789,12791
PO|12792,12794
DAILY|12795,12800
<EOL>|12801,12802
10.|12802,12805
Aspirin|12806,12813
325|12814,12817
mg|12818,12820
PO|12821,12823
DAILY|12824,12829
<EOL>|12830,12831
<EOL>|12831,12832
<EOL>|12833,12834
Discharge|12834,12843
Medications|12844,12855
:|12855,12856
<EOL>|12856,12857
1.|12857,12859
Aspirin|12860,12867
EC|12868,12870
81|12871,12873
mg|12874,12876
PO|12877,12879
DAILY|12880,12885
<EOL>|12886,12887
2.|12887,12889
Digoxin|12890,12897
0.125|12898,12903
mg|12904,12906
PO|12907,12909
DAILY|12910,12915
<EOL>|12916,12917
3.|12917,12919
Metoprolol|12920,12930
Succinate|12931,12940
XL|12941,12943
50|12944,12946
mg|12947,12949
PO|12950,12952
DAILY|12953,12958
<EOL>|12959,12960
4.|12960,12962
Atorvastatin|12963,12975
80|12976,12978
mg|12979,12981
PO|12982,12984
QPM|12985,12988
<EOL>|12989,12990
5.|12990,12992
Warfarin|12993,13001
4|13002,13003
mg|13004,13006
PO|13007,13009
DAILY16|13010,13017
<EOL>|13018,13019
6.|13019,13021
GlipiZIDE|13022,13031
2.5|13032,13035
mg|13036,13038
PO|13039,13041
BID|13042,13045
<EOL>|13046,13047
7.|13047,13049
Clopidogrel|13050,13061
75|13062,13064
mg|13065,13067
PO|13068,13070
DAILY|13071,13076
<EOL>|13077,13078
8.|13078,13080
Omeprazole|13081,13091
20|13092,13094
mg|13095,13097
PO|13098,13100
BID|13101,13104
<EOL>|13105,13106
9.|13106,13108
Vancomycin|13109,13119
Oral|13120,13124
Liquid|13125,13131
_|13132,13133
_|13133,13134
_|13134,13135
mg|13136,13138
PO|13139,13141
Q6H|13142,13145
<EOL>|13146,13147
10.|13147,13150
MetFORMIN|13151,13160
(|13161,13162
Glucophage|13162,13172
)|13172,13173
500|13174,13177
mg|13178,13180
PO|13181,13183
BID|13184,13187
<EOL>|13188,13189
11.|13189,13192
Gabapentin|13193,13203
600|13204,13207
mg|13208,13210
PO|13211,13213
TID|13214,13217
<EOL>|13218,13219
12.|13219,13222
Lisinopril|13223,13233
2.5|13234,13237
mg|13238,13240
PO|13241,13243
DAILY|13244,13249
<EOL>|13250,13251
13.|13251,13254
Furosemide|13255,13265
20|13266,13268
mg|13269,13271
PO|13272,13274
DAILY|13275,13280
<EOL>|13281,13282
<EOL>|13282,13283
<EOL>|13284,13285
Discharge|13285,13294
Disposition|13295,13306
:|13306,13307
<EOL>|13307,13308
Extended|13308,13316
Care|13317,13321
<EOL>|13321,13322
<EOL>|13323,13324
Facility|13324,13332
:|13332,13333
<EOL>|13333,13334
_|13334,13335
_|13335,13336
_|13336,13337
<EOL>|13337,13338
<EOL>|13339,13340
Discharge|13340,13349
Diagnosis|13350,13359
:|13359,13360
<EOL>|13360,13361
NSTEMI|13361,13367
s|13368,13369
/|13369,13370
p|13370,13371
_|13372,13373
_|13373,13374
_|13374,13375
,|13375,13376
likely|13377,13383
mixed|13384,13389
cardiogenic|13390,13401
/|13401,13402
distributive|13402,13414
<EOL>|13415,13416
Hematuria|13416,13425
<EOL>|13425,13426
Dyspnea|13426,13433
<EOL>|13433,13434
C.|13434,13436
dif|13437,13440
,|13440,13441
severe|13442,13448
<EOL>|13448,13449
GERD|13449,13453
<EOL>|13453,13454
Delirium|13454,13462
<EOL>|13462,13463
<EOL>|13463,13464
<EOL>|13465,13466
Mental|13487,13493
Status|13494,13500
:|13500,13501
Clear|13502,13507
and|13508,13511
coherent|13512,13520
.|13520,13521
<EOL>|13521,13522
Level|13522,13527
of|13528,13530
Consciousness|13531,13544
:|13544,13545
Alert|13546,13551
and|13552,13555
interactive|13556,13567
.|13567,13568
<EOL>|13568,13569
<EOL>|13570,13571
Dear|13595,13599
Mr.|13600,13603
_|13604,13605
_|13605,13606
_|13606,13607
,|13607,13608
<EOL>|13608,13609
<EOL>|13609,13610
You|13610,13613
were|13614,13618
admitted|13619,13627
to|13628,13630
_|13631,13632
_|13632,13633
_|13633,13634
because|13635,13642
you|13643,13646
were|13647,13651
experiencing|13652,13664
chest|13665,13670
<EOL>|13671,13672
pain|13672,13676
due|13677,13680
to|13681,13683
a|13684,13685
heart|13686,13691
attack|13692,13698
.|13698,13699
In|13700,13702
the|13703,13706
cath|13707,13711
lab|13712,13715
you|13716,13719
were|13720,13724
found|13725,13730
to|13731,13733
<EOL>|13734,13735
have|13735,13739
blockage|13740,13748
of|13749,13751
your|13752,13756
arteries|13757,13765
,|13765,13766
and|13767,13770
a|13771,13772
stent|13773,13778
was|13779,13782
placed|13783,13789
.|13789,13790
We|13791,13793
also|13794,13798
<EOL>|13799,13800
managed|13800,13807
your|13808,13812
low|13813,13816
blood|13817,13822
pressure|13823,13831
,|13831,13832
infectious|13833,13843
diarrhea|13844,13852
,|13852,13853
and|13854,13857
trauma|13858,13864
<EOL>|13865,13866
from|13866,13870
foley|13871,13876
placement|13877,13886
.|13886,13887
You|13888,13891
responded|13892,13901
well|13902,13906
.|13906,13907
<EOL>|13908,13909
<EOL>|13909,13910
Please|13910,13916
continue|13917,13925
taking|13926,13932
your|13933,13937
medications|13938,13949
as|13950,13952
prescribed|13953,13963
.|13963,13964
You|13966,13969
are|13970,13973
<EOL>|13974,13975
being|13975,13980
started|13981,13988
on|13989,13991
coumadin|13992,14000
.|14000,14001
Please|14003,14009
do|14010,14012
not|14013,14016
take|14017,14021
any|14022,14025
non-steroidal|14026,14039
<EOL>|14040,14041
antiinflammatory|14041,14057
drugs|14058,14063
(|14064,14065
NSAIDS|14065,14071
)|14071,14072
such|14073,14077
as|14078,14080
ibuprofen|14081,14090
,|14090,14091
advil|14092,14097
,|14097,14098
<EOL>|14099,14100
motrin|14100,14106
,|14106,14107
aleve|14108,14113
,|14113,14114
naproxen|14115,14123
.|14123,14124
Please|14126,14132
also|14133,14137
follow|14138,14144
-|14144,14145
up|14145,14147
with|14148,14152
your|14153,14157
<EOL>|14158,14159
cardiology|14159,14169
and|14170,14173
PCP|14174,14177
appointments|14178,14190
as|14191,14193
scheduled|14194,14203
<EOL>|14203,14204
<EOL>|14204,14205
It|14205,14207
was|14208,14211
a|14212,14213
pleasure|14214,14222
taking|14223,14229
care|14230,14234
of|14235,14237
you|14238,14241
,|14241,14242
<EOL>|14242,14243
Your|14243,14247
_|14248,14249
_|14249,14250
_|14250,14251
Care|14252,14256
Team|14257,14261
<EOL>|14261,14262
<EOL>|14263,14264
Followup|14264,14272
Instructions|14273,14285
:|14285,14286
<EOL>|14286,14287
_|14287,14288
_|14288,14289
_|14289,14290
<EOL>|14290,14291

