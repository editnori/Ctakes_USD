 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|26,30
No|31,33
:|33,34
_|37,38
_|38,39
_|39,40
<EOL>|40,41
<EOL>|42,43
Admission|43,52
Date|53,57
:|57,58
_|60,61
_|61,62
_|62,63
Discharge|77,86
Date|87,91
:|91,92
_|95,96
_|96,97
_|97,98
<EOL>|98,99
<EOL>|100,101
Date|101,105
of|106,108
Birth|109,114
:|114,115
_|117,118
_|118,119
_|119,120
Sex|133,136
:|136,137
F|140,141
<EOL>|141,142
<EOL>|143,144
Service|144,151
:|151,152
NEUROSURGERY|153,165
<EOL>|165,166
<EOL>|167,168
Penicillins|180,191
<EOL>|191,192
<EOL>|193,194
Attending|194,203
:|203,204
_|205,206
_|206,207
_|207,208
<EOL>|208,209
<EOL>|210,211
Wound|228,233
Infection|234,243
<EOL>|243,244
<EOL>|245,246
Major|246,251
Surgical|252,260
or|261,263
Invasive|264,272
Procedure|273,282
:|282,283
<EOL>|283,284
Right|284,289
Craniotomy|290,300
and|301,304
Evacuation|305,315
of|316,318
Abscess|319,326
on|327,329
_|330,331
_|331,332
_|332,333
<EOL>|333,334
<EOL>|335,336
Ms.|364,367
_|368,369
_|369,370
_|370,371
is|372,374
a|375,376
_|377,378
_|378,379
_|379,380
y|381,382
/|382,383
o|383,384
woman|385,390
with|391,395
a|396,397
past|398,402
medical|403,410
history|411,418
<EOL>|418,419
of|419,421
MS|422,424
,|424,425
and|426,429
a|430,431
right|432,437
parietal|438,446
brain|447,452
abscess|453,460
which|461,466
was|467,470
discovered|471,481
<EOL>|481,482
approxiamtely|482,495
one|496,499
month|500,505
ago|506,509
,|509,510
when|511,515
she|516,519
presented|520,529
with|530,534
left|535,539
arm|540,543
<EOL>|544,545
and|545,548
<EOL>|548,549
face|549,553
numbness|554,562
.|562,563
The|564,567
abscess|568,575
was|576,579
drained|580,587
in|588,590
the|591,594
OR|595,597
on|598,600
_|601,602
_|602,603
_|603,604
,|604,605
and|606,609
she|610,613
<EOL>|613,614
was|614,617
initially|618,627
started|628,635
on|636,638
broad|639,644
spectrum|645,653
antibiotics|654,665
until|666,671
<EOL>|672,673
culture|673,680
<EOL>|680,681
data|681,685
returned|686,694
with|695,699
S.|700,702
anginosus|703,712
and|713,716
fusobacterium|717,730
,|730,731
she|732,735
was|736,739
then|740,744
<EOL>|744,745
transitioned|745,757
to|758,760
Ceftriaxone|761,772
2g|773,775
IV|776,778
q12h|779,783
,|783,784
and|785,788
flagyl|789,795
500mg|796,801
TID|802,805
,|805,806
<EOL>|806,807
which|807,812
she|813,816
has|817,820
been|821,825
on|826,828
since|829,834
through|835,842
her|843,846
PICC|847,851
line|852,856
.|856,857
On|858,860
_|861,862
_|862,863
_|863,864
,|864,865
she|866,869
<EOL>|869,870
was|870,873
seen|874,878
in|879,881
_|882,883
_|883,884
_|884,885
clinic|886,892
and|893,896
a|897,898
repeat|899,905
MRI|906,909
was|910,913
performed|914,923
<EOL>|923,924
which|924,929
revealed|930,938
increased|939,948
edema|949,954
with|955,959
persistent|960,970
ring|971,975
enhancing|976,985
<EOL>|985,986
abnormality|986,997
at|998,1000
the|1001,1004
right|1005,1010
parietal|1011,1019
surgical|1020,1028
site|1029,1033
,|1033,1034
concerning|1035,1045
for|1046,1049
<EOL>|1049,1050
ongoing|1050,1057
abscess|1058,1065
.|1065,1066
She|1067,1070
was|1071,1074
therefore|1075,1084
scheduled|1085,1094
for|1095,1098
repeat|1099,1105
drainage|1106,1114
<EOL>|1114,1115
on|1115,1117
_|1118,1119
_|1119,1120
_|1120,1121
.|1121,1122
She|1123,1126
was|1127,1130
seen|1131,1135
as|1136,1138
an|1139,1141
outpatient|1142,1152
in|1153,1155
the|1156,1159
infectious|1160,1170
disease|1171,1178
<EOL>|1178,1179
office|1179,1185
today|1186,1191
,|1191,1192
_|1193,1194
_|1194,1195
_|1195,1196
,|1196,1197
and|1198,1201
it|1202,1204
was|1205,1208
recommended|1209,1220
that|1221,1225
she|1226,1229
be|1230,1232
admitted|1233,1241
<EOL>|1241,1242
to|1242,1244
the|1245,1248
hospital|1249,1257
one|1258,1261
day|1262,1265
early|1266,1271
for|1272,1275
broadening|1276,1286
of|1287,1289
her|1290,1293
antibiotic|1294,1304
<EOL>|1304,1305
regimen|1305,1312
prior|1313,1318
to|1319,1321
drainage|1322,1330
.|1330,1331
<EOL>|1331,1332
<EOL>|1332,1333
She|1333,1336
states|1337,1343
that|1344,1348
over|1349,1353
the|1354,1357
past|1358,1362
month|1363,1368
,|1368,1369
her|1370,1373
symptoms|1374,1382
,|1382,1383
including|1384,1393
<EOL>|1394,1395
left|1395,1399
<EOL>|1399,1400
upper|1400,1405
extremity|1406,1415
weakness|1416,1424
and|1425,1428
numbness|1429,1437
,|1437,1438
have|1439,1443
come|1444,1448
and|1449,1452
gone|1453,1457
,|1457,1458
<EOL>|1458,1459
although|1459,1467
she|1468,1471
thinks|1472,1478
that|1479,1483
overall|1484,1491
they|1492,1496
have|1497,1501
worsened|1502,1510
slightly|1511,1519
.|1519,1520
<EOL>|1521,1522
She|1522,1525
<EOL>|1525,1526
denies|1526,1532
any|1533,1536
fevers|1537,1543
/|1543,1544
chills|1544,1550
,|1550,1551
or|1552,1554
headaches|1555,1564
.|1564,1565
No|1566,1568
changes|1569,1576
in|1577,1579
vision|1580,1586
,|1586,1587
<EOL>|1588,1589
leg|1589,1592
<EOL>|1592,1593
weakness|1593,1601
or|1602,1604
trouble|1605,1612
with|1613,1617
coordination|1618,1630
or|1631,1633
balance|1634,1641
.|1641,1642
<EOL>|1642,1643
<EOL>|1643,1644
She|1644,1647
denies|1648,1654
shortness|1655,1664
of|1665,1667
breath|1668,1674
,|1674,1675
chest|1676,1681
pain|1682,1686
,|1686,1687
abdominal|1688,1697
pain|1698,1702
.|1702,1703
<EOL>|1703,1704
<EOL>|1704,1705
<EOL>|1706,1707
Multiple|1729,1737
sclerosis|1738,1747
<EOL>|1747,1748
<EOL>|1749,1750
:|1764,1765
<EOL>|1765,1766
_|1766,1767
_|1767,1768
_|1768,1769
<EOL>|1769,1770
:|1784,1785
<EOL>|1785,1786
Mother|1786,1792
with|1793,1797
pancreatic|1798,1808
cancer|1809,1815
,|1815,1816
brother|1817,1824
-|1824,1825
lung|1825,1829
cancer|1830,1836
,|1836,1837
two|1838,1841
sisters|1842,1849
<EOL>|1850,1851
with|1851,1855
brain|1856,1861
cancer|1862,1868
.|1868,1869
<EOL>|1869,1870
<EOL>|1870,1871
<EOL>|1872,1873
PHYSICAL|1888,1896
EXAMINATION|1897,1908
ON|1909,1911
ADMISSION|1912,1921
:|1921,1922
<EOL>|1922,1923
General|1946,1953
-|1954,1955
Appears|1956,1963
comfortable|1964,1975
<EOL>|1975,1976
HEENT|1976,1981
-|1982,1983
MMM|1984,1987
,|1987,1988
no|1989,1991
scleral|1992,1999
icterus|2000,2007
,|2007,2008
no|2009,2011
proptosis|2012,2021
,|2021,2022
sclera|2023,2029
and|2030,2033
<EOL>|2033,2034
conjunctiva|2034,2045
with|2046,2050
no|2051,2053
edema|2054,2059
/|2059,2060
injection|2060,2069
.|2069,2070
Neck|2071,2075
is|2076,2078
supple|2079,2085
.|2085,2086
<EOL>|2086,2087
CV|2087,2089
-|2090,2091
RRR|2092,2095
,|2095,2096
no|2097,2099
murmurs|2100,2107
,|2107,2108
rubs|2109,2113
,|2113,2114
or|2115,2117
gallops|2118,2125
.|2125,2126
No|2127,2129
carotid|2130,2137
bruits|2138,2144
<EOL>|2144,2145
Pulm|2145,2149
-|2150,2151
CTA|2152,2155
b|2156,2157
/|2157,2158
l|2158,2159
<EOL>|2159,2160
Abd|2160,2163
-|2164,2165
soft|2166,2170
,|2170,2171
non-tender|2172,2182
,|2182,2183
normal|2184,2190
bowel|2191,2196
sounds|2197,2203
<EOL>|2203,2204
Extremities|2204,2215
-|2216,2217
no|2218,2220
cyanosis|2221,2229
,|2229,2230
no|2231,2233
edema|2234,2239
<EOL>|2239,2240
Skin|2240,2244
-|2245,2246
warm|2247,2251
and|2252,2255
pink|2256,2260
with|2261,2265
no|2266,2268
rashes|2269,2275
<EOL>|2275,2276
Neurologic|2276,2286
Exam|2287,2291
:|2291,2292
<EOL>|2292,2293
MENTAL|2293,2299
STATUS|2300,2306
:|2306,2307
Awake|2308,2313
and|2314,2317
alert|2318,2323
,|2323,2324
oriented|2325,2333
x|2334,2335
3|2336,2337
,|2337,2338
responds|2339,2347
to|2348,2350
<EOL>|2350,2351
multi-step|2351,2361
commands|2362,2370
which|2371,2376
cross|2377,2382
the|2383,2386
midline|2387,2394
.|2394,2395
Knows|2396,2401
recent|2402,2408
and|2409,2412
<EOL>|2412,2413
distant|2413,2420
events|2421,2427
.|2427,2428
No|2429,2431
hemisensory|2432,2443
or|2444,2446
visual|2447,2453
neglect|2454,2461
.|2461,2462
<EOL>|2462,2463
<EOL>|2463,2464
PHYSICAL|2464,2472
EXAMINATION|2473,2484
ON|2485,2487
DISCHARGE|2488,2497
:|2497,2498
<EOL>|2498,2499
XXXXXX|2499,2505
<EOL>|2505,2506
<EOL>|2507,2508
Pertinent|2508,2517
Results|2518,2525
:|2525,2526
<EOL>|2526,2527
MRI|2527,2530
Brain|2531,2536
for|2537,2540
Operative|2541,2550
Planning|2551,2559
:|2559,2560
_|2561,2562
_|2562,2563
_|2563,2564
<EOL>|2564,2565
Decrease|2565,2573
in|2574,2576
size|2577,2581
of|2582,2584
known|2585,2590
right|2591,2596
frontal|2597,2604
vertex|2605,2611
rim|2612,2615
-|2615,2616
enhancing|2616,2625
<EOL>|2626,2627
lesion|2627,2633
,|2633,2634
but|2635,2638
unchanged|2639,2648
vasogenic|2649,2658
edema|2659,2664
and|2665,2668
mass|2669,2673
effect|2674,2680
.|2680,2681
<EOL>|2681,2682
<EOL>|2682,2683
Non-Contrast|2683,2695
Head|2696,2700
CT|2701,2703
:|2703,2704
_|2705,2706
_|2706,2707
_|2707,2708
<EOL>|2708,2709
POST-OP|2709,2716
SCAN|2717,2721
<EOL>|2722,2723
Status|2737,2743
post|2744,2748
redo|2749,2753
right|2754,2759
parietal|2760,2768
vertex|2769,2775
craniotomy|2776,2786
with|2787,2791
no|2792,2794
<EOL>|2795,2796
evidence|2796,2804
of|2805,2807
hemorrhage|2808,2818
.|2818,2819
Stable|2821,2827
vasogenic|2828,2837
edema|2838,2843
extending|2844,2853
in|2854,2856
the|2857,2860
<EOL>|2861,2862
right|2862,2867
frontal|2868,2875
and|2876,2879
parietal|2880,2888
lobes|2889,2894
.|2894,2895
<EOL>|2896,2897
<EOL>|2897,2898
<EOL>|2899,2900
Ms.|2923,2926
_|2927,2928
_|2928,2929
_|2929,2930
is|2931,2933
a|2934,2935
_|2936,2937
_|2937,2938
_|2938,2939
y|2940,2941
/|2941,2942
o|2942,2943
F|2944,2945
who|2946,2949
was|2950,2953
admitted|2954,2962
to|2963,2965
the|2966,2969
neurosurgery|2970,2982
<EOL>|2983,2984
service|2984,2991
on|2992,2994
the|2995,2998
day|2999,3002
of|3003,3005
admission|3006,3015
,|3015,3016
_|3017,3018
_|3018,3019
_|3019,3020
from|3021,3025
the|3026,3029
Infectious|3030,3040
<EOL>|3041,3042
Disease|3042,3049
Clinic|3050,3056
in|3057,3059
anticipation|3060,3072
for|3073,3076
evacuation|3077,3087
of|3088,3090
the|3091,3094
brain|3095,3100
<EOL>|3101,3102
abscess|3102,3109
.|3109,3110
She|3111,3114
underwent|3115,3124
a|3125,3126
MRI|3127,3130
prior|3131,3136
surgery|3137,3144
for|3145,3148
operative|3149,3158
<EOL>|3159,3160
planning|3160,3168
.|3168,3169
She|3170,3173
underwent|3174,3183
a|3184,3185
right|3186,3191
craniotomy|3192,3202
and|3203,3206
evacuation|3207,3217
of|3218,3220
<EOL>|3221,3222
abscess|3222,3229
on|3230,3232
_|3233,3234
_|3234,3235
_|3235,3236
.|3236,3237
She|3238,3241
tolerated|3242,3251
the|3252,3255
procedure|3256,3265
well|3266,3270
and|3271,3274
was|3275,3278
<EOL>|3279,3280
extubated|3280,3289
in|3290,3292
the|3293,3296
operating|3297,3306
room|3307,3311
.|3311,3312
She|3313,3316
was|3317,3320
then|3321,3325
transferred|3326,3337
to|3338,3340
the|3341,3344
<EOL>|3345,3346
ICU|3346,3349
for|3350,3353
recovery|3354,3362
.|3362,3363
She|3364,3367
underwent|3368,3377
a|3378,3379
post-operative|3380,3394
non-contrasat|3395,3408
<EOL>|3409,3410
head|3410,3414
CT|3415,3417
which|3418,3423
revealed|3424,3432
normal|3433,3439
post|3440,3444
operative|3445,3454
changes|3455,3462
and|3463,3466
no|3467,3469
new|3470,3473
<EOL>|3474,3475
hemorrahge|3475,3485
.|3485,3486
<EOL>|3487,3488
<EOL>|3488,3489
On|3489,3491
_|3492,3493
_|3493,3494
_|3494,3495
,|3495,3496
she|3497,3500
was|3501,3504
sitting|3505,3512
in|3513,3515
the|3516,3519
chair|3520,3525
,|3525,3526
hemodynamically|3527,3542
and|3543,3546
<EOL>|3547,3548
neurologically|3548,3562
intact|3563,3569
.|3569,3570
She|3571,3574
transfered|3575,3585
to|3586,3588
the|3589,3592
floor|3593,3598
in|3599,3601
stable|3602,3608
<EOL>|3609,3610
conditions|3610,3620
.|3620,3621
<EOL>|3622,3623
<EOL>|3623,3624
Mrs.|3624,3628
_|3629,3630
_|3630,3631
_|3631,3632
was|3633,3636
followed|3637,3645
by|3646,3648
Infectious|3649,3659
Disease|3660,3667
.|3667,3668
They|3670,3674
<EOL>|3675,3676
recommended|3676,3687
that|3688,3692
the|3693,3696
patient|3697,3704
be|3705,3707
started|3708,3715
on|3716,3718
vancomycin|3719,3729
and|3730,3733
<EOL>|3734,3735
meropenem|3735,3744
until|3745,3750
culture|3751,3758
data|3759,3763
from|3764,3768
her|3769,3772
head|3773,3777
wound|3778,3783
was|3784,3787
obtained|3788,3796
.|3796,3797
<EOL>|3799,3800
<EOL>|3800,3801
On|3801,3803
_|3804,3805
_|3805,3806
_|3806,3807
,|3807,3808
cultures|3809,3817
revealed|3818,3826
no|3827,3829
growth|3830,3836
.|3836,3837
The|3838,3841
patient|3842,3849
was|3850,3853
continued|3854,3863
<EOL>|3864,3865
on|3865,3867
Vancomycin|3868,3878
,|3878,3879
meropenem|3880,3889
was|3890,3893
changed|3894,3901
to|3902,3904
ertapenum|3905,3914
.|3914,3915
<EOL>|3915,3916
<EOL>|3916,3917
The|3917,3920
patient|3921,3928
continued|3929,3938
to|3939,3941
progress|3942,3950
well|3951,3955
,|3955,3956
although|3957,3965
she|3966,3969
had|3970,3973
some|3974,3978
<EOL>|3979,3980
residual|3980,3988
left|3989,3993
-|3993,3994
sided|3994,3999
weakness|4000,4008
.|4008,4009
She|4011,4014
also|4015,4019
complained|4020,4030
of|4031,4033
some|4034,4038
<EOL>|4039,4040
left|4040,4044
-|4044,4045
handed|4045,4051
numbness|4052,4060
and|4061,4064
pain|4065,4069
.|4069,4070
<EOL>|4072,4073
<EOL>|4073,4074
On|4074,4076
_|4077,4078
_|4078,4079
_|4079,4080
,|4080,4081
the|4082,4085
patient|4086,4093
had|4094,4097
a|4098,4099
MR|4100,4102
head|4103,4107
with|4108,4112
and|4113,4116
without|4117,4124
contrast|4125,4133
<EOL>|4134,4135
including|4135,4144
DWI|4145,4148
,|4148,4149
which|4150,4155
showed|4156,4162
slight|4163,4169
improvement|4170,4181
.|4181,4182
She|4183,4186
was|4187,4190
<EOL>|4191,4192
discharged|4192,4202
home|4203,4207
on|4208,4210
_|4211,4212
_|4212,4213
_|4213,4214
with|4215,4219
appropriate|4220,4231
follow|4232,4238
-|4238,4239
up|4239,4241
,|4241,4242
and|4243,4246
all|4247,4250
<EOL>|4251,4252
questions|4252,4261
were|4262,4266
answered|4267,4275
before|4276,4282
discharge|4283,4292
.|4292,4293
<EOL>|4293,4294
<EOL>|4295,4296
Medications|4296,4307
on|4308,4310
Admission|4311,4320
:|4320,4321
<EOL>|4321,4322
The|4322,4325
Preadmission|4326,4338
Medication|4339,4349
list|4350,4354
is|4355,4357
accurate|4358,4366
and|4367,4370
complete|4371,4379
.|4379,4380
<EOL>|4380,4381
1.|4381,4383
CeftriaXONE|4384,4395
1|4396,4397
gm|4398,4400
IV|4401,4403
Q12H|4404,4408
<EOL>|4409,4410
2.|4410,4412
MetRONIDAZOLE|4413,4426
(|4427,4428
FLagyl|4428,4434
)|4434,4435
500|4436,4439
mg|4440,4442
PO|4443,4445
TID|4446,4449
<EOL>|4450,4451
3.|4451,4453
OxycoDONE|4454,4463
(|4464,4465
Immediate|4465,4474
Release|4475,4482
)|4482,4483
5|4485,4486
mg|4487,4489
PO|4490,4492
Q6H|4493,4496
:|4496,4497
PRN|4497,4500
pain|4501,4505
<EOL>|4506,4507
4.|4507,4509
Acetaminophen|4510,4523
325|4524,4527
-|4527,4528
650|4528,4531
mg|4532,4534
PO|4535,4537
Q6H|4538,4541
:|4541,4542
PRN|4542,4545
pain|4546,4550
<EOL>|4551,4552
5.|4552,4554
LeVETiracetam|4555,4568
1000|4569,4573
mg|4574,4576
PO|4577,4579
BID|4580,4583
<EOL>|4584,4585
<EOL>|4585,4586
<EOL>|4587,4588
Discharge|4588,4597
Disposition|4598,4609
:|4609,4610
<EOL>|4610,4611
Home|4611,4615
With|4616,4620
Service|4621,4628
<EOL>|4628,4629
<EOL>|4630,4631
Facility|4631,4639
:|4639,4640
<EOL>|4640,4641
_|4641,4642
_|4642,4643
_|4643,4644
<EOL>|4644,4645
<EOL>|4646,4647
Discharge|4647,4656
Diagnosis|4657,4666
:|4666,4667
<EOL>|4667,4668
Brain|4668,4673
Abscess|4674,4681
<EOL>|4681,4682
<EOL>|4683,4684
Mental|4705,4711
Status|4712,4718
:|4718,4719
Clear|4720,4725
and|4726,4729
coherent|4730,4738
.|4738,4739
<EOL>|4739,4740
Level|4740,4745
of|4746,4748
Consciousness|4749,4762
:|4762,4763
Alert|4764,4769
and|4770,4773
interactive|4774,4785
.|4785,4786
<EOL>|4786,4787
Activity|4787,4795
Status|4796,4802
:|4802,4803
Ambulatory|4804,4814
-|4815,4816
Independent|4817,4828
.|4828,4829
<EOL>|4829,4830
<EOL>|4830,4831
<EOL>|4832,4833
|4857,4858
Your|4858,4862
staples|4863,4870
should|4871,4877
stay|4878,4882
clean|4883,4888
and|4889,4892
dry|4893,4896
until|4897,4902
they|4903,4907
are|4908,4911
removed|4912,4919
.|4919,4920
<EOL>|4921,4922
<EOL>|4922,4923
|4923,4924
Have|4924,4928
a|4929,4930
friend|4931,4937
or|4938,4940
family|4941,4947
member|4948,4954
check|4955,4960
the|4961,4964
wound|4965,4970
for|4971,4974
signs|4975,4980
of|4981,4983
<EOL>|4984,4985
infection|4985,4994
such|4995,4999
as|5000,5002
redness|5003,5010
or|5011,5013
drainage|5014,5022
daily|5023,5028
.|5028,5029
<EOL>|5030,5031
|5031,5032
Take|5032,5036
your|5037,5041
pain|5042,5046
medicine|5047,5055
as|5056,5058
prescribed|5059,5069
if|5070,5072
needed|5073,5079
.|5079,5080
You|5081,5084
do|5085,5087
not|5088,5091
<EOL>|5092,5093
need|5093,5097
to|5098,5100
take|5101,5105
it|5106,5108
if|5109,5111
you|5112,5115
do|5116,5118
not|5119,5122
have|5123,5127
pain|5128,5132
.|5132,5133
<EOL>|5133,5134
|5134,5135
Exercise|5135,5143
should|5144,5150
be|5151,5153
limited|5154,5161
to|5162,5164
walking|5165,5172
;|5172,5173
no|5174,5176
lifting|5177,5184
>|5185,5186
10lbs|5186,5191
,|5191,5192
<EOL>|5193,5194
straining|5194,5203
,|5203,5204
or|5205,5207
excessive|5208,5217
bending|5218,5225
.|5225,5226
<EOL>|5226,5227
|5227,5228
Increase|5228,5236
your|5237,5241
intake|5242,5248
of|5249,5251
fluids|5252,5258
and|5259,5262
fiber|5263,5268
,|5268,5269
as|5270,5272
narcotic|5273,5281
pain|5282,5286
<EOL>|5287,5288
medicine|5288,5296
can|5297,5300
cause|5301,5306
constipation|5307,5319
.|5319,5320
We|5321,5323
generally|5324,5333
recommend|5334,5343
taking|5344,5350
<EOL>|5351,5352
an|5352,5354
over|5355,5359
the|5360,5363
counter|5364,5371
stool|5372,5377
softener|5378,5386
,|5386,5387
such|5388,5392
as|5393,5395
Docusate|5396,5404
(|5405,5406
Colace|5406,5412
)|5412,5413
<EOL>|5414,5415
while|5415,5420
taking|5421,5427
narcotic|5428,5436
pain|5437,5441
medication|5442,5452
.|5452,5453
<EOL>|5453,5454
|5454,5455
DO|5455,5457
not|5458,5461
take|5462,5466
any|5467,5470
anti-inflammatory|5471,5488
medicines|5489,5498
such|5499,5503
as|5504,5506
Motrin|5507,5513
,|5513,5514
<EOL>|5515,5516
Aspirin|5516,5523
,|5523,5524
Advil|5525,5530
,|5530,5531
or|5532,5534
Ibuprofen|5535,5544
etc.|5545,5549
until|5550,5555
follow|5556,5562
up|5563,5565
.|5565,5566
<EOL>|5566,5567
|5568,5569
You|5569,5572
have|5573,5577
been|5578,5582
discharged|5583,5593
on|5594,5596
Keppra|5597,5603
(|5604,5605
Levetiracetam|5605,5618
)|5618,5619
for|5620,5623
<EOL>|5624,5625
anti-seizure|5625,5637
medicine|5638,5646
;|5646,5647
you|5648,5651
will|5652,5656
not|5657,5660
require|5661,5668
blood|5669,5674
work|5675,5679
<EOL>|5680,5681
monitoring|5681,5691
.|5691,5692
<EOL>|5692,5693
|5693,5694
Do|5694,5696
not|5697,5700
drive|5701,5706
until|5707,5712
your|5713,5717
follow|5718,5724
up|5725,5727
appointment|5728,5739
.|5739,5740
<EOL>|5740,5741
<EOL>|5741,5742
<EOL>|5743,5744
Followup|5744,5752
Instructions|5753,5765
:|5765,5766
<EOL>|5766,5767
_|5767,5768
_|5768,5769
_|5769,5770
<EOL>|5770,5771

