 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|25,29
No|30,32
:|32,33
_|36,37
_|37,38
_|38,39
<EOL>|39,40
<EOL>|41,42
Admission|42,51
Date|52,56
:|56,57
_|59,60
_|60,61
_|61,62
Discharge|76,85
Date|86,90
:|90,91
_|94,95
_|95,96
_|96,97
<EOL>|97,98
<EOL>|99,100
Date|100,104
of|105,107
Birth|108,113
:|113,114
_|116,117
_|117,118
_|118,119
Sex|132,135
:|135,136
F|139,140
<EOL>|140,141
<EOL>|142,143
Service|143,150
:|150,151
MEDICINE|152,160
<EOL>|160,161
<EOL>|162,163
No|175,177
Known|178,183
Allergies|184,193
/|194,195
Adverse|196,203
Drug|204,208
Reactions|209,218
<EOL>|218,219
<EOL>|220,221
Attending|221,230
:|230,231
_|232,233
_|233,234
_|234,235
.|235,236
<EOL>|236,237
<EOL>|238,239
Chest|256,261
Pain|262,266
<EOL>|268,269
<EOL>|270,271
Major|271,276
Surgical|277,285
or|286,288
Invasive|289,297
Procedure|298,307
:|307,308
<EOL>|308,309
None|309,313
<EOL>|313,314
<EOL>|314,315
<EOL>|316,317
Ms.|346,349
_|350,351
_|351,352
_|352,353
is|354,356
a|357,358
_|359,360
_|360,361
_|361,362
y|363,364
/|364,365
o|365,366
female|367,373
with|374,378
a|379,380
history|381,388
of|389,391
<EOL>|392,393
hypertension|393,405
,|405,406
asthma|407,413
and|414,417
recent|418,424
diagnosis|425,434
of|435,437
CAD|438,441
based|442,447
on|448,450
stress|451,457
<EOL>|458,459
echo|459,463
done|464,468
on|469,471
_|472,473
_|473,474
_|474,475
,|475,476
thought|477,484
to|485,487
be|488,490
single|491,497
vessel|498,504
disease|505,512
who|513,516
<EOL>|517,518
presents|518,526
with|527,531
intermittent|532,544
chest|545,550
pain|551,555
since|556,561
her|562,565
recent|566,572
discharge|573,582
<EOL>|583,584
on|584,586
_|587,588
_|588,589
_|589,590
.|590,591
During|592,598
her|599,602
recent|603,609
hospitalization|610,625
she|626,629
was|630,633
ruled|634,639
out|640,643
<EOL>|644,645
for|645,648
an|649,651
MI|652,654
with|655,659
three|660,665
negative|666,674
sets|675,679
of|680,682
cardiac|683,690
enzymes|691,698
,|698,699
she|700,703
had|704,707
a|708,709
<EOL>|710,711
stress|711,717
echo|718,722
which|723,728
showed|729,735
inducible|736,745
ischemia|746,754
at|755,757
the|758,761
achieved|762,770
<EOL>|771,772
workload|772,780
,|780,781
thought|782,789
to|790,792
be|793,795
single|796,802
vessel|803,809
disease|810,817
per|818,821
the|822,825
echo|826,830
<EOL>|831,832
report|832,838
.|838,839
At|840,842
that|843,847
time|848,852
the|853,856
plan|857,861
was|862,865
for|866,869
medical|870,877
management|878,888
,|888,889
given|890,895
<EOL>|896,897
her|897,900
severe|901,907
underlying|908,918
pulmonary|919,928
disease|929,936
she|937,940
was|941,944
not|945,948
started|949,956
on|957,959
a|960,961
<EOL>|962,963
beta|963,967
blocker|968,975
,|975,976
but|977,980
was|981,984
started|985,992
on|993,995
diltiazem|996,1005
120mg|1006,1011
daily|1012,1017
.|1017,1018
Also|1019,1023
<EOL>|1024,1025
during|1025,1031
that|1032,1036
admission|1037,1046
she|1047,1050
was|1051,1054
found|1055,1060
to|1061,1063
have|1064,1068
intermittent|1069,1081
<EOL>|1082,1083
episodes|1083,1091
of|1092,1094
MAT|1095,1098
.|1098,1099
Today|1100,1105
she|1106,1109
was|1110,1113
on|1114,1116
the|1117,1120
phone|1121,1126
with|1127,1131
her|1132,1135
_|1136,1137
_|1137,1138
_|1138,1139
year|1140,1144
<EOL>|1145,1146
old|1146,1149
aunt|1150,1154
,|1154,1155
who|1156,1159
is|1160,1162
very|1163,1167
hard|1168,1172
or|1173,1175
hearing|1176,1183
,|1183,1184
she|1185,1188
says|1189,1193
that|1194,1198
she|1199,1202
became|1203,1209
<EOL>|1210,1211
frustrated|1211,1221
when|1222,1226
her|1227,1230
aunt|1231,1235
was|1236,1239
_|1240,1241
_|1241,1242
_|1242,1243
to|1244,1246
hear|1247,1251
her|1252,1255
on|1256,1258
the|1259,1262
phone|1263,1268
and|1269,1272
<EOL>|1273,1274
she|1274,1277
started|1278,1285
to|1286,1288
have|1289,1293
some|1294,1298
chest|1299,1304
pain|1305,1309
.|1309,1310
The|1311,1314
pain|1315,1319
began|1320,1325
in|1326,1328
the|1329,1332
<EOL>|1333,1334
_|1334,1335
_|1335,1336
_|1336,1337
her|1338,1341
chest|1342,1347
,|1347,1348
as|1349,1351
a|1352,1353
dull|1354,1358
pain|1359,1363
then|1364,1368
moved|1369,1374
up|1375,1377
to|1378,1380
her|1381,1384
left|1385,1389
<EOL>|1390,1391
shoulder|1391,1399
and|1400,1403
under|1404,1409
her|1410,1413
left|1414,1418
breast|1419,1425
,|1425,1426
at|1427,1429
its|1430,1433
worst|1434,1439
was|1440,1443
a|1444,1445
_|1446,1447
_|1447,1448
_|1448,1449
.|1449,1450
<EOL>|1451,1452
She|1452,1455
took|1456,1460
three|1461,1466
SL|1467,1469
nitro|1470,1475
's|1475,1477
at|1478,1480
home|1481,1485
,|1485,1486
with|1487,1491
some|1492,1496
minor|1497,1502
improvement|1503,1514
<EOL>|1515,1516
in|1516,1518
her|1519,1522
CP|1523,1525
but|1526,1529
when|1530,1534
it|1535,1537
did|1538,1541
not|1542,1545
resolve|1546,1553
she|1554,1557
called|1558,1564
Dr.|1565,1568
_|1569,1570
_|1570,1571
_|1571,1572
<EOL>|1573,1574
referred|1574,1582
her|1583,1586
to|1587,1589
the|1590,1593
ER|1594,1596
.|1596,1597
She|1598,1601
denied|1602,1608
any|1609,1612
associated|1613,1623
SOB|1624,1627
,|1627,1628
<EOL>|1629,1630
nausea|1630,1636
/|1636,1637
vomiting|1637,1645
.|1645,1646
She|1647,1650
denies|1651,1657
any|1658,1661
orthopnea|1662,1671
,|1671,1672
PND|1673,1676
,|1676,1677
_|1678,1679
_|1679,1680
_|1680,1681
edema|1682,1687
or|1688,1690
<EOL>|1691,1692
palpitations|1692,1704
.|1704,1705
<EOL>|1707,1708
.|1708,1709
<EOL>|1711,1712
In|1712,1714
the|1715,1718
ED|1719,1721
,|1721,1722
initial|1723,1730
vitals|1731,1737
were|1738,1742
98.7|1743,1747
,|1747,1748
73|1749,1751
,|1751,1752
183|1753,1756
/|1756,1757
92|1757,1759
,|1759,1760
20|1761,1763
,|1763,1764
98|1765,1767
%|1767,1768
on|1769,1771
RA|1772,1774
.|1774,1775
<EOL>|1776,1777
Her|1777,1780
EKG|1781,1784
had|1785,1788
a|1789,1790
LBBB|1791,1795
that|1796,1800
was|1801,1804
unchanged|1805,1814
from|1815,1819
prior|1820,1825
,|1825,1826
CXR|1827,1830
with|1831,1835
no|1836,1838
<EOL>|1839,1840
acute|1840,1845
process|1846,1853
.|1853,1854
Patient|1855,1862
given|1863,1868
aspirin|1869,1876
243mg|1877,1882
since|1883,1888
she|1889,1892
had|1893,1896
already|1897,1904
<EOL>|1905,1906
taken|1906,1911
81mg|1912,1916
of|1917,1919
aspirin|1920,1927
at|1928,1930
home|1931,1935
.|1935,1936
She|1937,1940
was|1941,1944
not|1945,1948
given|1949,1954
anything|1955,1963
for|1964,1967
<EOL>|1968,1969
her|1969,1972
episodes|1973,1981
of|1982,1984
chest|1985,1990
pain|1991,1995
as|1996,1998
they|1999,2003
resolved|2004,2012
without|2013,2020
further|2021,2028
<EOL>|2029,2030
intervention|2030,2042
.|2042,2043
Vitals|2044,2050
on|2051,2053
transfer|2054,2062
were|2063,2067
71|2068,2070
,|2070,2071
121|2072,2075
/|2075,2076
56|2076,2078
,|2078,2079
22|2080,2082
,|2082,2083
100|2084,2087
%|2087,2088
on|2089,2091
<EOL>|2092,2093
RA|2093,2095
.|2095,2096
<EOL>|2098,2099
.|2099,2100
<EOL>|2102,2103
On|2103,2105
arrival|2106,2113
to|2114,2116
the|2117,2120
floor|2121,2126
,|2126,2127
patient|2128,2135
's|2135,2137
initial|2138,2145
VS|2146,2148
were|2149,2153
:|2153,2154
98.9|2155,2159
,|2159,2160
<EOL>|2161,2162
140|2162,2165
/|2165,2166
86|2166,2168
,|2168,2169
68|2170,2172
,|2172,2173
18|2174,2176
,|2176,2177
97|2178,2180
%|2180,2181
on|2182,2184
RA|2185,2187
.|2187,2188
She|2189,2192
says|2193,2197
that|2198,2202
she|2203,2206
currently|2207,2216
may|2217,2220
have|2221,2225
<EOL>|2226,2227
a|2227,2228
little|2229,2235
bit|2236,2239
of|2240,2242
cental|2243,2249
CP|2250,2252
,|2252,2253
but|2254,2257
otherwise|2258,2267
feels|2268,2273
well|2274,2278
and|2279,2282
has|2283,2286
no|2287,2289
<EOL>|2290,2291
complaints|2291,2301
.|2301,2302
<EOL>|2304,2305
<EOL>|2306,2307
HTN|2329,2332
<EOL>|2334,2335
Asthma|2335,2341
<EOL>|2343,2344
Diverticulitis|2344,2358
several|2359,2366
years|2367,2372
ago|2373,2376
<EOL>|2378,2379
R|2379,2380
hip|2381,2384
replacement|2385,2396
in|2397,2399
_|2400,2401
_|2401,2402
_|2402,2403
<EOL>|2405,2406
Exertional|2406,2416
Atypical|2417,2425
Chest|2426,2431
Pain|2432,2436
<EOL>|2436,2437
<EOL>|2438,2439
:|2453,2454
<EOL>|2454,2455
_|2455,2456
_|2456,2457
_|2457,2458
<EOL>|2458,2459
:|2473,2474
<EOL>|2474,2475
Mother|2475,2481
:|2481,2482
_|2483,2484
_|2484,2485
_|2485,2486
,|2486,2487
HTN|2488,2491
<EOL>|2493,2494
Father|2494,2500
:|2500,2501
_|2502,2503
_|2503,2504
_|2504,2505
CA|2506,2508
<EOL>|2510,2511
Brother|2511,2518
:|2518,2519
CA|2520,2522
?|2522,2523
<EOL>|2525,2526
Brother|2526,2533
:|2533,2534
_|2535,2536
_|2536,2537
_|2537,2538
<EOL>|2540,2541
<EOL>|2541,2542
<EOL>|2543,2544
Physical|2544,2552
_|2553,2554
_|2554,2555
_|2555,2556
:|2556,2557
<EOL>|2557,2558
On|2558,2560
Admission|2561,2570
:|2570,2571
<EOL>|2571,2572
VS|2572,2574
:|2574,2575
T|2576,2577
=|2577,2578
98.9|2578,2582
BP|2583,2585
=|2585,2586
140|2586,2589
/|2589,2590
86|2590,2592
HR|2593,2595
=|2595,2596
68|2596,2598
RR|2599,2601
=|2601,2602
18|2602,2604
O2|2605,2607
sat|2608,2611
=|2611,2612
97|2612,2614
%|2614,2615
on|2616,2618
RA|2619,2621
<EOL>|2623,2624
GENERAL|2624,2631
:|2631,2632
WDWN|2633,2637
female|2638,2644
in|2645,2647
NAD|2648,2651
.|2651,2652
Oriented|2653,2661
x3|2662,2664
.|2664,2665
Mood|2666,2670
,|2670,2671
affect|2672,2678
<EOL>|2679,2680
appropriate|2680,2691
.|2691,2692
<EOL>|2694,2695
HEENT|2695,2700
:|2700,2701
NCAT|2702,2706
.|2706,2707
Sclera|2708,2714
anicteric|2715,2724
.|2724,2725
Conjunctiva|2726,2737
were|2738,2742
pink|2743,2747
,|2747,2748
no|2749,2751
pallor|2752,2758
<EOL>|2759,2760
or|2760,2762
cyanosis|2763,2771
of|2772,2774
the|2775,2778
oral|2779,2783
mucosa|2784,2790
.|2790,2791
No|2792,2794
xanthalesma|2795,2806
.|2806,2807
<EOL>|2809,2810
NECK|2810,2814
:|2814,2815
Supple|2816,2822
<EOL>|2824,2825
CARDIAC|2825,2832
:|2832,2833
RR|2834,2836
,|2836,2837
normal|2838,2844
S1|2845,2847
,|2847,2848
S2|2849,2851
.|2851,2852
No|2853,2855
m|2856,2857
/|2857,2858
r|2858,2859
/|2859,2860
g|2860,2861
.|2861,2862
No|2863,2865
thrills|2866,2873
,|2873,2874
lifts|2875,2880
.|2880,2881
No|2882,2884
S3|2885,2887
<EOL>|2888,2889
or|2889,2891
S4|2892,2894
.|2894,2895
<EOL>|2897,2898
LUNGS|2898,2903
:|2903,2904
No|2905,2907
chest|2908,2913
wall|2914,2918
deformities|2919,2930
,|2930,2931
scoliosis|2932,2941
or|2942,2944
kyphosis|2945,2953
.|2953,2954
Resp|2955,2959
<EOL>|2960,2961
were|2961,2965
unlabored|2966,2975
,|2975,2976
no|2977,2979
accessory|2980,2989
muscle|2990,2996
use|2997,3000
.|3000,3001
decreased|3002,3011
breath|3012,3018
sounds|3019,3025
<EOL>|3026,3027
throughout|3027,3037
,|3037,3038
although|3039,3047
CTA|3048,3051
,|3051,3052
no|3053,3055
crackles|3056,3064
,|3064,3065
wheezes|3066,3073
or|3074,3076
rhonchi|3077,3084
.|3084,3085
<EOL>|3087,3088
ABDOMEN|3088,3095
:|3095,3096
Soft|3097,3101
,|3101,3102
NTND|3103,3107
.|3107,3108
No|3109,3111
tenderness|3112,3122
.|3122,3123
<EOL>|3125,3126
EXTREMITIES|3126,3137
:|3137,3138
No|3139,3141
c|3142,3143
/|3143,3144
c|3144,3145
/|3145,3146
e|3146,3147
.|3147,3148
<EOL>|3150,3151
SKIN|3151,3155
:|3155,3156
No|3157,3159
stasis|3160,3166
dermatitis|3167,3177
,|3177,3178
ulcers|3179,3185
,|3185,3186
scars|3187,3192
,|3192,3193
or|3194,3196
xanthomas|3197,3206
.|3206,3207
<EOL>|3209,3210
PULSES|3210,3216
:|3216,3217
<EOL>|3219,3220
Right|3220,3225
:|3225,3226
DP|3227,3229
2|3230,3231
+|3231,3232
_|3233,3234
_|3234,3235
_|3235,3236
2|3237,3238
+|3238,3239
<EOL>|3241,3242
Left|3242,3246
:|3246,3247
DP|3248,3250
2|3251,3252
+|3252,3253
_|3254,3255
_|3255,3256
_|3256,3257
2|3258,3259
+|3259,3260
<EOL>|3262,3263
<EOL>|3263,3264
<EOL>|3265,3266
Pertinent|3266,3275
Results|3276,3283
:|3283,3284
<EOL>|3284,3285
_|3285,3286
_|3286,3287
_|3287,3288
03|3289,3291
:|3291,3292
55PM|3292,3296
_|3299,3300
_|3300,3301
_|3301,3302
PTT|3303,3306
-|3306,3307
26.0|3307,3311
_|3312,3313
_|3313,3314
_|3314,3315
<EOL>|3315,3316
_|3316,3317
_|3317,3318
_|3318,3319
03|3320,3322
:|3322,3323
55PM|3323,3327
PLT|3330,3333
COUNT|3334,3339
-|3339,3340
215|3340,3343
<EOL>|3343,3344
_|3344,3345
_|3345,3346
_|3346,3347
03|3348,3350
:|3350,3351
55PM|3351,3355
NEUTS|3358,3363
-|3363,3364
53.2|3364,3368
_|3369,3370
_|3370,3371
_|3371,3372
MONOS|3373,3378
-|3378,3379
5.7|3379,3382
EOS|3383,3386
-|3386,3387
0.9|3387,3390
<EOL>|3391,3392
BASOS|3392,3397
-|3397,3398
0.5|3398,3401
<EOL>|3401,3402
_|3402,3403
_|3403,3404
_|3404,3405
03|3406,3408
:|3408,3409
55PM|3409,3413
WBC|3416,3419
-|3419,3420
5.6|3420,3423
RBC|3424,3427
-|3427,3428
4|3428,3429
.|3429,3430
66|3430,3432
HGB|3433,3436
-|3436,3437
13.2|3437,3441
HCT|3442,3445
-|3445,3446
39.4|3446,3450
MCV|3451,3454
-|3454,3455
85|3455,3457
<EOL>|3458,3459
MCH|3459,3462
-|3462,3463
28.3|3463,3467
MCHC|3468,3472
-|3472,3473
33.4|3473,3477
RDW|3478,3481
-|3481,3482
15.0|3482,3486
<EOL>|3486,3487
_|3487,3488
_|3488,3489
_|3489,3490
03|3491,3493
:|3493,3494
55PM|3494,3498
cTropnT|3501,3508
-|3508,3509
<|3509,3510
0|3510,3511
.|3511,3512
01|3512,3514
<EOL>|3514,3515
_|3515,3516
_|3516,3517
_|3517,3518
03|3519,3521
:|3521,3522
55PM|3522,3526
estGFR|3529,3535
-|3535,3536
Using|3536,3541
this|3542,3546
<EOL>|3546,3547
_|3547,3548
_|3548,3549
_|3549,3550
03|3551,3553
:|3553,3554
55PM|3554,3558
GLUCOSE|3561,3568
-|3568,3569
94|3569,3571
UREA|3572,3576
N|3577,3578
-|3578,3579
21|3579,3581
*|3581,3582
CREAT|3583,3588
-|3588,3589
0.9|3589,3592
SODIUM|3593,3599
-|3599,3600
138|3600,3603
<EOL>|3604,3605
POTASSIUM|3605,3614
-|3614,3615
4.0|3615,3618
CHLORIDE|3619,3627
-|3627,3628
100|3628,3631
TOTAL|3632,3637
CO2|3638,3641
-|3641,3642
27|3642,3644
ANION|3645,3650
GAP|3651,3654
-|3654,3655
15|3655,3657
<EOL>|3657,3658
_|3658,3659
_|3659,3660
_|3660,3661
04|3662,3664
:|3664,3665
04PM|3665,3669
GLUCOSE|3672,3679
-|3679,3680
91|3680,3682
K|3683,3684
+|3684,3685
-|3685,3686
4.1|3686,3689
<EOL>|3689,3690
_|3690,3691
_|3691,3692
_|3692,3693
12|3694,3696
:|3696,3697
00AM|3697,3701
CK|3704,3706
-|3706,3707
MB|3707,3709
-|3709,3710
3|3710,3711
cTropnT|3712,3719
-|3719,3720
<|3720,3721
0|3721,3722
.|3722,3723
01|3723,3725
<EOL>|3725,3726
_|3726,3727
_|3727,3728
_|3728,3729
12|3730,3732
:|3732,3733
00AM|3733,3737
CK|3740,3742
(|3742,3743
CPK|3743,3746
)|3746,3747
-|3747,3748
189|3748,3751
<EOL>|3751,3752
<EOL>|3752,3753
CXR|3753,3756
:|3756,3757
Emphysema|3758,3767
without|3768,3775
superimposed|3776,3788
pneumonia|3789,3798
or|3799,3801
CHF|3802,3805
.|3805,3806
<EOL>|3806,3807
<EOL>|3808,3809
ASSESSMENT|3832,3842
AND|3843,3846
PLAN|3847,3851
:|3851,3852
Ms|3853,3855
.|3855,3856
_|3857,3858
_|3858,3859
_|3859,3860
is|3861,3863
a|3864,3865
_|3866,3867
_|3867,3868
_|3868,3869
year|3870,3874
old|3875,3878
female|3879,3885
with|3886,3890
<EOL>|3891,3892
a|3892,3893
recent|3894,3900
diagnosis|3901,3910
of|3911,3913
CAD|3914,3917
,|3917,3918
HTN|3919,3922
and|3923,3926
asthma|3927,3933
who|3934,3937
presents|3938,3946
with|3947,3951
<EOL>|3952,3953
intermittent|3953,3965
episodes|3966,3974
of|3975,3977
chest|3978,3983
pain|3984,3988
since|3989,3994
her|3995,3998
recent|3999,4005
discharge|4006,4015
.|4015,4016
<EOL>|4018,4019
<EOL>|4019,4020
...|4020,4023
...|4023,4026
...|4026,4029
...|4029,4032
...|4032,4035
...|4035,4038
...|4038,4041
...|4041,4044
...|4044,4047
...|4047,4050
...|4050,4053
...|4053,4056
.|4056,4057
.|4057,4058
<EOL>|4058,4059
Active|4059,4065
Issues|4066,4072
:|4072,4073
<EOL>|4073,4074
.|4074,4075
<EOL>|4077,4078
#|4078,4079
CORONARIES|4080,4090
:|4090,4091
patient|4092,4099
with|4100,4104
intermittent|4105,4117
episodes|4118,4126
of|4127,4129
left|4130,4134
chest|4135,4140
<EOL>|4141,4142
burning|4142,4149
,|4149,4150
that|4151,4155
are|4156,4159
not|4160,4163
typical|4164,4171
of|4172,4174
angina|4175,4181
since|4182,4187
they|4188,4192
resolve|4193,4200
<EOL>|4201,4202
without|4202,4209
intervention|4210,4222
,|4222,4223
are|4224,4227
not|4228,4231
relieved|4232,4240
by|4241,4243
nitro|4244,4249
and|4250,4253
have|4254,4258
no|4259,4261
<EOL>|4262,4263
association|4263,4274
with|4275,4279
exercise|4280,4288
.|4288,4289
However|4290,4297
,|4297,4298
given|4299,4304
the|4305,4308
findings|4309,4317
on|4318,4320
her|4321,4324
<EOL>|4325,4326
recent|4326,4332
stress|4333,4339
echo|4340,4344
of|4345,4347
inducible|4348,4357
ischemia|4358,4366
it|4367,4369
is|4370,4372
concerning|4373,4383
that|4384,4388
<EOL>|4389,4390
her|4390,4393
current|4394,4401
symptoms|4402,4410
could|4411,4416
be|4417,4419
related|4420,4427
to|4428,4430
her|4431,4434
underlying|4435,4445
CAD|4446,4449
.|4449,4450
Her|4451,4454
<EOL>|4455,4456
troponins|4456,4465
were|4466,4470
negative|4471,4479
during|4480,4486
this|4487,4491
hospital|4492,4500
stay|4501,4505
.|4505,4506
On|4508,4510
this|4511,4515
<EOL>|4516,4517
admission|4517,4526
,|4526,4527
she|4528,4531
was|4532,4535
started|4536,4543
on|4544,4546
Imdur|4547,4552
30|4553,4555
in|4556,4558
addition|4559,4567
to|4568,4570
the|4571,4574
<EOL>|4575,4576
medications|4576,4587
started|4588,4595
on|4596,4598
last|4599,4603
discharge|4604,4613
as|4614,4616
it|4617,4619
was|4620,4623
decided|4624,4631
that|4632,4636
she|4637,4640
<EOL>|4641,4642
may|4642,4645
need|4646,4650
better|4651,4657
medical|4658,4665
management|4666,4676
prior|4677,4682
to|4683,4685
resorting|4686,4695
to|4696,4698
PCI|4699,4702
<EOL>|4703,4704
(|4704,4705
which|4705,4710
may|4711,4714
be|4715,4717
a|4718,4719
possibility|4720,4731
in|4732,4734
the|4735,4738
future|4739,4745
)|4745,4746
.|4746,4747
After|4748,4753
administration|4754,4768
<EOL>|4769,4770
of|4770,4772
IMDUR|4773,4778
,|4778,4779
we|4780,4782
walked|4783,4789
the|4790,4793
patient|4794,4801
down|4802,4806
the|4807,4810
hall|4811,4815
,|4815,4816
as|4817,4819
well|4820,4824
as|4825,4827
up|4828,4830
<EOL>|4831,4832
several|4832,4839
flights|4840,4847
of|4848,4850
stairs|4851,4857
.|4857,4858
She|4859,4862
denied|4863,4869
feeling|4870,4877
short|4878,4883
of|4884,4886
breath|4887,4893
,|4893,4894
<EOL>|4895,4896
nor|4896,4899
did|4900,4903
she|4904,4907
endorse|4908,4915
any|4916,4919
other|4920,4925
cardiac|4926,4933
symtpoms|4934,4942
,|4942,4943
such|4944,4948
as|4949,4951
chest|4952,4957
<EOL>|4958,4959
pain|4959,4963
.|4963,4964
In|4965,4967
fact|4968,4972
,|4972,4973
she|4974,4977
stated|4978,4984
that|4985,4989
she|4990,4993
felt|4994,4998
well|4999,5003
walking|5004,5011
.|5011,5012
<EOL>|5013,5014
.|5014,5015
<EOL>|5017,5018
#|5018,5019
RHYTHM|5020,5026
:|5026,5027
LBBB|5028,5032
on|5033,5035
EKG|5036,5039
from|5040,5044
yesterday|5045,5054
,|5054,5055
regular|5056,5063
.|5063,5064
patient|5065,5072
with|5073,5077
a|5078,5079
<EOL>|5080,5081
new|5081,5084
diagnosis|5085,5094
of|5095,5097
MAT|5098,5101
on|5102,5104
last|5105,5109
admission|5110,5119
.|5119,5120
We|5121,5123
continued|5124,5133
her|5134,5137
on|5138,5140
<EOL>|5141,5142
Diltiazem|5142,5151
.|5151,5152
She|5153,5156
had|5157,5160
several|5161,5168
episodes|5169,5177
of|5178,5180
MAT|5181,5184
on|5185,5187
tele|5188,5192
,|5192,5193
but|5194,5197
was|5198,5201
<EOL>|5202,5203
asymptomatic|5203,5215
.|5215,5216
Given|5217,5222
frequent|5223,5231
PAT|5232,5235
,|5235,5236
_|5237,5238
_|5238,5239
_|5239,5240
of|5241,5243
Hearts|5244,5250
monitor|5251,5258
was|5259,5262
<EOL>|5263,5264
arranged|5264,5272
for|5273,5276
her|5277,5280
on|5281,5283
discharge|5284,5293
to|5294,5296
exclude|5297,5304
the|5305,5308
possibility|5309,5320
that|5321,5325
<EOL>|5326,5327
symptoms|5327,5335
are|5336,5339
due|5340,5343
to|5344,5346
a|5347,5348
tachyarrhythmia|5349,5364
.|5364,5365
<EOL>|5366,5367
...|5367,5370
...|5370,5373
...|5373,5376
...|5376,5379
...|5379,5382
...|5382,5385
...|5385,5388
...|5388,5391
...|5391,5394
...|5394,5397
...|5397,5400
...|5400,5403
...|5403,5406
...|5406,5409
...|5409,5412
<EOL>|5412,5413
Inactive|5413,5421
Issues|5422,5428
:|5428,5429
<EOL>|5429,5430
#|5430,5431
Hypertension|5432,5444
:|5444,5445
continued|5446,5455
home|5456,5460
HCTZ|5461,5465
and|5466,5469
diltiazem|5470,5479
.|5479,5480
.|5480,5481
<EOL>|5483,5484
#|5484,5485
Asthma|5486,5492
:|5492,5493
continued|5493,5502
home|5503,5507
medications|5508,5519
.|5519,5520
<EOL>|5524,5525
#|5525,5526
GERD|5527,5531
:|5531,5532
continued|5533,5542
home|5543,5547
omeprazole|5548,5558
<EOL>|5560,5561
.|5561,5562
<EOL>|5566,5567
CODE|5567,5571
:|5571,5572
full|5573,5577
code|5578,5582
<EOL>|5584,5585
...|5585,5588
...|5588,5591
...|5591,5594
...|5594,5597
...|5597,5600
...|5600,5603
...|5603,5606
...|5606,5609
...|5609,5612
...|5612,5615
...|5615,5618
...|5618,5621
.|5621,5622
<EOL>|5624,5625
Transitional|5625,5637
Issues|5638,5644
:|5644,5645
<EOL>|5645,5646
1|5646,5647
)|5647,5648
Patient|5649,5656
was|5657,5660
started|5661,5668
on|5669,5671
Imdur|5672,5677
30mg|5678,5682
daily|5683,5688
in|5689,5691
additon|5692,5699
to|5700,5702
her|5703,5706
<EOL>|5707,5708
other|5708,5713
medications|5714,5725
.|5725,5726
She|5727,5730
is|5731,5733
being|5734,5739
medically|5740,5749
managed|5750,5757
for|5758,5761
her|5762,5765
<EOL>|5766,5767
coronary|5767,5775
artery|5776,5782
disease|5783,5790
but|5791,5794
may|5795,5798
be|5799,5801
a|5802,5803
candidate|5804,5813
for|5814,5817
PCI|5818,5821
in|5822,5824
the|5825,5828
<EOL>|5829,5830
future|5830,5836
if|5837,5839
the|5840,5843
symtpoms|5844,5852
of|5853,5855
chest|5856,5861
pain|5862,5866
return|5867,5873
.|5873,5874
<EOL>|5874,5875
2|5875,5876
)|5876,5877
Follow|5878,5884
-|5884,5885
up|5885,5887
event|5888,5893
monitor|5894,5901
for|5902,5905
evaluation|5906,5916
of|5917,5919
arrhythmias|5920,5931
<EOL>|5931,5932
<EOL>|5933,5934
Medications|5934,5945
on|5946,5948
Admission|5949,5958
:|5958,5959
<EOL>|5959,5960
-|5960,5961
acetaminophen|5961,5974
325|5975,5978
mg|5979,5981
Q4H|5982,5985
as|5986,5988
needed|5989,5995
for|5996,5999
pain|6000,6004
.|6004,6005
<EOL>|6007,6008
-|6008,6009
albuterol|6009,6018
sulfate|6019,6026
90|6027,6029
mcg|6030,6033
:|6033,6034
Two|6035,6038
(|6039,6040
2|6040,6041
)|6041,6042
Puff|6043,6047
Inhalation|6048,6058
Q6H|6059,6062
(|6063,6064
every|6064,6069
6|6070,6071
<EOL>|6072,6073
hours|6073,6078
)|6078,6079
as|6080,6082
needed|6083,6089
for|6090,6093
SOB|6094,6097
or|6098,6100
wheeze|6101,6107
.|6107,6108
<EOL>|6110,6111
-|6111,6112
fluticasone|6112,6123
-|6123,6124
salmeterol|6124,6134
500|6135,6138
-|6138,6139
50|6139,6141
mcg|6142,6145
:|6145,6146
Inhalation|6147,6157
BID|6158,6161
<EOL>|6163,6164
-|6164,6165
fluticasone|6165,6176
50|6177,6179
mcg|6180,6183
:|6183,6184
_|6185,6186
_|6186,6187
_|6187,6188
Nasal|6189,6194
once|6195,6199
a|6200,6201
day|6202,6205
<EOL>|6207,6208
-|6208,6209
hydrochlorothiazide|6209,6228
50|6229,6231
mg|6232,6234
once|6235,6239
a|6240,6241
day|6242,6245
.|6245,6246
<EOL>|6248,6249
-|6249,6250
omeprazole|6250,6260
20|6261,6263
mg|6264,6266
DAILY|6267,6272
<EOL>|6274,6275
-|6275,6276
simvastatin|6276,6287
20|6288,6290
mg|6291,6293
once|6294,6298
a|6299,6300
day|6301,6304
.|6304,6305
<EOL>|6307,6308
-|6308,6309
tiotropium|6309,6319
bromide|6320,6327
18|6328,6330
mcg|6331,6334
DAILY|6335,6340
<EOL>|6342,6343
-|6343,6344
aspirin|6344,6351
81|6352,6354
mg|6355,6357
once|6358,6362
a|6363,6364
day|6365,6368
.|6368,6369
<EOL>|6371,6372
-|6372,6373
multivitamin|6373,6385
1|6386,6387
Tablet|6388,6394
DAILY|6395,6400
<EOL>|6402,6403
-|6403,6404
diltiazem|6404,6413
HCl|6414,6417
120|6418,6421
mg|6422,6424
Tablet|6425,6431
Sustained|6432,6441
Release|6442,6449
24|6450,6452
hr|6453,6455
daily|6456,6461
<EOL>|6463,6464
-|6464,6465
singulair|6465,6474
10mg|6475,6479
QHS|6480,6483
<EOL>|6485,6486
<EOL>|6487,6488
Discharge|6488,6497
Medications|6498,6509
:|6509,6510
<EOL>|6510,6511
1.|6511,6513
acetaminophen|6514,6527
325|6528,6531
mg|6532,6534
Tablet|6535,6541
Sig|6542,6545
:|6545,6546
One|6547,6550
(|6551,6552
1|6552,6553
)|6553,6554
Tablet|6555,6561
PO|6562,6564
every|6565,6570
four|6571,6575
<EOL>|6576,6577
(|6577,6578
4|6578,6579
)|6579,6580
hours|6581,6586
as|6587,6589
needed|6590,6596
for|6597,6600
pain|6601,6605
.|6605,6606
<EOL>|6608,6609
2.|6609,6611
albuterol|6612,6621
sulfate|6622,6629
90|6630,6632
mcg|6633,6636
/|6636,6637
Actuation|6637,6646
HFA|6647,6650
Aerosol|6651,6658
Inhaler|6659,6666
Sig|6667,6670
:|6670,6671
<EOL>|6672,6673
Two|6673,6676
(|6677,6678
2|6678,6679
)|6679,6680
Puff|6681,6685
Inhalation|6686,6696
Q6H|6697,6700
(|6701,6702
every|6702,6707
6|6708,6709
hours|6710,6715
)|6715,6716
as|6717,6719
needed|6720,6726
for|6727,6730
sob|6731,6734
,|6734,6735
<EOL>|6736,6737
wheezing|6737,6745
.|6746,6747
<EOL>|6749,6750
3.|6750,6752
fluticasone|6753,6764
-|6764,6765
salmeterol|6765,6775
500|6776,6779
-|6779,6780
50|6780,6782
mcg|6783,6786
/|6786,6787
dose|6787,6791
Disk|6792,6796
with|6797,6801
Device|6802,6808
Sig|6809,6812
:|6812,6813
<EOL>|6814,6815
One|6815,6818
(|6819,6820
1|6820,6821
)|6821,6822
Disk|6823,6827
with|6828,6832
Device|6833,6839
Inhalation|6840,6850
BID|6851,6854
(|6855,6856
2|6856,6857
times|6858,6863
a|6864,6865
day|6866,6869
)|6869,6870
.|6870,6871
<EOL>|6873,6874
4.|6874,6876
fluticasone|6877,6888
50|6889,6891
mcg|6892,6895
/|6895,6896
Actuation|6896,6905
Spray|6906,6911
,|6911,6912
Suspension|6913,6923
Sig|6924,6927
:|6927,6928
One|6929,6932
(|6933,6934
1|6934,6935
)|6935,6936
<EOL>|6937,6938
Spray|6938,6943
Nasal|6944,6949
DAILY|6950,6955
(|6956,6957
Daily|6957,6962
)|6962,6963
.|6963,6964
<EOL>|6966,6967
5.|6967,6969
hydrochlorothiazide|6970,6989
12.5|6990,6994
mg|6995,6997
Capsule|6998,7005
Sig|7006,7009
:|7009,7010
One|7011,7014
(|7015,7016
1|7016,7017
)|7017,7018
Capsule|7019,7026
PO|7027,7029
<EOL>|7030,7031
once|7031,7035
a|7036,7037
day|7038,7041
.|7041,7042
<EOL>|7044,7045
6.|7045,7047
omeprazole|7048,7058
20|7059,7061
mg|7062,7064
Capsule|7065,7072
,|7072,7073
Delayed|7074,7081
Release|7082,7089
(|7089,7090
E.C|7090,7093
.|7093,7094
)|7094,7095
Sig|7096,7099
:|7099,7100
One|7101,7104
(|7105,7106
1|7106,7107
)|7107,7108
<EOL>|7109,7110
Capsule|7110,7117
,|7117,7118
Delayed|7119,7126
Release|7127,7134
(|7134,7135
E.C|7135,7138
.|7138,7139
)|7139,7140
PO|7141,7143
DAILY|7144,7149
(|7150,7151
Daily|7151,7156
)|7156,7157
.|7157,7158
<EOL>|7160,7161
7.|7161,7163
simvastatin|7164,7175
20|7176,7178
mg|7179,7181
Tablet|7182,7188
Sig|7189,7192
:|7192,7193
One|7194,7197
(|7198,7199
1|7199,7200
)|7200,7201
Tablet|7202,7208
PO|7209,7211
once|7212,7216
a|7217,7218
day|7219,7222
.|7222,7223
<EOL>|7225,7226
8.|7226,7228
tiotropium|7229,7239
bromide|7240,7247
18|7248,7250
mcg|7251,7254
Capsule|7255,7262
,|7262,7263
w|7264,7265
/|7265,7266
Inhalation|7266,7276
Device|7277,7283
Sig|7284,7287
:|7287,7288
<EOL>|7289,7290
One|7290,7293
(|7294,7295
1|7295,7296
)|7296,7297
Cap|7298,7301
Inhalation|7302,7312
DAILY|7313,7318
(|7319,7320
Daily|7320,7325
)|7325,7326
.|7326,7327
<EOL>|7329,7330
9.|7330,7332
aspirin|7333,7340
81|7341,7343
mg|7344,7346
Tablet|7347,7353
Sig|7354,7357
:|7357,7358
One|7359,7362
(|7363,7364
1|7364,7365
)|7365,7366
Tablet|7367,7373
PO|7374,7376
once|7377,7381
a|7382,7383
day|7384,7387
.|7387,7388
<EOL>|7390,7391
10.|7391,7394
multivitamin|7395,7407
Tablet|7412,7418
Sig|7419,7422
:|7422,7423
One|7424,7427
(|7428,7429
1|7429,7430
)|7430,7431
Tablet|7432,7438
PO|7439,7441
DAILY|7442,7447
<EOL>|7448,7449
(|7449,7450
Daily|7450,7455
)|7455,7456
.|7456,7457
<EOL>|7459,7460
11.|7460,7463
montelukast|7464,7475
10|7476,7478
mg|7479,7481
Tablet|7482,7488
Sig|7489,7492
:|7492,7493
One|7494,7497
(|7498,7499
1|7499,7500
)|7500,7501
Tablet|7502,7508
PO|7509,7511
QHS|7512,7515
(|7516,7517
once|7517,7521
a|7522,7523
<EOL>|7524,7525
day|7525,7528
(|7529,7530
at|7530,7532
bedtime|7533,7540
)|7540,7541
)|7541,7542
.|7542,7543
<EOL>|7545,7546
12.|7546,7549
isosorbide|7550,7560
mononitrate|7561,7572
30|7573,7575
mg|7576,7578
Tablet|7579,7585
Sustained|7586,7595
Release|7596,7603
24|7604,7606
hr|7607,7609
<EOL>|7610,7611
Sig|7611,7614
:|7614,7615
One|7616,7619
(|7620,7621
1|7621,7622
)|7622,7623
Tablet|7624,7630
Sustained|7631,7640
Release|7641,7648
24|7649,7651
hr|7652,7654
PO|7655,7657
once|7658,7662
a|7663,7664
day|7665,7668
.|7668,7669
<EOL>|7669,7670
Disp|7670,7674
:|7674,7675
*|7675,7676
30|7676,7678
Tablet|7679,7685
Sustained|7686,7695
Release|7696,7703
24|7704,7706
hr|7707,7709
(|7709,7710
s|7710,7711
)|7711,7712
*|7712,7713
Refills|7714,7721
:|7721,7722
*|7722,7723
2|7723,7724
*|7724,7725
<EOL>|7725,7726
13.|7726,7729
diltiazem|7730,7739
HCl|7740,7743
180|7744,7747
mg|7748,7750
Capsule|7751,7758
,|7758,7759
Sust|7760,7764
.|7764,7765
Release|7766,7773
24|7774,7776
hr|7777,7779
Sig|7780,7783
:|7783,7784
One|7785,7788
<EOL>|7789,7790
(|7790,7791
1|7791,7792
)|7792,7793
Capsule|7794,7801
,|7801,7802
Sust|7803,7807
.|7807,7808
Release|7809,7816
24|7817,7819
hr|7820,7822
PO|7823,7825
once|7826,7830
a|7831,7832
day|7833,7836
.|7836,7837
<EOL>|7837,7838
Disp|7838,7842
:|7842,7843
*|7843,7844
30|7844,7846
Capsule|7847,7854
,|7854,7855
Sust|7856,7860
.|7860,7861
Release|7862,7869
24|7870,7872
hr|7873,7875
(|7875,7876
s|7876,7877
)|7877,7878
*|7878,7879
Refills|7880,7887
:|7887,7888
*|7888,7889
2|7889,7890
*|7890,7891
<EOL>|7891,7892
<EOL>|7892,7893
<EOL>|7894,7895
Discharge|7895,7904
Disposition|7905,7916
:|7916,7917
<EOL>|7917,7918
Home|7918,7922
<EOL>|7922,7923
<EOL>|7924,7925
Discharge|7925,7934
Diagnosis|7935,7944
:|7944,7945
<EOL>|7945,7946
PRIMARY|7946,7953
:|7953,7954
<EOL>|7954,7955
1.|7955,7957
atypical|7958,7966
chest|7967,7972
pain|7973,7977
<EOL>|7977,7978
<EOL>|7978,7979
Secondary|7979,7988
:|7988,7989
<EOL>|7990,7991
1.|7991,7993
Hypertension|7994,8006
<EOL>|8006,8007
2.|8007,8009
Asthma|8010,8016
<EOL>|8016,8017
3.|8017,8019
Diverticulitis|8020,8034
<EOL>|8034,8035
<EOL>|8035,8036
<EOL>|8037,8038
Mental|8059,8065
Status|8066,8072
:|8072,8073
Clear|8074,8079
and|8080,8083
coherent|8084,8092
.|8092,8093
<EOL>|8093,8094
Level|8094,8099
of|8100,8102
Consciousness|8103,8116
:|8116,8117
Alert|8118,8123
and|8124,8127
interactive|8128,8139
.|8139,8140
<EOL>|8140,8141
Activity|8141,8149
Status|8150,8156
:|8156,8157
Ambulatory|8158,8168
-|8169,8170
Independent|8171,8182
.|8182,8183
<EOL>|8183,8184
<EOL>|8184,8185
<EOL>|8186,8187
You|8211,8214
were|8215,8219
admitted|8220,8228
to|8229,8231
the|8232,8235
hospital|8236,8244
for|8245,8248
atypical|8249,8257
chest|8258,8263
pain|8264,8268
.|8268,8269
You|8270,8273
<EOL>|8274,8275
were|8275,8279
monitored|8280,8289
on|8290,8292
telemetry|8293,8302
.|8302,8303
Your|8304,8308
EKG|8309,8312
was|8313,8316
unchanged|8317,8326
.|8326,8327
Your|8328,8332
<EOL>|8333,8334
cardiac|8334,8341
enzymes|8342,8349
were|8350,8354
normal|8355,8361
,|8361,8362
without|8363,8370
evidence|8371,8379
for|8380,8383
heart|8384,8389
damage|8390,8396
<EOL>|8397,8398
or|8398,8400
heart|8401,8406
attack|8407,8413
.|8413,8414
We|8415,8417
have|8418,8422
started|8423,8430
you|8431,8434
on|8435,8437
a|8438,8439
long|8440,8444
acting|8445,8451
nitrate|8452,8459
<EOL>|8460,8461
medication|8461,8471
to|8472,8474
control|8475,8482
your|8483,8487
chest|8488,8493
pain|8494,8498
symptoms|8499,8507
.|8507,8508
We|8509,8511
also|8512,8516
<EOL>|8517,8518
increased|8518,8527
your|8528,8532
diltiazem|8533,8542
for|8543,8546
better|8547,8553
blood|8554,8559
pressure|8560,8568
and|8569,8572
heart|8573,8578
<EOL>|8579,8580
rate|8580,8584
control|8585,8592
.|8592,8593
<EOL>|8593,8594
.|8594,8595
<EOL>|8595,8596
Finally|8596,8603
,|8603,8604
we|8605,8607
have|8608,8612
set|8613,8616
you|8617,8620
up|8621,8623
with|8624,8628
a|8629,8630
48|8631,8633
hour|8634,8638
holter|8639,8645
monitor|8646,8653
to|8654,8656
get|8657,8660
<EOL>|8661,8662
a|8662,8663
better|8664,8670
idea|8671,8675
of|8676,8678
your|8679,8683
heart|8684,8689
rhythm|8690,8696
over|8697,8701
time|8702,8706
.|8706,8707
Please|8708,8714
discuss|8715,8722
<EOL>|8723,8724
these|8724,8729
results|8730,8737
with|8738,8742
_|8743,8744
_|8744,8745
_|8745,8746
.|8746,8747
_|8748,8749
_|8749,8750
_|8750,8751
at|8752,8754
your|8755,8759
upcoming|8760,8768
<EOL>|8769,8770
cardiology|8770,8780
appointment|8781,8792
.|8792,8793
<EOL>|8793,8794
.|8794,8795
<EOL>|8795,8796
MEDICATION|8796,8806
CHANGES|8807,8814
:|8814,8815
<EOL>|8815,8816
-|8816,8817
START|8818,8823
imdur|8824,8829
30|8830,8832
mg|8833,8835
daily|8836,8841
<EOL>|8841,8842
-|8842,8843
INCREASE|8844,8852
diltiazem|8853,8862
to|8863,8865
180|8866,8869
mg|8870,8872
daily|8873,8878
<EOL>|8878,8879
.|8879,8880
<EOL>|8880,8881
Please|8881,8887
continue|8888,8896
your|8897,8901
other|8902,8907
medications|8908,8919
as|8920,8922
prescribed|8923,8933
.|8933,8934
<EOL>|8934,8935
.|8935,8936
<EOL>|8936,8937
Please|8937,8943
seek|8944,8948
medical|8949,8956
attention|8957,8966
for|8967,8970
worsening|8971,8980
chest|8981,8986
pain|8987,8991
,|8991,8992
<EOL>|8993,8994
shortness|8994,9003
of|9004,9006
breath|9007,9013
,|9013,9014
or|9015,9017
any|9018,9021
other|9022,9027
symptoms|9028,9036
.|9036,9037
<EOL>|9037,9038
<EOL>|9039,9040
Followup|9040,9048
Instructions|9049,9061
:|9061,9062
<EOL>|9062,9063
_|9063,9064
_|9064,9065
_|9065,9066
<EOL>|9066,9067

