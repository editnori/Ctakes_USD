 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|45,54|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|45,54|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|45,59|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|79,88|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|79,88|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|79,88|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|79,93|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|111,116|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|135,138|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|135,138|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|146,153|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|146,153|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Attribute|Clinical Attribute|Allergies|188,197|false|false|false|C1717415||Allergies
Event|Event|Allergies|188,197|false|false|false|||Allergies
Finding|Pathologic Function|Allergies|188,197|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|200,222|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|208,212|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|208,212|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|208,222|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Event|Event|Allergies|213,222|false|false|false|||Reactions
Event|Event|Allergies|225,234|false|false|false|||Attending
Finding|Functional Concept|Allergies|225,234|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|268,274|false|false|false|||speech
Finding|Organism Function|Chief Complaint|268,274|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Chief Complaint|268,274|false|false|false|C0846595|Speech assessment|speech
Finding|Classification|Chief Complaint|277,282|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|283,291|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|295,313|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|304,313|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|304,313|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|304,313|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|304,313|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|304,313|false|false|false|C0184661|Interventional procedure|Procedure
Finding|Idea or Concept|History of Present Illness|354,358|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|354,358|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Functional Concept|History of Present Illness|363,368|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|393,399|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|History of Present Illness|393,412|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|393,412|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|History of Present Illness|393,412|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|History of Present Illness|400,412|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|History of Present Illness|400,412|false|false|false|||fibrillation
Drug|Organic Chemical|History of Present Illness|417,424|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|History of Present Illness|417,424|false|false|false|C3530466|Eliquis|Eliquis
Event|Event|History of Present Illness|417,424|false|false|false|||Eliquis
Finding|Intellectual Product|History of Present Illness|431,435|false|false|false|C1720092|Once - dosing instruction fragment|once
Disorder|Disease or Syndrome|History of Present Illness|444,456|false|false|false|C0020538|Hypertensive disease|hypertension
Event|Event|History of Present Illness|444,456|false|false|false|||hypertension
Disorder|Disease or Syndrome|History of Present Illness|458,472|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|History of Present Illness|458,472|false|false|false|||hyperlipidemia
Finding|Finding|History of Present Illness|458,472|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Anatomy|Body Space or Junction|History of Present Illness|474,477|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|History of Present Illness|474,477|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|History of Present Illness|474,477|false|false|false|||CHF
Event|Event|History of Present Illness|478,486|false|false|false|||presents
Event|Event|History of Present Illness|490,498|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|490,498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|490,498|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|490,498|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|History of Present Illness|504,507|false|false|false|||OSH
Finding|Intellectual Product|History of Present Illness|522,527|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Intellectual Product|History of Present Illness|522,533|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|acute onset
Event|Event|History of Present Illness|528,533|false|false|false|||onset
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|535,545|false|false|false|C0013362|Dysarthria|dysarthria
Event|Event|History of Present Illness|535,545|false|false|false|||dysarthria
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|550,553|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|History of Present Illness|550,553|false|false|false|||CTA
Finding|Gene or Genome|History of Present Illness|550,553|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|History of Present Illness|550,553|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Event|Event|History of Present Illness|554,560|false|false|false|||showed
Finding|Finding|History of Present Illness|561,569|false|false|false|C0332149|Possible|possible
Finding|Idea or Concept|History of Present Illness|570,577|false|true|false|C1550516|Target Awareness - partial|partial
Event|Event|History of Present Illness|578,586|false|false|false|||thrombus
Finding|Pathologic Function|History of Present Illness|578,586|false|true|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Event|Event|History of Present Illness|590,598|false|false|false|||stenosis
Finding|Pathologic Function|History of Present Illness|590,598|false|false|false|C1261287|Stenosis|stenosis
Event|Activity|History of Present Illness|612,620|false|false|false|C2919031|Division (action)|division
Event|Event|History of Present Illness|612,620|false|false|false|||division
Finding|Idea or Concept|History of Present Illness|612,620|false|false|false|C1547541|Organization Unit Type - Division|division
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|612,620|false|false|false|C0152060;C1293097|Division (surgical procedure);Transection (procedure)|division
Event|Event|History of Present Illness|631,642|false|false|false|||Transferred
Event|Activity|History of Present Illness|660,670|false|false|false|C1283169||monitoring
Event|Event|History of Present Illness|660,670|false|false|false|||monitoring
Procedure|Health Care Activity|History of Present Illness|660,670|false|false|false|C0150369|Preventive monitoring|monitoring
Finding|Finding|History of Present Illness|675,683|false|false|false|C0332149|Possible|possible
Event|Event|History of Present Illness|684,696|false|false|false|||thrombectomy
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|684,696|false|false|false|C0162578|Thrombectomy|thrombectomy
Event|Event|History of Present Illness|704,708|false|false|false|||exam
Finding|Functional Concept|History of Present Illness|704,708|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|History of Present Illness|704,708|false|false|false|C0582103|Medical Examination|exam
Event|Event|History of Present Illness|718,725|false|false|false|||worsens
Event|Event|History of Present Illness|728,735|false|false|false|||History
Finding|Conceptual Entity|History of Present Illness|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Finding|History of Present Illness|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Finding|Functional Concept|History of Present Illness|728,735|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|History
Event|Event|History of Present Illness|736,744|false|false|false|||obtained
Finding|Body Substance|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|750,757|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Body Substance|History of Present Illness|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|History of Present Illness|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|History of Present Illness|783,790|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|History of Present Illness|808,817|false|false|false|||historian
Event|Event|History of Present Illness|837,843|false|false|false|||dinner
Finding|Daily or Recreational Activity|History of Present Illness|837,843|false|false|false|C4048877|Dinner|dinner
Event|Event|History of Present Illness|849,856|false|false|false|||friends
Finding|Intellectual Product|History of Present Illness|861,865|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|History of Present Illness|866,874|false|false|false|||returned
Event|Event|History of Present Illness|883,892|false|false|false|||apartment
Event|Event|History of Present Illness|901,908|false|false|false|||fooling
Finding|Finding|History of Present Illness|945,949|false|false|false|C5575035|Well (answer to question)|well
Finding|Intellectual Product|History of Present Illness|971,975|false|false|false|C1720594|Then - dosing instruction fragment|Then
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|988,991|false|false|false|C0029121|Oppositional Defiant Disorder|odd
Finding|Gene or Genome|History of Present Illness|988,991|false|false|false|C1415068;C1418191|GJA1 gene;OSR1 gene|odd
Event|Event|History of Present Illness|992,1001|false|false|false|||sensation
Finding|Finding|History of Present Illness|992,1001|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|History of Present Illness|992,1001|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|History of Present Illness|992,1001|false|false|false|C2229507|sensory exam|sensation
Event|Event|History of Present Illness|1006,1013|false|false|false|||started
Event|Event|History of Present Illness|1015,1023|false|false|false|||throwing
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1028,1032|false|false|false|C0446516|Upper arm|arms
Attribute|Clinical Attribute|History of Present Illness|1028,1032|false|false|false|C5782111||arms
Disorder|Neoplastic Process|History of Present Illness|1028,1032|false|false|false|C0206655|Alveolar rhabdomyosarcoma|arms
Event|Event|History of Present Illness|1028,1032|false|false|false|||arms
Finding|Gene or Genome|History of Present Illness|1028,1032|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Finding|Intellectual Product|History of Present Illness|1028,1032|false|false|false|C2681631;C5575339|Adherence to Refills and Medications Scale;KIDINS220 gene|arms
Event|Event|History of Present Illness|1068,1071|false|false|false|||sit
Event|Event|History of Present Illness|1082,1087|false|false|false|||tried
Event|Event|History of Present Illness|1091,1095|false|false|false|||read
Event|Event|History of Present Illness|1110,1113|false|false|false|||see
Finding|Intellectual Product|History of Present Illness|1138,1142|false|false|false|C1720594|Then - dosing instruction fragment|Then
Finding|Classification|History of Present Illness|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|1149,1155|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|History of Present Illness|1169,1177|false|false|false|||knocking
Event|Event|History of Present Illness|1204,1209|false|false|false|||tough
Finding|Finding|History of Present Illness|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|1211,1215|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|History of Present Illness|1216,1224|false|false|false|||standing
Event|Event|History of Present Illness|1250,1254|false|false|false|||able
Finding|Finding|History of Present Illness|1250,1254|false|false|false|C1299581|Able (qualifier value)|able
Finding|Gene or Genome|History of Present Illness|1284,1289|false|false|false|C1424898|RXFP2 gene|great
Event|Event|History of Present Illness|1290,1300|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1290,1300|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|1305,1311|false|false|false|||walked
Finding|Finding|History of Present Illness|1333,1340|false|false|false|C3888388|Usually|usually
Event|Event|History of Present Illness|1342,1347|false|false|false|||walks
Event|Event|History of Present Illness|1355,1361|false|false|false|||walker
Anatomy|Body Location or Region|History of Present Illness|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|History of Present Illness|1373,1377|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|History of Present Illness|1373,1377|false|false|false|C0562271|Examination of knee joint|knee
Attribute|Clinical Attribute|History of Present Illness|1373,1389|false|false|false|C5575606||knee replacement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1373,1389|false|false|false|C0086511|Knee Replacement Arthroplasty|knee replacement
Event|Event|History of Present Illness|1378,1389|false|false|false|||replacement
Finding|Functional Concept|History of Present Illness|1378,1389|false|false|false|C0559956|Replacement|replacement
Procedure|Health Care Activity|History of Present Illness|1378,1389|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1378,1389|false|false|false|C0035139;C1555302|Replacement - supply;Surgical Replantation|replacement
Event|Event|History of Present Illness|1404,1406|false|false|false|||up
Event|Event|History of Present Illness|1437,1443|false|false|false|||walked
Event|Event|History of Present Illness|1459,1465|false|false|false|||unlock
Finding|Idea or Concept|History of Present Illness|1459,1465|false|false|false|C1550031|Unlock|unlock
Event|Event|History of Present Illness|1480,1488|false|false|false|||problems
Finding|Idea or Concept|History of Present Illness|1480,1488|false|false|false|C1546466|Problems - What subject filter|problems
Event|Event|History of Present Illness|1489,1496|false|false|false|||talking
Finding|Classification|History of Present Illness|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|1500,1506|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|History of Present Illness|1524,1534|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1524,1534|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|1544,1549|false|false|false|||words
Event|Event|History of Present Illness|1566,1571|false|false|false|||words
Event|Event|History of Present Illness|1573,1579|false|false|false|||Denies
Finding|Idea or Concept|History of Present Illness|1580,1584|false|false|false|C1705313|Term (lexical)|word
Event|Event|History of Present Illness|1585,1592|false|false|false|||finding
Finding|Finding|History of Present Illness|1585,1592|true|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|History of Present Illness|1585,1592|true|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Event|Event|History of Present Illness|1594,1604|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1594,1604|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Event|Event|History of Present Illness|1616,1620|false|false|false|||tell
Event|Event|History of Present Illness|1628,1635|false|false|false|||slurred
Attribute|Clinical Attribute|History of Present Illness|1643,1649|false|false|true|C5890614||person
Finding|Intellectual Product|History of Present Illness|1643,1649|false|false|true|C1522390|Person Info|person
Finding|Finding|History of Present Illness|1659,1667|false|false|false|C3843660|Too much|too much
Event|Event|History of Present Illness|1663,1667|false|false|false|||much
Finding|Finding|History of Present Illness|1663,1667|false|false|false|C4281574|Much|much
Event|Event|History of Present Illness|1671,1676|false|false|false|||drink
Event|Event|History of Present Illness|1683,1688|false|false|false|||asked
Event|Event|History of Present Illness|1700,1711|false|false|false|||intoxicated
Event|Event|History of Present Illness|1743,1748|false|false|false|||aware
Finding|Mental Process|History of Present Illness|1743,1748|false|false|false|C0004448|Awareness|aware
Disorder|Mental or Behavioral Dysfunction|History of Present Illness|1756,1766|false|false|false|C0013362|Dysarthria|dysarthria
Event|Event|History of Present Illness|1756,1766|false|false|false|||dysarthria
Event|Event|History of Present Illness|1771,1775|false|false|false|||told
Event|Event|History of Present Illness|1780,1789|false|false|false|||daughters
Event|Event|History of Present Illness|1800,1806|false|false|false|||thinks
Event|Event|History of Present Illness|1810,1812|false|false|false|||'s
Disorder|Disease or Syndrome|History of Present Illness|1822,1828|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|History of Present Illness|1822,1828|false|false|false|||stroke
Finding|Finding|History of Present Illness|1822,1828|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|History of Present Illness|1830,1834|false|false|false|C1720594|Then - dosing instruction fragment|Then
Event|Event|History of Present Illness|1840,1844|false|false|false|||said
Event|Event|History of Present Illness|1862,1869|false|false|false|||sitting
Event|Event|History of Present Illness|1886,1890|false|false|false|||idea
Event|Event|History of Present Illness|1899,1906|false|false|false|||thought
Event|Event|History of Present Illness|1945,1949|false|false|false|||able
Finding|Finding|History of Present Illness|1945,1949|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|1953,1957|false|false|false|||walk
Event|Event|History of Present Illness|1963,1969|false|false|false|||walker
Event|Event|History of Present Illness|1978,1982|false|false|false|||felt
Event|Event|History of Present Illness|2004,2008|false|false|false|||fell
Finding|Functional Concept|History of Present Illness|2013,2019|false|false|false|C0234621|Visual|visual
Finding|Finding|History of Present Illness|2013,2027|true|false|false|C0750280|Visual changes|visual changes
Event|Event|History of Present Illness|2020,2027|false|false|false|||changes
Finding|Functional Concept|History of Present Illness|2020,2027|true|false|false|C0392747|Changing|changes
Event|Event|History of Present Illness|2032,2040|false|false|false|||numbness
Finding|Finding|History of Present Illness|2032,2040|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|2032,2040|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|History of Present Illness|2045,2053|false|false|false|C0030554|Paresthesia|tingling
Event|Event|History of Present Illness|2045,2053|false|false|false|||tingling
Finding|Sign or Symptom|History of Present Illness|2045,2053|false|false|false|C2242996|Has tingling sensation|tingling
Event|Event|History of Present Illness|2055,2061|false|false|false|||Denies
Event|Event|History of Present Illness|2068,2076|false|false|false|||weakness
Finding|Sign or Symptom|History of Present Illness|2068,2076|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Event|Event|History of Present Illness|2091,2098|false|false|false|||trouble
Event|Event|History of Present Illness|2121,2125|false|false|false|||able
Finding|Finding|History of Present Illness|2121,2125|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|History of Present Illness|2129,2135|false|false|false|||unlock
Event|Event|History of Present Illness|2140,2144|false|false|false|||door
Event|Activity|History of Present Illness|2153,2158|true|false|false|C5966184|Issue (action)|issue
Event|Event|History of Present Illness|2153,2158|false|false|false|||issue
Finding|Finding|History of Present Illness|2153,2158|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Finding|Intellectual Product|History of Present Illness|2153,2158|true|false|false|C0033213;C1706387|Issue (document);Problem|issue
Event|Event|History of Present Illness|2167,2171|false|false|false|||felt
Event|Event|History of Present Illness|2173,2178|false|false|false|||shaky
Finding|Finding|History of Present Illness|2173,2178|false|false|false|C0392703|Shakes|shaky
Event|Event|History of Present Illness|2190,2197|false|false|false|||brought
Drug|Hazardous or Poisonous Substance|History of Present Illness|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|History of Present Illness|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|History of Present Illness|2201,2204|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Event|Event|History of Present Illness|2201,2204|false|false|false|||EMS
Finding|Gene or Genome|History of Present Illness|2201,2204|false|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|History of Present Illness|2201,2204|false|false|false|C0013961|Emergency Medical Services|EMS
Event|Event|History of Present Illness|2218,2223|false|false|false|||NIHSS
Finding|Intellectual Product|History of Present Illness|2218,2223|false|false|false|C1697238|NIH stroke scale|NIHSS
Event|Event|History of Present Illness|2235,2242|false|false|false|||slurred
Event|Event|History of Present Illness|2243,2249|false|false|false|||speech
Finding|Organism Function|History of Present Illness|2243,2249|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|History of Present Illness|2243,2249|false|false|false|C0846595|Speech assessment|speech
Event|Event|History of Present Illness|2262,2266|false|false|false|||felt
Event|Event|History of Present Illness|2284,2292|false|false|false|||symptoms
Finding|Functional Concept|History of Present Illness|2284,2292|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|History of Present Illness|2284,2292|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|History of Present Illness|2294,2301|false|false|false|||started
Event|Event|History of Present Illness|2305,2312|false|false|false|||improve
Event|Event|History of Present Illness|2322,2329|false|false|false|||started
Event|Event|History of Present Illness|2336,2347|false|false|false|||transferred
Event|Event|History of Present Illness|2361,2365|false|false|false|||said
Event|Event|History of Present Illness|2370,2376|false|false|false|||speech
Finding|Organism Function|History of Present Illness|2370,2376|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|History of Present Illness|2370,2376|false|false|false|C0846595|Speech assessment|speech
Event|Event|History of Present Illness|2381,2390|false|false|false|||improving
Finding|Idea or Concept|History of Present Illness|2417,2422|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Finding|Intellectual Product|History of Present Illness|2417,2422|false|false|false|C1561541;C1561542|Precision - month;Transaction counts and value totals - month|month
Event|Event|History of Present Illness|2424,2431|false|false|false|||started
Drug|Organic Chemical|History of Present Illness|2440,2444|false|false|false|C0067518|N-(4-aminophenethyl)spiroperidol|naps
Event|Event|History of Present Illness|2440,2444|false|false|false|||naps
Event|Event|History of Present Illness|2450,2457|false|false|false|||hearing
Finding|Finding|History of Present Illness|2450,2457|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|History of Present Illness|2450,2457|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Event|Event|History of Present Illness|2461,2465|false|false|false|||poor
Finding|Intellectual Product|History of Present Illness|2461,2465|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Drug|Biomedical or Dental Material|History of Present Illness|2470,2478|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|2470,2478|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|2470,2478|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|History of Present Illness|2501,2508|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|History of Present Illness|2501,2508|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|History of Present Illness|2509,2513|false|false|false|C0001175|Acquired Immunodeficiency Syndrome|aids
Event|Event|History of Present Illness|2509,2513|false|false|false|||aids
Event|Event|History of Present Illness|2567,2574|false|false|false|||nightly
Event|Event|History of Present Illness|2580,2587|false|false|false|||dysuria
Finding|Sign or Symptom|History of Present Illness|2580,2587|false|false|false|C0013428|Dysuria|dysuria
Event|Event|History of Present Illness|2599,2606|false|false|false|||noticed
Finding|Sign or Symptom|History of Present Illness|2612,2630|false|false|false|C0948396|Frequent headache|frequent headaches
Event|Event|History of Present Illness|2621,2630|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|2621,2630|false|false|false|C0018681|Headache|headaches
Event|Event|History of Present Illness|2668,2676|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2668,2676|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|2681,2690|false|false|false|||yesterday
Drug|Organic Chemical|History of Present Illness|2702,2710|false|false|false|C0040610|tramadol|tramadol
Drug|Pharmacologic Substance|History of Present Illness|2702,2710|false|false|false|C0040610|tramadol|tramadol
Event|Event|History of Present Illness|2702,2710|false|false|false|||tramadol
Procedure|Laboratory Procedure|History of Present Illness|2702,2710|false|false|false|C1266765|Tramadol measurement (procedure)|tramadol
Drug|Organic Chemical|History of Present Illness|2716,2729|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Drug|Pharmacologic Substance|History of Present Illness|2716,2729|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|acetaminophen
Event|Event|History of Present Illness|2716,2729|false|false|false|||acetaminophen
Procedure|Laboratory Procedure|History of Present Illness|2716,2729|false|false|false|C0373527|Acetaminophen measurement|acetaminophen
Event|Event|History of Present Illness|2738,2744|false|false|false|||couple
Finding|Functional Concept|History of Present Illness|2738,2744|false|false|false|C1948027|Couple (action)|couple
Event|Event|History of Present Illness|2764,2771|false|false|false|||reports
Event|Event|History of Present Illness|2773,2782|false|false|false|||headaches
Finding|Sign or Symptom|History of Present Illness|2773,2782|false|false|false|C0018681|Headache|headaches
Event|Event|History of Present Illness|2798,2802|false|false|false|||wake
Event|Event|History of Present Illness|2815,2821|false|false|false|||denies
Event|Event|History of Present Illness|2832,2840|false|false|false|||headache
Finding|Sign or Symptom|History of Present Illness|2832,2840|false|false|false|C0018681|Headache|headache
Event|Event|History of Present Illness|2844,2854|false|false|false|||positional
Finding|Finding|History of Present Illness|2844,2854|false|false|false|C0240795|positional|positional
Event|Event|History of Present Illness|2871,2878|false|false|false|||sitting
Event|Event|History of Present Illness|2885,2890|false|false|false|||lying
Attribute|Clinical Attribute|History of Present Illness|2923,2929|false|false|false|C0944911||weight
Event|Event|History of Present Illness|2923,2929|false|false|false|||weight
Finding|Finding|History of Present Illness|2923,2929|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|History of Present Illness|2923,2929|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|History of Present Illness|2923,2929|false|false|false|C1305866|Weighing patient|weight
Finding|Finding|History of Present Illness|2923,2934|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Finding|Intellectual Product|History of Present Illness|2923,2934|false|false|false|C1262477;C3540682|Losing Weight (question);Weight Loss|weight loss
Event|Event|History of Present Illness|2930,2934|false|false|false|||loss
Finding|Finding|History of Present Illness|2930,2934|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Idea or Concept|History of Present Illness|2965,2969|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|History of Present Illness|2965,2969|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Gene or Genome|History of Present Illness|2970,2973|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|History of Present Illness|2994,2997|false|false|false|||lbs
Procedure|Laboratory Procedure|History of Present Illness|2994,2997|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|History of Present Illness|3018,3021|false|false|false|||lbs
Procedure|Laboratory Procedure|History of Present Illness|3018,3021|false|false|false|C3161851|liquid-based cytology (procedure)|lbs
Event|Event|History of Present Illness|3027,3035|false|false|false|||appetite
Finding|Organism Function|History of Present Illness|3027,3035|false|false|false|C0003618|Desire for food|appetite
Disorder|Disease or Syndrome|History of Present Illness|3040,3045|false|false|false|C1410088|Still|still
Event|Event|History of Present Illness|3046,3050|false|false|false|||good
Finding|Idea or Concept|History of Present Illness|3046,3050|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|History of Present Illness|3059,3065|false|false|false|||enjoys
Event|Event|History of Present Illness|3066,3072|false|false|false|||eating
Event|Event|History of Present Illness|3089,3095|false|false|false|||hungry
Finding|Sign or Symptom|History of Present Illness|3089,3095|false|false|false|C0020175|Hunger|hungry
Event|Event|History of Present Illness|3106,3110|false|false|false|||used
Event|Event|History of Present Illness|3130,3134|false|false|false|||says
Event|Event|History of Present Illness|3159,3166|false|false|false|||decline
Event|Event|History of Present Illness|3170,3176|false|false|false|||memory
Finding|Finding|History of Present Illness|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|History of Present Illness|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|3170,3176|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Event|Event|History of Present Illness|3242,3247|false|false|false|||plans
Disorder|Disease or Syndrome|History of Present Illness|3250,3255|false|false|false|C5975557|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|times
Event|Event|History of Present Illness|3250,3255|false|false|false|||times
Event|Event|History of Present Illness|3260,3267|false|false|false|||pickpup
Finding|Daily or Recreational Activity|History of Present Illness|3273,3279|false|false|false|C4048877|Dinner|dinner
Event|Event|History of Present Illness|3280,3285|false|false|false|||plans
Event|Event|History of Present Illness|3297,3303|false|false|false|||become
Event|Event|History of Present Illness|3304,3310|false|false|false|||normal
Finding|Classification|History of Present Illness|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|History of Present Illness|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|History of Present Illness|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|History of Present Illness|3338,3344|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Event|Event|History of Present Illness|3349,3356|false|false|false|||noticed
Event|Event|History of Present Illness|3366,3375|false|false|false|||worsening
Event|Event|History of Present Illness|3390,3398|false|false|false|||remember
Event|Event|History of Present Illness|3405,3414|false|false|false|||grandkids
Event|Event|History of Present Illness|3420,3426|false|false|false|||coming
Event|Event|History of Present Illness|3430,3435|false|false|false|||visit
Finding|Social Behavior|History of Present Illness|3430,3435|false|false|false|C0545082|Visit|visit
Event|Event|History of Present Illness|3446,3452|false|false|false|||bought
Finding|Gene or Genome|History of Present Illness|3457,3462|false|false|false|C4321205|MELTF-AS1 gene|plane
Event|Event|History of Present Illness|3463,3470|false|false|false|||tickets
Event|Event|History of Present Illness|3485,3493|false|false|false|||endorses
Event|Event|History of Present Illness|3503,3512|false|false|false|||orthopnea
Finding|Finding|History of Present Illness|3503,3512|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Finding|Sign or Symptom|History of Present Illness|3503,3512|false|false|false|C0085619;C2188830|Orthopnea;sleeping upright or using specific number of extra pillows (orthopnea)|orthopnea
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|3554,3560|false|false|false|C0018792|Heart Atrium|Atrial
Attribute|Clinical Attribute|Past Medical History|3554,3573|false|false|false|C2926591||Atrial fibrillation
Disorder|Disease or Syndrome|Past Medical History|3554,3573|false|false|false|C0004238|Atrial Fibrillation|Atrial fibrillation
Lab|Laboratory or Test Result|Past Medical History|3554,3573|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Atrial fibrillation
Disorder|Disease or Syndrome|Past Medical History|3561,3573|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Past Medical History|3561,3573|false|false|false|||fibrillation
Drug|Organic Chemical|Past Medical History|3577,3584|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|Past Medical History|3577,3584|false|false|false|C3530466|Eliquis|Eliquis
Event|Event|Past Medical History|3577,3584|false|false|false|||Eliquis
Anatomy|Body Space or Junction|Past Medical History|3585,3588|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Past Medical History|3585,3588|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Past Medical History|3585,3588|false|false|false|||CHF
Disorder|Disease or Syndrome|Past Medical History|3589,3609|false|false|false|C0020443|Hypercholesterolemia|Hypercholesterolemia
Event|Event|Past Medical History|3589,3609|false|false|false|||Hypercholesterolemia
Finding|Finding|Past Medical History|3589,3609|false|false|false|C1522133|Hypercholesterolemia result|Hypercholesterolemia
Disorder|Disease or Syndrome|Past Medical History|3610,3622|false|false|false|C0020538|Hypertensive disease|Hypertension
Event|Event|Past Medical History|3610,3622|false|false|false|||Hypertension
Finding|Conceptual Entity|Family Medical History|3661,3667|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|3661,3667|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Finding|Family Medical History|3670,3676|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Family Medical History|3670,3676|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Event|Event|Family Medical History|3677,3686|false|false|false|||alcoholic
Disorder|Mental or Behavioral Dysfunction|Family Medical History|3688,3701|false|false|false|C0036341|Schizophrenia|schizophrenia
Event|Event|Family Medical History|3688,3701|false|false|false|||schizophrenia
Finding|Idea or Concept|Family Medical History|3702,3708|false|false|false|C1546508|Relationship - Mother|Mother
Anatomy|Body Space or Junction|Family Medical History|3711,3714|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Family Medical History|3711,3714|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Family Medical History|3711,3714|false|false|false|||CHF
Finding|Conceptual Entity|Family Medical History|3715,3722|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Finding|Idea or Concept|Family Medical History|3715,3722|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|Brother
Disorder|Disease or Syndrome|Family Medical History|3725,3731|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Family Medical History|3725,3731|false|false|false|||stroke
Finding|Finding|Family Medical History|3725,3731|false|false|false|C5977286|Stroke (heart beat)|stroke
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|3733,3740|false|false|false|C0007272|Carotid Arteries|carotid
Disorder|Disease or Syndrome|Family Medical History|3733,3749|false|false|false|C0007282|Carotid Stenosis|carotid stenosis
Event|Event|Family Medical History|3741,3749|false|false|false|||stenosis
Finding|Pathologic Function|Family Medical History|3741,3749|false|false|false|C1261287|Stenosis|stenosis
Procedure|Health Care Activity|General Exam|3767,3776|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3777,3781|false|false|false|||EXAM
Finding|Functional Concept|General Exam|3777,3781|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3777,3781|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3849,3856|false|false|false|||General
Finding|Classification|General Exam|3849,3856|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3849,3856|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|3858,3863|false|false|false|||Awake
Finding|Finding|General Exam|3858,3863|false|false|false|C0234422|Awake (finding)|Awake
Disorder|Disease or Syndrome|General Exam|3892,3895|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|3892,3895|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|3892,3895|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|3892,3895|false|false|false|||NAD
Finding|Finding|General Exam|3892,3895|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|3897,3902|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3914,3921|false|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|3914,3929|true|false|false|C0240962|Scleral icterus|scleral icterus
Event|Event|General Exam|3922,3929|false|false|false|||icterus
Finding|Sign or Symptom|General Exam|3922,3929|true|false|false|C0022346|Icterus|icterus
Event|Event|General Exam|3930,3935|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|3937,3940|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3937,3940|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|3945,3952|false|false|false|||lesions
Finding|Finding|General Exam|3945,3952|true|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|3953,3958|false|false|false|||noted
Anatomy|Body Location or Region|General Exam|3962,3972|false|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Location or Region|General Exam|3974,3978|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3974,3978|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3974,3978|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|3980,3986|false|false|false|||Supple
Finding|Functional Concept|General Exam|3980,3986|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|3991,4006|true|false|false|C1320474|Nuchal Rigidity|nuchal rigidity
Event|Event|General Exam|3998,4006|false|false|false|||rigidity
Finding|Sign or Symptom|General Exam|3998,4006|true|false|false|C0026837|Muscle Rigidity|rigidity
Phenomenon|Natural Phenomenon or Process|General Exam|3998,4006|true|false|false|C0700109|plastic property - rigidity|rigidity
Anatomy|Body Part, Organ, or Organ Component|General Exam|4008,4017|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|General Exam|4008,4017|false|false|false|C2707265||Pulmonary
Finding|Finding|General Exam|4008,4017|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|General Exam|4026,4030|false|false|false|||work
Event|Occupational Activity|General Exam|4026,4030|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|4026,4043|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|4034,4043|false|false|false|C5885990||breathing
Event|Event|General Exam|4034,4043|false|false|false|||breathing
Finding|Finding|General Exam|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|4034,4043|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|4034,4043|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Part, Organ, or Organ Component|General Exam|4045,4052|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|General Exam|4045,4052|false|false|false|C1314974|Cardiac attachment|Cardiac
Event|Event|General Exam|4054,4057|false|false|false|||RRR
Event|Event|General Exam|4059,4063|false|false|false|||warm
Finding|Finding|General Exam|4059,4063|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|4059,4063|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|4065,4069|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|4070,4078|false|false|false|||perfused
Anatomy|Body Location or Region|General Exam|4080,4087|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|4080,4087|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|4080,4087|false|false|false|||Abdomen
Finding|Finding|General Exam|4080,4087|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|4089,4093|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|4089,4093|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|4110,4121|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|General Exam|4130,4135|false|false|false|C1717255||edema
Event|Event|General Exam|4130,4135|false|false|false|||edema
Finding|Pathologic Function|General Exam|4130,4135|false|false|false|C0013604|Edema|edema
Anatomy|Body System|General Exam|4137,4141|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|4137,4141|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|4137,4141|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|4137,4141|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|4137,4141|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|4143,4153|false|false|false|||ecchymoses
Finding|Pathologic Function|General Exam|4143,4153|false|false|false|C0013491|Ecchymosis|ecchymoses
Anatomy|Body Location or Region|General Exam|4159,4163|false|false|false|C0230444|Shin|shin
Event|Event|General Exam|4170,4179|false|false|false|||extensive
Anatomy|Body Location or Region|General Exam|4185,4189|false|false|false|C0230444|Shin|shin
Finding|Mental Process|General Exam|4207,4213|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|4207,4220|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|General Exam|4207,4220|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|General Exam|4214,4220|false|false|false|C5889824||Status
Event|Event|General Exam|4214,4220|false|false|false|||Status
Finding|Idea or Concept|General Exam|4214,4220|false|false|false|C1546481|What subject filter - Status|Status
Attribute|Clinical Attribute|General Exam|4222,4227|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|4222,4227|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|4222,4227|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|4222,4227|false|false|false|||Alert
Finding|Finding|General Exam|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|4222,4227|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|4229,4237|false|false|false|||oriented
Finding|Finding|General Exam|4243,4247|false|false|false|C1299581|Able (qualifier value)|Able
Event|Event|General Exam|4258,4265|false|false|false|||history
Finding|Conceptual Entity|General Exam|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|4258,4265|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|General Exam|4297,4301|false|false|false|||able
Finding|Finding|General Exam|4297,4301|false|false|false|C1299581|Able (qualifier value)|able
Finding|Intellectual Product|General Exam|4305,4309|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Attribute|Clinical Attribute|General Exam|4343,4351|true|false|false|C2706915||Language
Event|Event|General Exam|4343,4351|false|false|false|||Language
Finding|Intellectual Product|General Exam|4343,4351|true|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|4355,4361|false|false|false|||fluent
Finding|Finding|General Exam|4367,4373|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|4374,4384|false|false|false|||repetition
Finding|Finding|General Exam|4374,4384|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Finding|Functional Concept|General Exam|4374,4384|false|false|false|C0205341;C2018025|Repeat;speech fluency repetition (physical finding)|repetition
Event|Event|General Exam|4389,4402|false|false|false|||comprehension
Finding|Mental Process|General Exam|4389,4402|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|4411,4418|false|false|false|||prosody
Finding|Finding|General Exam|4411,4418|false|false|false|C0233743|Prosody|prosody
Event|Event|General Exam|4445,4451|false|false|false|||errors
Finding|Finding|General Exam|4453,4457|false|false|false|C1299581|Able (qualifier value)|Able
Finding|Intellectual Product|General Exam|4461,4465|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|name
Finding|Finding|General Exam|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|General Exam|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|General Exam|4471,4475|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|General Exam|4480,4483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|4480,4483|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|General Exam|4484,4493|false|false|false|||frequency
Finding|Intellectual Product|General Exam|4484,4493|false|false|false|C3898838;C4321352|Frequency;How Often|frequency
Event|Event|General Exam|4494,4501|false|false|false|||objects
Finding|Finding|General Exam|4504,4508|false|false|false|C1299581|Able (qualifier value)|Able
Event|Event|General Exam|4512,4516|false|false|false|||read
Event|Event|General Exam|4525,4535|false|false|false|||difficulty
Finding|Finding|General Exam|4525,4535|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Disorder|Mental or Behavioral Dysfunction|General Exam|4540,4550|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|4540,4550|false|false|false|||dysarthria
Finding|Finding|General Exam|4552,4556|false|false|false|C1299581|Able (qualifier value)|Able
Event|Event|General Exam|4561,4567|false|false|false|||follow
Anatomy|Cell Component|General Exam|4573,4580|false|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|4598,4606|false|false|false|||commands
Event|Event|General Exam|4621,4629|false|false|false|||evidence
Finding|Idea or Concept|General Exam|4621,4629|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|4621,4632|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|General Exam|4633,4640|true|false|false|C0003635|Apraxias|apraxia
Event|Event|General Exam|4633,4640|false|false|false|||apraxia
Event|Event|General Exam|4644,4651|false|false|false|||neglect
Event|Event|General Exam|4644,4651|false|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|General Exam|4644,4651|false|false|false|C0521874|Victim of neglect (finding)|neglect
Anatomy|Body Part, Organ, or Organ Component|General Exam|4655,4662|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4655,4669|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|4655,4669|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|4663,4669|false|false|false|C0027740|Nerve|Nerves
Finding|Finding|General Exam|4689,4694|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|4715,4719|false|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|4728,4737|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|4728,4737|false|false|false|||nystagmus
Event|Event|General Exam|4746,4754|false|false|false|||saccades
Finding|Finding|General Exam|4746,4754|false|false|false|C0036019|Saccades|saccades
Event|Event|General Exam|4756,4759|false|false|false|||VFF
Event|Event|General Exam|4763,4776|false|false|false|||confrontation
Finding|Finding|General Exam|4763,4776|false|false|false|C0518608|Social confrontation skill|confrontation
Procedure|Diagnostic Procedure|General Exam|4763,4776|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Procedure|Therapeutic or Preventive Procedure|General Exam|4763,4776|false|false|false|C0700282;C1444674|Confrontation;Confrontation visual field test|confrontation
Anatomy|Body Location or Region|General Exam|4782,4788|false|false|false|C0015450|Face|Facial
Finding|Finding|General Exam|4782,4798|false|false|false|C0517999|facial sensation|Facial sensation
Event|Event|General Exam|4789,4798|false|false|false|||sensation
Finding|Finding|General Exam|4789,4798|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|4789,4798|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|4789,4798|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|4799,4805|false|false|false|||intact
Finding|Finding|General Exam|4799,4805|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|General Exam|4809,4814|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|4809,4814|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|4809,4814|false|false|false|||light
Finding|Finding|General Exam|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|4809,4814|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|4809,4814|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|4809,4814|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|4809,4820|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|4815,4820|false|false|false|||touch
Finding|Mental Process|General Exam|4815,4820|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|4815,4820|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|4815,4820|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|4825,4833|false|false|false|||pinprick
Anatomy|Body Part, Organ, or Organ Component|General Exam|4835,4838|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|4835,4838|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|4843,4849|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|General Exam|4843,4855|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|General Exam|4843,4855|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|General Exam|4850,4855|false|false|false|||droop
Anatomy|Body Location or Region|General Exam|4857,4863|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4864,4875|false|false|false|C1995013|Set of muscles|musculature
Event|Event|General Exam|4876,4885|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|4876,4885|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|4876,4885|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|4887,4891|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|4887,4891|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|4887,4891|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|General Exam|4893,4900|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|4893,4900|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|4901,4907|false|false|false|||intact
Finding|Finding|General Exam|4901,4907|false|false|false|C1554187|Gender Status - Intact|intact
Anatomy|Body Part, Organ, or Organ Component|General Exam|4911,4917|false|false|false|C0016129;C0851278;C4299059|Fingers;Fingers not including thumb;Upper extremity>Finger|finger
Drug|Biomedical or Dental Material|General Exam|4918,4926|false|false|false|C1177045|Snap brand of resin|snapping
Event|Event|General Exam|4918,4926|false|false|false|||snapping
Event|Event|General Exam|4940,4945|false|false|false|||bring
Finding|Finding|General Exam|4950,4957|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Finding|Physiologic Function|General Exam|4950,4957|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|hearing
Disorder|Disease or Syndrome|General Exam|4958,4962|false|false|false|C0001175|Acquired Immunodeficiency Syndrome|aids
Event|Event|General Exam|4958,4962|false|false|false|||aids
Anatomy|Body Part, Organ, or Organ Component|General Exam|4972,4978|false|false|false|C0700374|Palate|Palate
Event|Event|General Exam|4979,4987|false|false|false|||elevates
Event|Event|General Exam|5011,5019|false|false|false|||strength
Finding|Idea or Concept|General Exam|5011,5019|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|5050,5056|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|5050,5056|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Event|Event|General Exam|5050,5056|false|false|false|||Tongue
Procedure|Health Care Activity|General Exam|5050,5056|false|false|false|C0872394|Procedure on tongue|Tongue
Event|Event|General Exam|5057,5066|false|false|false|||protrudes
Anatomy|Cell Component|General Exam|5070,5077|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|General Exam|5083,5087|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|5088,5098|false|false|false|||excursions
Finding|Idea or Concept|General Exam|5100,5108|false|false|false|C0808080|Strength (attribute)|Strength
Event|Event|General Exam|5109,5113|false|false|false|||full
Anatomy|Body Part, Organ, or Organ Component|General Exam|5119,5125|false|false|false|C0040408|Tongue|tongue
Disorder|Neoplastic Process|General Exam|5119,5125|false|false|false|C0153933|Benign neoplasm of tongue|tongue
Event|Event|General Exam|5119,5125|false|false|false|||tongue
Procedure|Health Care Activity|General Exam|5119,5125|false|false|false|C0872394|Procedure on tongue|tongue
Anatomy|Body Location or Region|General Exam|5129,5134|false|false|false|C0007966|Cheek structure|cheek
Event|Event|General Exam|5135,5142|false|false|false|||testing
Finding|Functional Concept|General Exam|5135,5142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Intellectual Product|General Exam|5135,5142|false|false|false|C0039593;C0392366|Testing;Tests (qualifier value)|testing
Finding|Functional Concept|General Exam|5146,5151|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|5160,5164|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|5160,5164|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|5169,5173|false|false|false|||tone
Finding|Pathologic Function|General Exam|5189,5203|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|5198,5203|false|false|false|||drift
Event|Event|General Exam|5221,5230|false|false|false|||movements
Finding|Organism Function|General Exam|5221,5230|false|false|false|C0026649|Movement|movements
Event|Event|General Exam|5240,5246|false|false|false|||tremor
Finding|Sign or Symptom|General Exam|5240,5246|false|false|false|C0040822|Tremor|tremor
Event|Event|General Exam|5250,5259|false|false|false|||asterixis
Finding|Sign or Symptom|General Exam|5250,5259|false|false|false|C0232766|Asterixis|asterixis
Event|Event|General Exam|5260,5265|false|false|false|||noted
Event|Event|General Exam|5409,5417|false|false|false|||deficits
Drug|Amino Acid, Peptide, or Protein|General Exam|5421,5426|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|5421,5426|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|5421,5426|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|5421,5426|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|5421,5426|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|5421,5432|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|5427,5432|false|false|false|||touch
Finding|Mental Process|General Exam|5427,5432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|5427,5432|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|5427,5432|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|5434,5442|false|false|false|||pinprick
Event|Event|General Exam|5444,5455|false|false|false|||temperature
Procedure|Health Care Activity|General Exam|5444,5455|false|false|false|C0886414|Body temperature measurement|temperature
Finding|Finding|General Exam|5468,5477|false|false|false|C0392756;C0442797|Decreasing;Reduced|Decreased
Finding|Finding|General Exam|5468,5493|false|false|false|C1295585|Decreased vibratory sense|Decreased vibratory sense
Finding|Organism Function|General Exam|5478,5493|false|false|false|C0234198||vibratory sense
Event|Event|General Exam|5488,5493|false|false|false|||sense
Finding|Organ or Tissue Function|General Exam|5488,5493|false|false|false|C0036658|Sensory perception|sense
Anatomy|Body Part, Organ, or Organ Component|General Exam|5501,5505|false|false|false|C0016504|Foot|feet
Anatomy|Body Location or Region|General Exam|5512,5518|false|false|false|C0003086|Ankle|ankles
Anatomy|Body Space or Junction|General Exam|5520,5525|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Anatomy|Body System|General Exam|5520,5525|false|false|false|C0022417;C0392905;C1269611|Articular system;Joints|Joint
Finding|Finding|General Exam|5520,5525|false|false|false|C0575044|Joint problem|Joint
Finding|Physiologic Function|General Exam|5520,5540|false|false|false|C0423561|Joint position sense|Joint position sense
Finding|Organism Function|General Exam|5526,5540|false|false|false|C0234219|Position Sense|position sense
Event|Event|General Exam|5535,5540|false|false|false|||sense
Finding|Organ or Tissue Function|General Exam|5535,5540|false|false|false|C0036658|Sensory perception|sense
Event|Event|General Exam|5541,5547|false|false|false|||intact
Finding|Finding|General Exam|5541,5547|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Gene or Genome|General Exam|5555,5560|false|false|false|C1424898|RXFP2 gene|great
Anatomy|Body Part, Organ, or Organ Component|General Exam|5555,5565|false|false|false|C0018534|Hallux structure|great toes
Anatomy|Body Part, Organ, or Organ Component|General Exam|5561,5565|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Event|Event|General Exam|5570,5580|false|false|false|||extinction
Finding|Mental Process|General Exam|5570,5580|true|false|false|C0015347|Extinction, Psychological|extinction
Disorder|Disease or Syndrome|General Exam|5584,5587|false|false|false|C0011195;C1848296|DOSAGE-SENSITIVE SEX REVERSAL;Dejerine-Sottas Disease|DSS
Drug|Organic Chemical|General Exam|5584,5587|false|false|false|C0719637|DSS brand of docusate sodium|DSS
Drug|Pharmacologic Substance|General Exam|5584,5587|false|false|false|C0719637|DSS brand of docusate sodium|DSS
Event|Event|General Exam|5584,5587|false|false|false|||DSS
Finding|Gene or Genome|General Exam|5584,5587|false|false|false|C1417820;C2698419;C2698698;C5890838|MPZ wt Allele;NR0B1 gene;NR0B1 wt Allele;PMP22 wt Allele|DSS
Disorder|Disease or Syndrome|General Exam|5589,5596|false|false|false|C0015458|Facial Hemiatrophy|Romberg
Event|Event|General Exam|5589,5596|false|false|false|||Romberg
Finding|Functional Concept|General Exam|5597,5603|false|false|false|C0332197|Absent|absent
Lab|Laboratory or Test Result|General Exam|5597,5603|false|false|false|C5237010|Expression Negative|absent
Event|Event|General Exam|5607,5615|false|false|false|||Reflexes
Finding|Finding|General Exam|5607,5615|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Finding|Organ or Tissue Function|General Exam|5607,5615|false|false|false|C0034929;C0596002|Observation of reflex;Reflex action|Reflexes
Procedure|Diagnostic Procedure|General Exam|5607,5615|false|false|false|C0436145|Examination of reflexes|Reflexes
Anatomy|Body Part, Organ, or Organ Component|General Exam|5620,5623|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|General Exam|5620,5623|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|General Exam|5620,5623|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|General Exam|5620,5623|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|General Exam|5620,5623|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|General Exam|5626,5629|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|5626,5629|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Disorder|Disease or Syndrome|General Exam|5638,5641|false|false|false|C0030587|Paroxysmal atrial tachycardia|Pat
Drug|Organic Chemical|General Exam|5638,5641|false|false|false|C2825250|Fenamole|Pat
Drug|Pharmacologic Substance|General Exam|5638,5641|false|false|false|C2825250|Fenamole|Pat
Event|Event|General Exam|5638,5641|false|false|false|||Pat
Finding|Molecular Function|General Exam|5638,5641|false|false|false|C2247344;C2247346;C2248827|aspartate-prephenate aminotransferase activity;glutamate-prephenate aminotransferase activity;protein acetyltransferase activity|Pat
Procedure|Diagnostic Procedure|General Exam|5638,5641|false|false|false|C3897364|Thermoacoustic Computed Tomography|Pat
Disorder|Congenital Abnormality|General Exam|5644,5647|false|false|false|C0001080|Achondroplasia|Ach
Drug|Biologically Active Substance|General Exam|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Drug|Organic Chemical|General Exam|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Drug|Pharmacologic Substance|General Exam|5644,5647|false|false|false|C0001041|acetylcholine|Ach
Event|Event|General Exam|5644,5647|false|false|false|||Ach
Finding|Gene or Genome|General Exam|5644,5647|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Finding|Sign or Symptom|General Exam|5644,5647|false|false|false|C0234238;C1333543;C1705145|Ache;FGFR3 gene;FGFR3 wt Allele|Ach
Anatomy|Body Location or Region|General Exam|5714,5721|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|Plantar
Event|Event|General Exam|5722,5730|false|false|false|||response
Finding|Finding|General Exam|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Intellectual Product|General Exam|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Finding|Mental Process|General Exam|5722,5730|false|false|false|C1704632;C1706817;C2911692|Answer (statement);Communication Response;Disease Response|response
Anatomy|Body Location or Region|General Exam|5735,5741|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Event|Event|General Exam|5757,5769|false|false|false|||Coordination
Finding|Functional Concept|General Exam|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|5757,5769|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|General Exam|5774,5783|false|false|false|||intention
Finding|Mental Process|General Exam|5774,5783|false|false|false|C0162425||intention
Finding|Sign or Symptom|General Exam|5774,5790|true|false|false|C0234376;C4551520|Action Tremor;Intention tremor|intention tremor
Event|Event|General Exam|5784,5790|false|false|false|||tremor
Finding|Sign or Symptom|General Exam|5784,5790|true|false|false|C0040822|Tremor|tremor
Event|Event|General Exam|5796,5805|false|false|false|||dysmetria
Finding|Finding|General Exam|5796,5805|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Drug|Organic Chemical|General Exam|5809,5812|false|false|false|C0033228|fenofibrate|FNF
Drug|Pharmacologic Substance|General Exam|5809,5812|false|false|false|C0033228|fenofibrate|FNF
Event|Event|General Exam|5809,5812|false|false|false|||FNF
Event|Event|General Exam|5826,5829|false|false|false|||HKS
Anatomy|Body Part, Organ, or Organ Component|General Exam|5837,5841|false|false|false|C0018870|Heel|heel
Event|Event|General Exam|5850,5859|false|false|false|||dysmetria
Finding|Finding|General Exam|5850,5859|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Event|Event|General Exam|5861,5867|false|false|false|||Unable
Finding|Finding|General Exam|5861,5867|false|false|false|C1299582|Unable|Unable
Event|Event|General Exam|5871,5875|false|false|false|||bend
Anatomy|Body Location or Region|General Exam|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|5878,5882|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|5878,5882|false|false|false|C0562271|Examination of knee joint|knee
Anatomy|Body Location or Region|General Exam|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Anatomy|Body Space or Junction|General Exam|5890,5894|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|knee
Procedure|Diagnostic Procedure|General Exam|5890,5894|false|false|false|C0562271|Examination of knee joint|knee
Procedure|Therapeutic or Preventive Procedure|General Exam|5890,5902|false|false|false|C0187769|Operative procedure on knee|knee surgery
Event|Event|General Exam|5895,5902|false|false|false|||surgery
Finding|Finding|General Exam|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|General Exam|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|General Exam|5895,5902|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|General Exam|5895,5902|false|false|false|C0543467|Operative Surgical Procedures|surgery
Finding|Finding|General Exam|5907,5911|false|false|false|C0016928|Gait|Gait
Event|Event|General Exam|5913,5919|false|false|false|||unable
Finding|Finding|General Exam|5913,5919|false|false|false|C1299582|Unable|unable
Event|Event|General Exam|5923,5929|false|false|false|||assess
Finding|Body Substance|General Exam|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5933,5940|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5941,5946|false|false|false|||needs
Event|Event|General Exam|5949,5955|false|false|false|||walker
Drug|Biomedical or Dental Material|General Exam|5959,5967|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|5959,5967|false|false|false|||baseline
Finding|Idea or Concept|General Exam|5959,5967|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Body Substance|General Exam|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|5969,5978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|5969,5978|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|5979,5983|false|false|false|||EXAM
Finding|Functional Concept|General Exam|5979,5983|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|5979,5983|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|5991,5995|false|false|false|||Data
Finding|Idea or Concept|General Exam|5991,5995|false|false|false|C1511726|Data|Data
Event|Event|General Exam|6002,6009|false|false|false|||updated
Event|Event|General Exam|6021,6025|false|false|false|||Temp
Finding|Gene or Genome|General Exam|6021,6025|false|false|false|C1823816|C1orf210 gene|Temp
Procedure|Therapeutic or Preventive Procedure|General Exam|6021,6025|false|false|false|C0279848|Tamoxifen/Etoposide/Mitoxantrone/Cisplatin Regimen|Temp
Event|Event|General Exam|6088,6090|false|false|false|||RR
Event|Event|General Exam|6126,6134|false|false|false|||delivery
Finding|Finding|General Exam|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Functional Concept|General Exam|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Finding|Organism Function|General Exam|6126,6134|false|false|false|C1314680;C1705822;C2053584|Transfer Technique;delivery (history)|delivery
Procedure|Therapeutic or Preventive Procedure|General Exam|6126,6134|false|false|false|C0011209|Obstetric Delivery|delivery
Event|Event|General Exam|6140,6147|false|false|false|||General
Finding|Classification|General Exam|6140,6147|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|6140,6147|false|false|false|C3812897|General medical service|General
Event|Event|General Exam|6149,6154|false|false|false|||Awake
Finding|Finding|General Exam|6149,6154|false|false|false|C0234422|Awake (finding)|Awake
Disorder|Disease or Syndrome|General Exam|6183,6186|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|6183,6186|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|6183,6186|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Event|Event|General Exam|6183,6186|false|false|false|||NAD
Finding|Finding|General Exam|6183,6186|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|6188,6193|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|6205,6212|false|false|false|C0036410|Sclera|scleral
Finding|Finding|General Exam|6205,6220|true|false|false|C0240962|Scleral icterus|scleral icterus
Event|Event|General Exam|6213,6220|false|false|false|||icterus
Finding|Sign or Symptom|General Exam|6213,6220|true|false|false|C0022346|Icterus|icterus
Event|Event|General Exam|6221,6226|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|6228,6231|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|6228,6231|false|false|false|C0026987|Myelofibrosis|MMM
Event|Event|General Exam|6236,6243|false|false|false|||lesions
Finding|Finding|General Exam|6236,6243|true|false|false|C0221198|Lesion|lesions
Event|Event|General Exam|6244,6249|false|false|false|||noted
Anatomy|Body Location or Region|General Exam|6253,6263|false|false|false|C0521367|Oropharyngeal|oropharynx
Anatomy|Body Location or Region|General Exam|6265,6269|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|6265,6269|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|6265,6269|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|6271,6277|false|false|false|||Supple
Finding|Functional Concept|General Exam|6271,6277|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|6282,6297|true|false|false|C1320474|Nuchal Rigidity|nuchal rigidity
Event|Event|General Exam|6289,6297|false|false|false|||rigidity
Finding|Sign or Symptom|General Exam|6289,6297|true|false|false|C0026837|Muscle Rigidity|rigidity
Phenomenon|Natural Phenomenon or Process|General Exam|6289,6297|true|false|false|C0700109|plastic property - rigidity|rigidity
Anatomy|Body Part, Organ, or Organ Component|General Exam|6299,6308|false|false|false|C0024109|Lung|Pulmonary
Attribute|Clinical Attribute|General Exam|6299,6308|false|false|false|C2707265||Pulmonary
Finding|Finding|General Exam|6299,6308|false|false|false|C4522268|Pulmonary (intended site)|Pulmonary
Event|Event|General Exam|6317,6321|false|false|false|||work
Event|Occupational Activity|General Exam|6317,6321|false|false|false|C0043227|Work|work
Finding|Organ or Tissue Function|General Exam|6317,6334|false|false|false|C0043229|Work of Breathing|work of breathing
Attribute|Clinical Attribute|General Exam|6325,6334|false|false|false|C5885990||breathing
Event|Event|General Exam|6325,6334|false|false|false|||breathing
Finding|Finding|General Exam|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|General Exam|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|General Exam|6325,6334|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|General Exam|6325,6334|false|false|false|C1160636|respiratory system process|breathing
Anatomy|Body Part, Organ, or Organ Component|General Exam|6336,6343|false|false|false|C0018787|Heart|Cardiac
Finding|Intellectual Product|General Exam|6336,6343|false|false|false|C1314974|Cardiac attachment|Cardiac
Finding|Finding|General Exam|6353,6357|false|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|6353,6357|false|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|6359,6363|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|6364,6372|false|false|false|||perfused
Anatomy|Body Location or Region|General Exam|6374,6381|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|6374,6381|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Event|Event|General Exam|6374,6381|false|false|false|||Abdomen
Finding|Finding|General Exam|6374,6381|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|6383,6387|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|6383,6387|false|false|false|||Soft
Anatomy|Body Part, Organ, or Organ Component|General Exam|6404,6415|false|false|false|C0015385;C0278454|All extremities;Limb structure|Extremities
Attribute|Clinical Attribute|General Exam|6424,6429|false|false|false|C1717255||edema
Event|Event|General Exam|6424,6429|false|false|false|||edema
Finding|Pathologic Function|General Exam|6424,6429|false|false|false|C0013604|Edema|edema
Anatomy|Body System|General Exam|6431,6435|false|false|false|C1123023;C4520765|Skin;Skin, Human|Skin
Disorder|Disease or Syndrome|General Exam|6431,6435|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Disorder|Neoplastic Process|General Exam|6431,6435|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|Skin
Finding|Body Substance|General Exam|6431,6435|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Finding|Intellectual Product|General Exam|6431,6435|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|Skin
Event|Event|General Exam|6437,6447|false|false|false|||ecchymoses
Finding|Pathologic Function|General Exam|6437,6447|false|false|false|C0013491|Ecchymosis|ecchymoses
Anatomy|Body Location or Region|General Exam|6453,6457|false|false|false|C0230444|Shin|shin
Event|Event|General Exam|6464,6473|false|false|false|||extensive
Anatomy|Body Location or Region|General Exam|6479,6483|false|false|false|C0230444|Shin|shin
Finding|Mental Process|General Exam|6501,6507|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|6501,6514|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|General Exam|6501,6514|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|General Exam|6508,6514|false|false|false|C5889824||Status
Event|Event|General Exam|6508,6514|false|false|false|||Status
Finding|Idea or Concept|General Exam|6508,6514|false|false|false|C1546481|What subject filter - Status|Status
Attribute|Clinical Attribute|General Exam|6516,6521|false|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|6516,6521|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|6516,6521|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|6516,6521|false|false|false|||Alert
Finding|Finding|General Exam|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|6516,6521|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|6523,6531|false|false|false|||oriented
Attribute|Clinical Attribute|General Exam|6535,6541|false|false|false|C5890614||person
Event|Event|General Exam|6535,6541|false|false|false|||person
Finding|Intellectual Product|General Exam|6535,6541|false|false|false|C1522390|Person Info|person
Event|Event|General Exam|6546,6555|false|false|false|||situation
Finding|Finding|General Exam|6557,6561|false|false|false|C1299581|Able (qualifier value)|Able
Drug|Organic Chemical|General Exam|6565,6571|false|false|false|C0163712|Relate - vinyl resin|relate
Event|Event|General Exam|6572,6579|false|false|false|||history
Finding|Conceptual Entity|General Exam|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|General Exam|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|General Exam|6572,6579|false|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Event|Event|General Exam|6600,6609|false|false|false|||Attentive
Event|Event|General Exam|6613,6621|false|false|false|||examiner
Attribute|Clinical Attribute|General Exam|6623,6631|false|false|false|C2706915||Language
Event|Event|General Exam|6623,6631|false|false|false|||Language
Finding|Intellectual Product|General Exam|6623,6631|false|false|false|C0033348|Programming Languages|Language
Event|Event|General Exam|6635,6641|false|false|false|||fluent
Event|Event|General Exam|6647,6653|false|false|false|||intact
Finding|Finding|General Exam|6647,6653|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|6654,6667|false|false|false|||comprehension
Finding|Mental Process|General Exam|6654,6667|false|false|false|C0162340|Comprehension|comprehension
Event|Event|General Exam|6676,6683|false|false|false|||prosody
Finding|Finding|General Exam|6676,6683|false|false|false|C0233743|Prosody|prosody
Event|Event|General Exam|6710,6716|false|false|false|||errors
Disorder|Mental or Behavioral Dysfunction|General Exam|6721,6731|true|false|false|C0013362|Dysarthria|dysarthria
Event|Event|General Exam|6721,6731|false|false|false|||dysarthria
Event|Event|General Exam|6733,6737|false|false|false|||Able
Finding|Finding|General Exam|6733,6737|false|false|false|C1299581|Able (qualifier value)|Able
Event|Event|General Exam|6741,6747|false|false|false|||follow
Finding|Functional Concept|General Exam|6741,6747|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Finding|Intellectual Product|General Exam|6741,6747|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|follow
Anatomy|Cell Component|General Exam|6753,6760|false|false|false|C1660780|midline cell component|midline
Event|Event|General Exam|6778,6786|false|false|false|||commands
Event|Event|General Exam|6801,6809|false|false|false|||evidence
Finding|Idea or Concept|General Exam|6801,6809|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|6801,6812|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Mental or Behavioral Dysfunction|General Exam|6813,6820|false|false|false|C0003635|Apraxias|apraxia
Event|Event|General Exam|6813,6820|false|false|false|||apraxia
Event|Event|General Exam|6824,6831|false|false|false|||neglect
Event|Event|General Exam|6824,6831|false|false|false|C5969868|Neglect (event)|neglect
Finding|Finding|General Exam|6824,6831|false|false|false|C0521874|Victim of neglect (finding)|neglect
Anatomy|Body Part, Organ, or Organ Component|General Exam|6835,6842|false|false|false|C0037303|Bone structure of cranium|Cranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|6835,6849|false|false|false|C0010268|Cranial Nerves|Cranial Nerves
Disorder|Neoplastic Process|General Exam|6835,6849|false|false|false|C0004992;C0496937|Benign neoplasm of cranial nerves;Neoplasm of uncertain or unknown behavior of cranial nerves|Cranial Nerves
Anatomy|Body Part, Organ, or Organ Component|General Exam|6843,6849|false|false|false|C0027740|Nerve|Nerves
Finding|Finding|General Exam|6869,6874|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Event|Event|General Exam|6895,6899|false|false|false|||EOMI
Disorder|Disease or Syndrome|General Exam|6908,6917|false|false|false|C0028738|Nystagmus|nystagmus
Event|Event|General Exam|6908,6917|false|false|false|||nystagmus
Event|Event|General Exam|6926,6934|false|false|false|||saccades
Finding|Finding|General Exam|6926,6934|false|false|false|C0036019|Saccades|saccades
Anatomy|Body Location or Region|General Exam|6939,6945|false|false|false|C0015450|Face|Facial
Finding|Finding|General Exam|6939,6955|false|false|false|C0517999|facial sensation|Facial sensation
Event|Event|General Exam|6946,6955|false|false|false|||sensation
Finding|Finding|General Exam|6946,6955|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|6946,6955|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|6946,6955|false|false|false|C2229507|sensory exam|sensation
Event|Event|General Exam|6956,6962|false|false|false|||intact
Finding|Finding|General Exam|6956,6962|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Amino Acid, Peptide, or Protein|General Exam|6966,6971|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|6966,6971|false|false|false|C1570446|TNFSF14 protein, human|light
Event|Event|General Exam|6966,6971|false|false|false|||light
Finding|Finding|General Exam|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|6966,6971|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|6966,6971|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|6966,6971|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|6966,6977|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|6972,6977|false|false|false|||touch
Finding|Mental Process|General Exam|6972,6977|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|6972,6977|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|6972,6977|false|false|false|C0152054|Therapeutic Touch|touch
Anatomy|Body Part, Organ, or Organ Component|General Exam|6979,6982|false|false|false|C2338708;C3496273;C3496274|Lamina VII of gray matter of spinal cord;layer VII (Cajal);lobule VII|VII
Finding|Intellectual Product|General Exam|6979,6982|false|false|false|C0445385|Roman numeral VII|VII
Anatomy|Body Location or Region|General Exam|6987,6993|false|false|false|C0015450|Face|facial
Disorder|Disease or Syndrome|General Exam|6987,6999|true|false|false|C0427055|Facial Paresis|facial droop
Finding|Finding|General Exam|6987,6999|true|false|false|C4022719|Unilateral facial palsy|facial droop
Event|Event|General Exam|6994,6999|false|false|false|||droop
Anatomy|Body Location or Region|General Exam|7001,7007|false|false|false|C0015450|Face|facial
Anatomy|Body Part, Organ, or Organ Component|General Exam|7008,7019|false|false|false|C1995013|Set of muscles|musculature
Event|Event|General Exam|7020,7029|false|false|false|||symmetric
Finding|Conceptual Entity|General Exam|7020,7029|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Finding|Finding|General Exam|7020,7029|false|false|false|C0332516;C2699744|Symmetric Relationship;Symmetrical|symmetric
Anatomy|Body Part, Organ, or Organ Component|General Exam|7031,7035|false|false|false|C0228488;C2327388|Cerebellar pyramis;Lamina VIII of gray matter of spinal cord|VIII
Finding|Gene or Genome|General Exam|7031,7035|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Intellectual Product|General Exam|7031,7035|false|false|false|C0445599;C1413661|COX8A gene;Roman numeral VIII|VIII
Finding|Finding|General Exam|7037,7044|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Finding|Physiologic Function|General Exam|7037,7044|false|false|false|C0018767;C1455844;C2015933|Hearing;Hearing finding;outcomes otolaryngology hearing|Hearing
Event|Event|General Exam|7045,7051|false|false|false|||intact
Finding|Finding|General Exam|7045,7051|false|false|false|C1554187|Gender Status - Intact|intact
Event|Event|General Exam|7055,7067|false|false|false|||conversation
Finding|Social Behavior|General Exam|7055,7067|false|false|false|C0871703|conversation|conversation
Anatomy|Body Part, Organ, or Organ Component|General Exam|7076,7082|false|false|false|C0700374|Palate|Palate
Event|Event|General Exam|7083,7091|false|false|false|||elevates
Event|Event|General Exam|7115,7123|false|false|false|||strength
Finding|Idea or Concept|General Exam|7115,7123|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|7154,7160|false|false|false|C0040408|Tongue|Tongue
Disorder|Neoplastic Process|General Exam|7154,7160|false|false|false|C0153933|Benign neoplasm of tongue|Tongue
Event|Event|General Exam|7154,7160|false|false|false|||Tongue
Procedure|Health Care Activity|General Exam|7154,7160|false|false|false|C0872394|Procedure on tongue|Tongue
Event|Event|General Exam|7161,7170|false|false|false|||protrudes
Anatomy|Cell Component|General Exam|7174,7181|false|false|false|C1660780|midline cell component|midline
Finding|Idea or Concept|General Exam|7187,7191|false|false|false|C1551023;C1610541|Language Ability Proficiency - Good;Language Proficiency - Good|good
Event|Event|General Exam|7192,7202|false|false|false|||excursions
Finding|Functional Concept|General Exam|7206,7211|false|false|false|C1513492|motor movement|Motor
Drug|Biomedical or Dental Material|General Exam|7220,7224|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Drug|Food|General Exam|7220,7224|false|false|false|C0012173;C1337615|Bulk (conceptual);Dietary Fiber|bulk
Event|Event|General Exam|7229,7233|false|false|false|||tone
Finding|Pathologic Function|General Exam|7249,7263|true|false|false|C1504476|Pronator drift|pronator drift
Event|Event|General Exam|7258,7263|false|false|false|||drift
Event|Event|General Exam|7281,7290|false|false|false|||movements
Finding|Organism Function|General Exam|7281,7290|false|false|false|C0026649|Movement|movements
Event|Event|General Exam|7300,7306|false|false|false|||tremor
Finding|Sign or Symptom|General Exam|7300,7306|false|false|false|C0040822|Tremor|tremor
Event|Event|General Exam|7310,7319|false|false|false|||asterixis
Finding|Sign or Symptom|General Exam|7310,7319|false|false|false|C0232766|Asterixis|asterixis
Event|Event|General Exam|7320,7325|false|false|false|||noted
Anatomy|Body Part, Organ, or Organ Component|General Exam|7330,7334|false|false|false|C0224234|Structure of deltoid muscle|Delt
Anatomy|Body Part, Organ, or Organ Component|General Exam|7336,7339|false|false|false|C0175372;C3495985|Structure of inferior brachium of corpora quadrigemina;nucleus of the brachium of the inferior colliculus|Bic
Drug|Organic Chemical|General Exam|7336,7339|false|false|false|C0063382|imidazole mustard|Bic
Drug|Pharmacologic Substance|General Exam|7336,7339|false|false|false|C0063382|imidazole mustard|Bic
Finding|Gene or Genome|General Exam|7336,7339|false|false|false|C1537811;C2681931|MIR155 gene;MIR155HG gene|Bic
Procedure|Therapeutic or Preventive Procedure|General Exam|7336,7339|false|false|false|C5202575|BIC Regimen|Bic
Finding|Gene or Genome|General Exam|7341,7344|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Intellectual Product|General Exam|7341,7344|false|false|false|C0814229;C3891460|TRI-AAT9-1 gene;Temptation and Restraint Inventory|Tri
Finding|Gene or Genome|General Exam|7351,7354|false|false|false|C1537570;C3539626|LGR5 gene;LGR5 wt Allele|FEx
Disorder|Disease or Syndrome|General Exam|7370,7373|false|false|false|C0030481|Tropical Spastic Paraparesis|Ham
Drug|Amino Acid, Peptide, or Protein|General Exam|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Drug|Biologically Active Substance|General Exam|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Drug|Food|General Exam|7370,7373|false|false|false|C1570167;C3853311|ATF7IP protein, human;Ham|Ham
Event|Event|General Exam|7370,7373|false|false|false|||Ham
Procedure|Therapeutic or Preventive Procedure|General Exam|7370,7373|false|false|false|C0279477|altretamine/doxorubicin/melphalan protocol|Ham
Drug|Biomedical or Dental Material|General Exam|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Drug|Chemical Viewed Structurally|General Exam|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Drug|Substance|General Exam|7379,7382|false|false|false|C0017110;C1550641;C1704673|Gas - SpecimenType;Gas Dosage Form;Gases|Gas
Finding|Gene or Genome|General Exam|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Intellectual Product|General Exam|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Molecular Function|General Exam|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Finding|Sign or Symptom|General Exam|7379,7382|false|false|false|C0596601;C1414950;C1439341;C1540252;C1546643;C2266618;C2986619;C3812826;C5890923|GALNS gene;GALNS wt Allele;GAST gene;GAST wt Allele;Gas - Specimen Source Codes;PAGR1 gene;PAGR1 wt Allele;gastrointestinal gas;germacrene-A synthase activity|Gas
Event|Event|General Exam|7496,7497|false|false|false|||5
Anatomy|Body Location or Region|General Exam|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Part, Organ, or Organ Component|General Exam|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Anatomy|Body Space or Junction|General Exam|7503,7507|false|false|false|C0022742;C0022745;C1963703;C4299094|Knee;Knee joint;Knee region structure;Lower extremity>Knee|Knee
Procedure|Diagnostic Procedure|General Exam|7503,7507|false|false|false|C0562271|Examination of knee joint|Knee
Event|Event|General Exam|7515,7519|false|false|false|||bend
Finding|Finding|General Exam|7526,7539|false|true|false|C0455610|History of surgery|prior surgery
Event|Event|General Exam|7532,7539|false|false|false|||surgery
Finding|Finding|General Exam|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Functional Concept|General Exam|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Finding|Idea or Concept|General Exam|7532,7539|false|false|false|C0038895;C1457907;C1547138|Level of Care - Surgery;Surgical aspects;Surgical procedure finding|surgery
Procedure|Therapeutic or Preventive Procedure|General Exam|7532,7539|false|false|false|C0543467|Operative Surgical Procedures|surgery
Event|Event|General Exam|7554,7562|false|false|false|||deficits
Drug|Amino Acid, Peptide, or Protein|General Exam|7566,7571|false|false|false|C1570446|TNFSF14 protein, human|light
Drug|Biologically Active Substance|General Exam|7566,7571|false|false|false|C1570446|TNFSF14 protein, human|light
Finding|Finding|General Exam|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Functional Concept|General Exam|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Finding|Gene or Genome|General Exam|7566,7571|false|false|false|C1306462;C1420817;C3842678;C4521367|Light - subjective measurement;Light color;TNFSF14 gene;TNFSF14 wt Allele|light
Phenomenon|Natural Phenomenon or Process|General Exam|7566,7571|false|false|false|C0023693|Light|light
Procedure|Therapeutic or Preventive Procedure|General Exam|7566,7571|false|false|false|C0031765|Phototherapy|light
Finding|Physiologic Function|General Exam|7566,7577|false|false|false|C0423553|Light touch|light touch
Event|Event|General Exam|7572,7577|false|false|false|||touch
Finding|Mental Process|General Exam|7572,7577|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|7572,7577|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|7572,7577|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|General Exam|7592,7604|false|false|false|||Coordination
Finding|Functional Concept|General Exam|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Idea or Concept|General Exam|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Finding|Physiologic Function|General Exam|7592,7604|false|false|false|C0242414;C0700114;C1549570|Coordinated;Coordination of Benefits - Coordination;Physiologic Coordination|Coordination
Event|Event|General Exam|7609,7618|false|false|false|||intention
Finding|Mental Process|General Exam|7609,7618|false|false|false|C0162425||intention
Finding|Sign or Symptom|General Exam|7609,7625|true|false|false|C0234376;C4551520|Action Tremor;Intention tremor|intention tremor
Event|Event|General Exam|7619,7625|false|false|false|||tremor
Finding|Sign or Symptom|General Exam|7619,7625|true|false|false|C0040822|Tremor|tremor
Event|Event|General Exam|7631,7640|false|false|false|||dysmetria
Finding|Finding|General Exam|7631,7640|true|false|false|C0234162|Cerebellar Dysmetria|dysmetria
Drug|Organic Chemical|General Exam|7644,7647|false|false|false|C0033228|fenofibrate|FNF
Drug|Pharmacologic Substance|General Exam|7644,7647|false|false|false|C0033228|fenofibrate|FNF
Event|Event|General Exam|7644,7647|false|false|false|||FNF
Finding|Finding|General Exam|7664,7668|false|false|false|C0016928|Gait|Gait
Event|Event|General Exam|7670,7675|false|false|false|||needs
Event|Event|General Exam|7678,7684|false|false|false|||walker
Drug|Biomedical or Dental Material|General Exam|7688,7696|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|7688,7696|false|false|false|||baseline
Finding|Idea or Concept|General Exam|7688,7696|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|General Exam|7730,7735|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7730,7735|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7730,7735|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|7736,7739|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|7744,7747|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|7744,7747|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|7744,7747|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|7753,7756|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|7753,7756|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|7753,7756|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|7753,7756|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|7762,7765|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|7762,7765|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|7773,7776|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|7773,7776|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|7773,7776|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|7773,7776|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|7773,7776|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|7780,7783|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|7780,7783|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|7780,7783|false|false|false|||MCH
Finding|Gene or Genome|General Exam|7780,7783|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|7780,7783|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|7780,7783|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Event|Event|General Exam|7789,7793|false|false|false|||MCHC
Procedure|Laboratory Procedure|General Exam|7789,7793|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|7820,7823|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|7840,7845|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7840,7845|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7840,7845|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Antibiotic|General Exam|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|7861,7866|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|7871,7874|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Event|Event|General Exam|7871,7874|false|false|false|||Eos
Finding|Gene or Genome|General Exam|7871,7874|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|7973,7978|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|7973,7978|false|false|false|||BLOOD
Finding|Body Substance|General Exam|7973,7978|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|7983,7986|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|7983,7986|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|7983,7986|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|8008,8013|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8008,8013|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8008,8013|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|8008,8021|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|8008,8021|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|8008,8021|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|8014,8021|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|8014,8021|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|8014,8021|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|8014,8021|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|8014,8021|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|8014,8021|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|8065,8069|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|8065,8069|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|8065,8069|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|8094,8099|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8094,8099|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8094,8099|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|8100,8105|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Drug|Enzyme|General Exam|8100,8105|false|false|false|C0010290|Creatine Kinase MB Isoenzyme|CK-MB
Finding|Molecular Function|General Exam|8100,8105|false|false|false|C1150462|creatine kinase activity|CK-MB
Procedure|Laboratory Procedure|General Exam|8100,8105|false|false|false|C0455293;C0523584|Creatine kinase MB measurement;Serum creatine phosphokinase MB isoenzyme measurement|CK-MB
Disorder|Disease or Syndrome|General Exam|8134,8139|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8134,8139|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8134,8139|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|8134,8147|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|8140,8147|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|8140,8147|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|8140,8147|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|8140,8147|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|8193,8198|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8193,8198|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8193,8198|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|8210,8213|false|false|false|C0023821|High Density Lipoproteins|HDL
Drug|Biologically Active Substance|General Exam|8210,8213|false|false|false|C0023821|High Density Lipoproteins|HDL
Event|Event|General Exam|8210,8213|false|false|false|||HDL
Finding|Gene or Genome|General Exam|8210,8213|false|false|false|C3715113|HSD11B1 wt Allele|HDL
Procedure|Laboratory Procedure|General Exam|8210,8213|false|false|false|C0392885|High density lipoprotein measurement|HDL
Event|Event|General Exam|8217,8221|false|false|false|||CHOL
Disorder|Disease or Syndrome|General Exam|8253,8258|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8253,8258|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8253,8258|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|8260,8265|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Drug|Biologically Active Substance|General Exam|8260,8265|false|false|false|C0019018|Glycosylated hemoglobin A|HbA1c
Event|Event|General Exam|8260,8265|false|false|false|||HbA1c
Procedure|Laboratory Procedure|General Exam|8260,8265|false|false|false|C0202054|Glucohemoglobin measurement|HbA1c
Finding|Gene or Genome|General Exam|8270,8273|false|false|false|C1416571|KCNH1 gene|eAG
Disorder|Disease or Syndrome|General Exam|8290,8295|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8290,8295|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8290,8295|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Disease or Syndrome|General Exam|8319,8324|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8319,8324|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8319,8324|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Attribute|Clinical Attribute|General Exam|8325,8328|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|General Exam|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|General Exam|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|General Exam|8325,8328|false|false|false|C0040160|thyrotropin|TSH
Event|Event|General Exam|8325,8328|false|false|false|||TSH
Procedure|Laboratory Procedure|General Exam|8325,8328|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Disorder|Disease or Syndrome|General Exam|8346,8351|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|8346,8351|false|false|false|||BLOOD
Finding|Body Substance|General Exam|8346,8351|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Event|Event|General Exam|8360,8363|false|false|false|||NEG
Finding|Finding|General Exam|8360,8363|false|false|false|C5848551|Neg - answer|NEG
Finding|Body Substance|General Exam|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|8376,8381|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Finding|General Exam|8376,8387|false|false|false|C0278030|Color of urine|URINE Color
Drug|Biomedical or Dental Material|General Exam|8382,8387|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Indicator, Reagent, or Diagnostic Aid|General Exam|8382,8387|false|false|false|C1550604;C1705245|Coloring Excipient;color additive|Color
Drug|Organic Chemical|General Exam|8388,8393|false|false|false|C4047917|Cereal plant straw|Straw
Finding|Idea or Concept|General Exam|8401,8406|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Body Substance|General Exam|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Functional Concept|General Exam|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Finding|Intellectual Product|General Exam|8426,8431|false|false|false|C0042036;C0042037;C1547942;C1610733;C2963137|In Urine;Portion of urine;Urine;Urine specimen|URINE
Disorder|Disease or Syndrome|General Exam|8426,8437|false|false|false|C0018965|Hematuria|URINE Blood
Disorder|Disease or Syndrome|General Exam|8432,8437|false|false|false|C0851353|Blood and lymphatic system disorders|Blood
Finding|Body Substance|General Exam|8432,8437|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|Blood
Event|Event|General Exam|8438,8441|false|false|false|||NEG
Finding|Finding|General Exam|8438,8441|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Inorganic Chemical|General Exam|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Drug|Pharmacologic Substance|General Exam|8442,8449|false|false|false|C0028137;C3848529|Nitrites;nitrite ion|Nitrite
Event|Event|General Exam|8450,8453|false|false|false|||NEG
Finding|Finding|General Exam|8450,8453|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|8454,8461|false|false|false|C0033684|Proteins|Protein
Drug|Biologically Active Substance|General Exam|8454,8461|false|false|false|C0033684|Proteins|Protein
Event|Event|General Exam|8454,8461|false|false|false|||Protein
Finding|Conceptual Entity|General Exam|8454,8461|false|false|false|C1521746|Protein Info|Protein
Procedure|Laboratory Procedure|General Exam|8454,8461|false|false|false|C0202202|Protein measurement|Protein
Event|Event|General Exam|8462,8465|false|false|false|||NEG
Finding|Finding|General Exam|8462,8465|false|false|false|C5848551|Neg - answer|NEG
Drug|Biologically Active Substance|General Exam|8467,8474|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|8467,8474|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|8467,8474|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|8467,8474|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|8467,8474|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|8467,8474|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|8475,8478|false|false|false|||NEG
Finding|Finding|General Exam|8475,8478|false|false|false|C5848551|Neg - answer|NEG
Drug|Organic Chemical|General Exam|8479,8485|false|false|false|C0022634|Ketones|Ketone
Event|Event|General Exam|8486,8489|false|false|false|||NEG
Finding|Finding|General Exam|8486,8489|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|8498,8501|false|false|false|C5848551|Neg - answer|NEG
Finding|Finding|General Exam|8510,8513|false|false|false|C5848551|Neg - answer|NEG
Event|Event|General Exam|8527,8530|false|false|false|||NEG
Finding|Finding|General Exam|8527,8530|false|false|false|C5848551|Neg - answer|NEG
Drug|Amino Acid, Peptide, or Protein|General Exam|8540,8543|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|General Exam|8540,8543|false|false|false|||CTA
Finding|Gene or Genome|General Exam|8540,8543|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|General Exam|8540,8543|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|General Exam|8544,8548|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|8544,8548|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|General Exam|8544,8548|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|General Exam|8544,8548|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|General Exam|8549,8553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|General Exam|8549,8553|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|General Exam|8549,8553|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|General Exam|8558,8565|false|false|false|||opinion
Finding|Idea or Concept|General Exam|8558,8565|false|false|false|C0871010|Opinions|opinion
Finding|Functional Concept|Impression|8599,8603|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|8599,8620|false|false|false|C0226231|Structure of left vertebral artery|left vertebral artery
Finding|Pathologic Function|Impression|8599,8630|false|false|false|C4536452|Occlusion of left vertebral artery (disorder)|left vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|Impression|8604,8613|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Location or Region|Impression|8604,8620|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Anatomy|Body Part, Organ, or Organ Component|Impression|8604,8620|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Finding|Pathologic Function|Impression|8604,8630|false|false|false|C0265104|Vertebral artery obstruction (disorder)|vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|Impression|8614,8620|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Impression|8614,8620|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Pathologic Function|Impression|8614,8630|false|false|false|C0264995|Occlusion of artery (disorder)|artery occlusion
Disorder|Acquired Abnormality|Impression|8621,8630|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|Impression|8621,8630|false|false|false|||occlusion
Finding|Finding|Impression|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Impression|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Impression|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Impression|8621,8630|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|Impression|8634,8647|false|false|false|||indeterminate
Event|Event|Impression|8649,8659|false|false|false|||chronicity
Event|Event|Impression|8665,8673|false|false|false|||evidence
Finding|Idea or Concept|Impression|8665,8673|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|8665,8676|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Event|Event|Impression|8677,8685|false|false|false|||ischemia
Finding|Pathologic Function|Impression|8677,8685|true|false|false|C0022116|Ischemia|ischemia
Procedure|Therapeutic or Preventive Procedure|Impression|8677,8685|true|false|false|C4321499|Ischemia Procedure|ischemia
Finding|Finding|Impression|8691,8699|false|false|false|C2984079|Somewhat|Somewhat
Event|Activity|Impression|8714,8724|false|false|false|C0599946|Attenuation|attenuated
Finding|Functional Concept|Impression|8725,8729|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Social Behavior|Impression|8733,8741|false|false|false|C0678975|inferiority|inferior
Drug|Chemical Viewed Structurally|Impression|8742,8748|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|Impression|8742,8748|false|false|false|||branch
Event|Event|Impression|8759,8767|false|false|false|||evidence
Finding|Idea or Concept|Impression|8759,8767|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|8759,8770|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Acquired Abnormality|Impression|8777,8786|true|false|false|C0001168|Complete obstruction|occlusion
Event|Event|Impression|8777,8786|false|false|false|||occlusion
Finding|Finding|Impression|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Impression|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Impression|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Impression|8777,8786|true|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Intellectual Product|Impression|8795,8800|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|8801,8813|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Impression|8801,8813|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|Impression|8814,8825|false|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Impression|8814,8825|false|false|false|||abnormality
Finding|Finding|Impression|8814,8825|false|false|false|C1704258|Abnormality|abnormality
Attribute|Clinical Attribute|Impression|8841,8848|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|Impression|8841,8848|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|Impression|8844,8848|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Impression|8844,8848|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Impression|8844,8848|false|false|false|C0362076|Problems with head|head
Event|Event|Impression|8844,8848|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Impression|8844,8848|false|false|false|C0876917|Procedure on head|head
Event|Event|Impression|8855,8858|false|false|false|||MRI
Finding|Gene or Genome|Impression|8855,8858|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Impression|8855,8858|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Impression|8855,8858|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Impression|8855,8863|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|Impression|8859,8863|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Impression|8859,8863|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Impression|8859,8863|false|false|false|C0362076|Problems with head|head
Event|Event|Impression|8859,8863|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Impression|8859,8863|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|8868,8876|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Impression|8868,8876|false|false|false|||contrast
Finding|Intellectual Product|Impression|8895,8900|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|Impression|8901,8913|false|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|Impression|8901,8913|false|false|false|C1522213|Intracranial Route of Administration|intracranial
Disorder|Congenital Abnormality|Impression|8914,8925|true|false|false|C0000768|Congenital Abnormality|abnormality
Event|Event|Impression|8914,8925|false|false|false|||abnormality
Finding|Finding|Impression|8914,8925|true|false|false|C1704258|Abnormality|abnormality
Event|Event|Impression|8945,8950|false|false|false|||large
Finding|Gene or Genome|Impression|8945,8950|true|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Event|Event|Impression|8962,8972|false|false|false|||infarction
Finding|Pathologic Function|Impression|8962,8972|false|false|false|C0021308|Infarction|infarction
Event|Event|Impression|8976,8986|false|false|false|||hemorrhage
Finding|Pathologic Function|Impression|8976,8986|false|false|false|C0019080|Hemorrhage|hemorrhage
Event|Event|Impression|9001,9005|false|false|false|||foci
Finding|Finding|Impression|9001,9005|false|false|false|C4321394|Foci|foci
Finding|Finding|Impression|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Impression|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Impression|9012,9016|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Phenomenon|Phenomenon or Process|Impression|9017,9023|false|false|false|C1710082|Signal|signal
Event|Event|Impression|9024,9033|false|false|false|||intensity
Anatomy|Body Location or Region|Impression|9041,9052|false|false|false|C0815275|Subcortical|subcortical
Anatomy|Body Part, Organ, or Organ Component|Impression|9058,9086|false|false|false|C0228157|Periventricular white matter|periventricular white matter
Anatomy|Tissue|Impression|9074,9086|false|false|false|C0682708|White matter|white matter
Event|Event|Impression|9091,9102|false|false|false|||nonspecific
Event|Event|Impression|9111,9118|false|false|false|||reflect
Event|Event|Impression|9120,9127|false|false|false|||changes
Finding|Functional Concept|Impression|9120,9127|false|false|false|C0392747|Changing|changes
Event|Event|Impression|9135,9142|false|false|false|||chronic
Finding|Intellectual Product|Impression|9135,9142|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Impression|9135,9142|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Anatomy|Body Part, Organ, or Organ Component|Impression|9143,9155|false|false|false|C0225988|Structure of small blood vessel (organ)|small vessel
Anatomy|Body Location or Region|Impression|9149,9155|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Impression|9149,9155|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Disorder|Disease or Syndrome|Impression|9156,9163|false|false|false|C0012634|Disease|disease
Event|Event|Impression|9156,9163|false|false|false|||disease
Event|Event|Impression|9170,9173|false|false|false|||TTE
Procedure|Diagnostic Procedure|Impression|9170,9173|false|false|false|C0430462|Transthoracic echocardiography|TTE
Event|Event|Impression|9174,9184|false|false|false|||IMPRESSION
Finding|Intellectual Product|Impression|9174,9184|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Impression|9174,9184|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Event|Event|Impression|9200,9206|false|false|false|||source
Finding|Finding|Impression|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Functional Concept|Impression|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Finding|Intellectual Product|Impression|9200,9206|true|false|false|C0449416;C1705919;C4521696|Source;Source (property) (qualifier value);Term Source|source
Event|Event|Impression|9210,9225|false|false|false|||thromboembolism
Finding|Pathologic Function|Impression|9210,9225|true|false|false|C0040038|Thromboembolism|thromboembolism
Event|Event|Impression|9226,9236|false|false|false|||identified
Finding|Finding|Impression|9250,9256|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|Impression|9250,9256|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|Impression|9257,9268|false|false|false|||predisposes
Finding|Pathologic Function|Impression|9272,9280|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|thrombus
Finding|Finding|Impression|9272,9290|false|false|false|C4717432|Thrombus formation|thrombus formation
Event|Event|Impression|9281,9290|false|false|false|||formation
Finding|Functional Concept|Impression|9281,9290|false|false|false|C1522492|Formation|formation
Phenomenon|Biologic Function|Impression|9281,9290|false|false|false|C0220781|Anabolism|formation
Finding|Functional Concept|Impression|9304,9308|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|9309,9320|false|false|false|C0018827|Heart Ventricle|ventricular
Finding|Organ or Tissue Function|Impression|9321,9329|false|false|false|C0039155|Systole|systolic
Event|Event|Impression|9330,9338|false|false|false|||function
Finding|Finding|Impression|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Functional Concept|Impression|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Intellectual Product|Impression|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Physiologic Function|Impression|9330,9338|false|true|false|C0031843;C0542341;C0598463;C1705273|Function (attribute);Functional Status;Mathematical Operator;physiological aspects|function
Finding|Mental Process|Impression|9346,9353|false|false|false|C0542559|contextual factors|setting
Event|Event|Impression|9358,9362|false|false|false|||beat
Event|Event|Impression|9371,9382|false|false|false|||variability
Finding|Conceptual Entity|Impression|9371,9382|false|false|false|C2827666|Variability|variability
Disorder|Disease or Syndrome|Impression|9390,9400|false|false|false|C0003811|Cardiac Arrhythmia|arrhythmia
Event|Event|Impression|9390,9400|false|false|false|||arrhythmia
Event|Event|Impression|9402,9406|false|false|false|||Mild
Finding|Intellectual Product|Impression|9402,9406|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Event|Event|Impression|9410,9418|false|false|false|||moderate
Finding|Finding|Impression|9410,9418|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Finding|Intellectual Product|Impression|9410,9418|false|false|false|C1547226;C5201148|Moderate;Moderate - Severity of Illness Code|moderate
Disorder|Disease or Syndrome|Impression|9431,9454|false|false|false|C0040961|Tricuspid Valve Insufficiency|tricuspid regurgitation
Event|Event|Impression|9441,9454|false|false|false|||regurgitation
Finding|Finding|Impression|9441,9454|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Finding|Sign or Symptom|Impression|9441,9454|false|false|false|C0232605;C2004489|Regurgitates after swallowing;Regurgitation|regurgitation
Phenomenon|Biologic Function|Impression|9441,9454|false|false|false|C0460152|Regurgitation - mechanism|regurgitation
Anatomy|Body Part, Organ, or Organ Component|Impression|9463,9472|false|false|false|C0024109|Lung|pulmonary
Attribute|Clinical Attribute|Impression|9463,9472|false|false|false|C2707265||pulmonary
Finding|Finding|Impression|9463,9472|false|false|false|C4522268|Pulmonary (intended site)|pulmonary
Event|Event|Impression|9473,9481|false|false|false|||pressure
Finding|Finding|Impression|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Impression|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Impression|9473,9481|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Impression|9473,9481|false|false|false|C0033095||pressure
Anatomy|Body Location or Region|Impression|9495,9506|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Anatomy|Body Part, Organ, or Organ Component|Impression|9495,9506|false|false|false|C0031050;C0442031|Pericardial (qualifier value);Pericardial sac structure|pericardial
Disorder|Disease or Syndrome|Impression|9495,9515|false|false|false|C0031039|Pericardial effusion|pericardial effusion
Finding|Body Substance|Impression|9495,9515|false|false|false|C1253937|Pericardial effusion body substance|pericardial effusion
Event|Event|Impression|9507,9515|false|false|false|||effusion
Finding|Body Substance|Impression|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Intellectual Product|Impression|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Pathologic Function|Impression|9507,9515|false|false|false|C0013687;C1546613;C2317432|Effusion (substance);effusion|effusion
Finding|Idea or Concept|Hospital Course|9558,9562|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Finding|Intellectual Product|Hospital Course|9558,9562|false|false|false|C1561543;C1561544|Precision - year;Transaction counts and value totals - year|year
Event|Event|Hospital Course|9563,9566|false|false|false|||old
Disorder|Disease or Syndrome|Hospital Course|9579,9583|false|false|false|C0004238|Atrial Fibrillation|AFib
Event|Event|Hospital Course|9579,9583|false|false|false|||AFib
Lab|Laboratory or Test Result|Hospital Course|9579,9583|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|AFib
Drug|Organic Chemical|Hospital Course|9587,9594|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|Hospital Course|9587,9594|false|false|false|C3530466|Eliquis|Eliquis
Event|Event|Hospital Course|9587,9594|false|false|false|||Eliquis
Anatomy|Body Space or Junction|Hospital Course|9596,9599|false|false|false|C0262212|Choroidal fissure|CHF
Disorder|Disease or Syndrome|Hospital Course|9596,9599|false|false|false|C0018802|Congestive heart failure|CHF
Event|Event|Hospital Course|9596,9599|false|false|false|||CHF
Event|Event|Hospital Course|9602,9605|false|false|false|||HLD
Disorder|Disease or Syndrome|Hospital Course|9607,9610|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Hospital Course|9607,9610|false|false|false|||HTN
Event|Event|Hospital Course|9615,9624|false|false|false|||presented
Finding|Intellectual Product|Hospital Course|9628,9640|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9641,9651|false|false|false|C0013362|Dysarthria|dysarthria
Event|Event|Hospital Course|9641,9651|false|false|false|||dysarthria
Finding|Finding|Hospital Course|9653,9661|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Finding|Idea or Concept|Hospital Course|9653,9661|false|false|false|C0205161;C1550458|Abnormal;Observation Interpretation - Abnormal|abnormal
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9662,9665|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|9662,9665|false|false|false|C3495676|Anorectal Malformations|arm
Event|Event|Hospital Course|9662,9665|false|false|false|||arm
Finding|Gene or Genome|Hospital Course|9662,9665|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9662,9665|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Event|Event|Hospital Course|9667,9676|false|false|false|||movements
Finding|Organism Function|Hospital Course|9667,9676|false|false|false|C0026649|Movement|movements
Finding|Intellectual Product|Hospital Course|9682,9686|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Finding|Hospital Course|9682,9694|false|false|false|C0234964|Poor balance (finding)|poor balance
Drug|Organic Chemical|Hospital Course|9687,9694|false|false|false|C4319618|Balance (substance)|balance
Drug|Pharmacologic Substance|Hospital Course|9687,9694|false|false|false|C4319618|Balance (substance)|balance
Event|Event|Hospital Course|9687,9694|false|false|false|||balance
Finding|Finding|Hospital Course|9687,9694|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Finding|Organism Function|Hospital Course|9687,9694|false|false|false|C0014653;C0560184|Ability to balance;Equilibrium|balance
Procedure|Diagnostic Procedure|Hospital Course|9687,9694|false|false|false|C2174421|examination of balance|balance
Event|Event|Hospital Course|9696,9702|false|false|false|||walker
Drug|Biomedical or Dental Material|Hospital Course|9706,9714|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|Hospital Course|9706,9714|false|false|false|||baseline
Finding|Idea or Concept|Hospital Course|9706,9714|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Intellectual Product|Hospital Course|9717,9722|false|false|false|C1697238|NIH stroke scale|NIHSS
Event|Event|Hospital Course|9730,9737|false|false|false|||slurred
Event|Event|Hospital Course|9738,9744|false|false|false|||speech
Finding|Organism Function|Hospital Course|9738,9744|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Hospital Course|9738,9744|false|false|false|C0846595|Speech assessment|speech
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9762,9765|false|false|false|C3813556|Cancer/Testis Antigen|CTA
Event|Event|Hospital Course|9762,9765|false|false|false|||CTA
Finding|Gene or Genome|Hospital Course|9762,9765|false|false|false|C3540513;C4554671|CERNA3 gene;PCYT1A wt Allele|CTA
Procedure|Diagnostic Procedure|Hospital Course|9762,9765|false|false|false|C3272310|Cardiac Computerized Tomographic Angiography|CTA
Anatomy|Body Location or Region|Hospital Course|9766,9770|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|9766,9770|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|9766,9770|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9766,9770|false|false|false|C0876917|Procedure on head|head
Anatomy|Body Location or Region|Hospital Course|9766,9779|false|false|false|C0460004|Head and neck structure|head and neck
Anatomy|Body Location or Region|Hospital Course|9775,9779|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Anatomy|Cell Component|Hospital Course|9775,9779|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|neck
Finding|Finding|Hospital Course|9775,9779|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|neck
Event|Event|Hospital Course|9784,9793|false|false|false|||completed
Event|Event|Hospital Course|9810,9817|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|9810,9817|false|false|false|C2699424|Concern|concern
Finding|Functional Concept|Hospital Course|9822,9826|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Drug|Chemical Viewed Structurally|Hospital Course|9830,9836|false|false|false|C1881507|Macromolecular Branch|branch
Event|Activity|Hospital Course|9837,9848|false|false|false|C0599946|Attenuation|attenuation
Event|Event|Hospital Course|9849,9859|false|false|false|||concerning
Event|Event|Hospital Course|9865,9873|false|false|false|||stenosis
Finding|Pathologic Function|Hospital Course|9865,9873|false|false|false|C1261287|Stenosis|stenosis
Disorder|Acquired Abnormality|Hospital Course|9877,9886|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|Hospital Course|9877,9886|false|false|false|||occlusion
Finding|Finding|Hospital Course|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Hospital Course|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Hospital Course|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Hospital Course|9877,9886|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Event|Event|Hospital Course|9913,9924|false|false|false|||transferred
Event|Event|Hospital Course|9930,9943|false|false|false|||consideration
Finding|Finding|Hospital Course|9930,9943|false|false|false|C0518609|Consideration|consideration
Event|Event|Hospital Course|9947,9959|false|false|false|||thrombectomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9947,9959|false|false|false|C0162578|Thrombectomy|thrombectomy
Finding|Intellectual Product|Hospital Course|9964,9969|false|false|false|C1697238|NIH stroke scale|NIHSS
Event|Activity|Hospital Course|9975,9982|false|false|false|C1706079||arrival
Event|Event|Hospital Course|9975,9982|false|false|false|||arrival
Finding|Functional Concept|Hospital Course|9975,9982|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|Hospital Course|9999,10005|false|false|false|||deemed
Event|Event|Hospital Course|10008,10017|false|false|false|||candidate
Finding|Conceptual Entity|Hospital Course|10008,10017|false|false|false|C4527371|Candidate|candidate
Event|Event|Hospital Course|10027,10035|false|false|false|||admitted
Disorder|Disease or Syndrome|Hospital Course|10054,10060|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|10054,10060|false|false|false|||stroke
Finding|Finding|Hospital Course|10054,10060|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Occupational Activity|Hospital Course|10061,10068|false|false|false|C0557854|Services|service
Finding|Idea or Concept|Hospital Course|10061,10068|false|false|false|C3245478|ActInformationPrivacyReason - service|service
Event|Event|Hospital Course|10081,10091|false|false|false|||evaluation
Finding|Idea or Concept|Hospital Course|10081,10091|false|false|false|C1550157|Processing type - Evaluation|evaluation
Procedure|Health Care Activity|Hospital Course|10081,10091|false|false|false|C0220825;C1261322|Evaluation;Evaluation procedure|evaluation
Finding|Finding|Hospital Course|10095,10103|false|false|false|C0332149|Possible|possible
Disorder|Disease or Syndrome|Hospital Course|10104,10107|false|true|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|Hospital Course|10104,10107|false|false|false|||TIA
Disorder|Disease or Syndrome|Hospital Course|10111,10117|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|10111,10117|false|false|false|||stroke
Finding|Finding|Hospital Course|10111,10117|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Hospital Course|10131,10139|false|false|false|||symptoms
Finding|Functional Concept|Hospital Course|10131,10139|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Hospital Course|10131,10139|true|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Hospital Course|10140,10145|false|false|false|||noted
Event|Event|Hospital Course|10153,10162|false|false|false|||admission
Procedure|Health Care Activity|Hospital Course|10153,10162|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|Hospital Course|10164,10167|false|false|false|||MRI
Finding|Gene or Genome|Hospital Course|10164,10167|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Hospital Course|10164,10167|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Hospital Course|10164,10167|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Diagnostic Procedure|Hospital Course|10164,10172|false|false|false|C0412674|MRI of head|MRI head
Anatomy|Body Location or Region|Hospital Course|10168,10172|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|10168,10172|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Hospital Course|10168,10172|false|false|false|C0362076|Problems with head|head
Event|Event|Hospital Course|10168,10172|false|false|false|||head
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10168,10172|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|10178,10186|false|false|false|C0009924|Contrast Media|contrast
Event|Event|Hospital Course|10178,10186|false|false|false|||contrast
Event|Event|Hospital Course|10200,10208|false|false|false|||evidence
Finding|Idea or Concept|Hospital Course|10200,10208|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|10200,10211|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Hospital Course|10212,10218|true|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|10212,10218|false|false|false|||stroke
Finding|Finding|Hospital Course|10212,10218|true|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Hospital Course|10220,10227|false|false|false|||Reports
Finding|Intellectual Product|Hospital Course|10220,10227|false|false|false|C0684224|Report (document)|Reports
Procedure|Health Care Activity|Hospital Course|10220,10227|false|false|false|C0700287|Reporting|Reports
Event|Event|Hospital Course|10236,10250|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|Hospital Course|10236,10250|false|false|false|C0013516|Echocardiography|echocardiogram
Finding|Classification|Hospital Course|10255,10265|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|10255,10265|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|Hospital Course|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|10266,10269|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|10266,10269|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|10266,10269|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|10266,10269|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|10266,10269|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Hospital Course|10284,10292|false|false|false|||reported
Finding|Intellectual Product|Hospital Course|10300,10305|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Attribute|Clinical Attribute|Hospital Course|10306,10314|false|false|false|C2926606||findings
Event|Event|Hospital Course|10306,10314|false|false|false|||findings
Finding|Functional Concept|Hospital Course|10306,10314|false|false|false|C2607943|findings aspects|findings
Event|Event|Hospital Course|10335,10343|false|false|false|||repeated
Event|Event|Hospital Course|10360,10367|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|10360,10367|false|false|false|C2699424|Concern|concern
Event|Event|Hospital Course|10384,10390|false|false|false|||memory
Finding|Finding|Hospital Course|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|Hospital Course|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|Hospital Course|10384,10390|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Event|Event|Hospital Course|10396,10400|false|false|false|||able
Finding|Finding|Hospital Course|10396,10400|false|false|false|C1299581|Able (qualifier value)|able
Event|Event|Hospital Course|10412,10416|false|false|false|||ADLs
Finding|Daily or Recreational Activity|Hospital Course|10412,10416|false|false|false|C0001288|Activity of daily living (function)|ADLs
Event|Event|Hospital Course|10421,10426|false|false|false|||meals
Finding|Daily or Recreational Activity|Hospital Course|10421,10426|false|false|false|C1998602|Meal (occasion for eating)|meals
Event|Event|Hospital Course|10436,10444|false|false|false|||provided
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10448,10451|false|false|false|C1431931|ALF protein, human|ALF
Drug|Biologically Active Substance|Hospital Course|10448,10451|false|false|false|C1431931|ALF protein, human|ALF
Event|Event|Hospital Course|10448,10451|false|false|false|||ALF
Finding|Gene or Genome|Hospital Course|10448,10451|false|false|false|C1332077;C1704942|GTF2A1L gene;GTF2A1L wt Allele|ALF
Event|Event|Hospital Course|10453,10458|false|false|false|||moved
Finding|Gene or Genome|Hospital Course|10469,10472|false|false|false|C1333533;C1704938|FBXW7 gene;FBXW7 wt Allele|ago
Event|Event|Hospital Course|10478,10485|false|false|false|||appears
Finding|Intellectual Product|Hospital Course|10505,10510|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|Hospital Course|10511,10517|false|false|false|||change
Finding|Functional Concept|Hospital Course|10511,10517|true|false|false|C0392747|Changing|change
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10511,10517|true|false|false|C4319952|Change - procedure|change
Event|Event|Hospital Course|10527,10533|false|false|false|||taking
Finding|Intellectual Product|Hospital Course|10550,10554|false|false|false|C1720092|Once - dosing instruction fragment|once
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10587,10590|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10587,10590|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10587,10590|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10587,10590|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10587,10590|false|false|false|C1332410|BID gene|BID
Drug|Pharmacologic Substance|Hospital Course|10591,10601|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Hospital Course|10591,10601|false|false|false|||medication
Finding|Intellectual Product|Hospital Course|10591,10601|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Event|Event|Hospital Course|10616,10620|false|false|false|||dose
Event|Event|Hospital Course|10625,10634|false|false|false|||increased
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10644,10647|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10644,10647|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10644,10647|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10644,10647|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10644,10647|false|false|false|C1332410|BID gene|BID
Event|Event|Hospital Course|10663,10672|false|false|false|||candidate
Finding|Conceptual Entity|Hospital Course|10663,10672|false|false|false|C4527371|Candidate|candidate
Disorder|Mental or Behavioral Dysfunction|Hospital Course|10682,10685|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10682,10685|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|10682,10685|false|false|false|C1530795|BID protein, human|BID
Event|Event|Hospital Course|10682,10685|false|false|false|||BID
Finding|Gene or Genome|Hospital Course|10682,10685|false|false|false|C1332410|BID gene|BID
Attribute|Clinical Attribute|Hospital Course|10697,10700|false|false|false|C1114365||age
Drug|Biologically Active Substance|Hospital Course|10697,10700|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Hospital Course|10697,10700|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Hospital Course|10697,10700|false|false|false|||age
Attribute|Clinical Attribute|Hospital Course|10705,10711|false|false|false|C0944911||weight
Event|Event|Hospital Course|10705,10711|false|false|false|||weight
Finding|Finding|Hospital Course|10705,10711|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Hospital Course|10705,10711|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Hospital Course|10705,10711|false|false|false|C1305866|Weighing patient|weight
Event|Event|Hospital Course|10722,10729|false|false|false|||started
Drug|Organic Chemical|Hospital Course|10733,10745|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|10733,10745|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|10733,10745|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|Hospital Course|10755,10769|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|hyperlipidemia
Event|Event|Hospital Course|10755,10769|false|false|false|||hyperlipidemia
Finding|Finding|Hospital Course|10755,10769|false|false|false|C0428465|Serum lipids high (finding)|hyperlipidemia
Drug|Biologically Active Substance|Hospital Course|10771,10774|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Hospital Course|10771,10774|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Hospital Course|10771,10774|false|false|false|||LDL
Procedure|Laboratory Procedure|Hospital Course|10771,10774|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Anatomy|Body System|Hospital Course|10784,10794|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Hospital Course|10799,10808|false|false|false|||consulted
Anatomy|Body Space or Junction|Hospital Course|10823,10828|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Hospital Course|10823,10828|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Hospital Course|10823,10828|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Hospital Course|10823,10828|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Attribute|Clinical Attribute|Hospital Course|10829,10835|false|false|false|C0488347||pauses
Event|Event|Hospital Course|10829,10835|false|false|false|||pauses
Event|Event|Hospital Course|10836,10841|false|false|false|||noted
Event|Event|Hospital Course|10845,10854|false|false|false|||telemetry
Procedure|Diagnostic Procedure|Hospital Course|10845,10854|false|false|false|C0039451|Telemetry|telemetry
Event|Event|Hospital Course|10860,10869|false|false|false|||persisted
Finding|Idea or Concept|Hospital Course|10887,10891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10887,10891|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10887,10891|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10892,10900|false|false|false|C0004147|atenolol|atenolol
Drug|Pharmacologic Substance|Hospital Course|10892,10900|false|false|false|C0004147|atenolol|atenolol
Event|Event|Hospital Course|10892,10900|false|false|false|||atenolol
Event|Event|Hospital Course|10902,10914|false|false|false|||recommending
Event|Event|Hospital Course|10929,10933|false|false|false|||home
Finding|Idea or Concept|Hospital Course|10929,10933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10929,10933|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10929,10933|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|10935,10942|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|Hospital Course|10935,10942|false|false|false|C0012265|digoxin|digoxin
Event|Event|Hospital Course|10935,10942|false|false|false|||digoxin
Procedure|Laboratory Procedure|Hospital Course|10935,10942|false|false|false|C0337449|Digoxin measurement|digoxin
Finding|Finding|Hospital Course|10947,10952|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|10947,10952|false|false|false|C0587267;C3810854|Close;Closed|close
Anatomy|Body System|Hospital Course|10953,10963|false|false|false|C0007226|Cardiovascular system|cardiology
Event|Event|Hospital Course|10969,10979|false|false|false|||Discharged
Event|Event|Hospital Course|10983,10987|false|false|false|||home
Finding|Idea or Concept|Hospital Course|10983,10987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10983,10987|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10983,10987|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|11006,11011|false|false|false|C0587267;C3810854|Close;Closed|close
Finding|Functional Concept|Hospital Course|11006,11011|false|false|false|C0587267;C3810854|Close;Closed|close
Disorder|Disease or Syndrome|Hospital Course|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Hospital Course|11012,11015|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Hospital Course|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Hospital Course|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Hospital Course|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Hospital Course|11012,11015|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Hospital Course|11012,11015|false|false|false|||PCP
Finding|Gene or Genome|Hospital Course|11012,11015|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Hospital Course|11012,11015|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Finding|Hospital Course|11023,11032|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|Transient
Event|Event|Hospital Course|11041,11047|false|false|false|||speech
Finding|Organism Function|Hospital Course|11041,11047|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Hospital Course|11041,11047|false|false|false|C0846595|Speech assessment|speech
Event|Event|Hospital Course|11052,11063|false|false|false|||instability
Finding|Finding|Hospital Course|11052,11063|false|false|false|C1444783|Instability|instability
Disorder|Disease or Syndrome|Hospital Course|11069,11072|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|Hospital Course|11069,11072|false|false|false|||TIA
Event|Event|Hospital Course|11079,11086|false|false|false|||consult
Procedure|Health Care Activity|Hospital Course|11079,11086|false|false|false|C0009818|Consultation|consult
Event|Event|Hospital Course|11089,11096|false|false|false|||cleared
Event|Event|Hospital Course|11101,11105|false|false|false|||home
Finding|Idea or Concept|Hospital Course|11101,11105|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11101,11105|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11101,11105|false|false|false|C1553498|home health encounter|home
Finding|Idea or Concept|Hospital Course|11111,11115|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11111,11115|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11111,11115|false|false|false|C1553498|home health encounter|home
Procedure|Health Care Activity|Hospital Course|11111,11124|false|false|false|C0020043|Home visit (procedure)|home services
Event|Event|Hospital Course|11116,11124|false|false|false|||services
Event|Occupational Activity|Hospital Course|11116,11124|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Hospital Course|11116,11124|false|false|false|C1704289|Clinical Service|services
Event|Event|Hospital Course|11127,11134|false|false|false|||Started
Drug|Organic Chemical|Hospital Course|11138,11150|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11138,11150|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Hospital Course|11138,11150|false|false|false|||atorvastatin
Event|Event|Hospital Course|11155,11158|false|false|false|||HLD
Finding|Idea or Concept|Hospital Course|11173,11177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|11173,11177|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|11173,11177|false|false|false|C1553498|home health encounter|home
Drug|Organic Chemical|Hospital Course|11178,11186|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Hospital Course|11178,11186|false|false|false|C1831808|apixaban|apixaban
Event|Event|Hospital Course|11178,11186|false|false|false|||apixaban
Drug|Organic Chemical|Hospital Course|11191,11202|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Hospital Course|11191,11202|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Finding|Functional Concept|Hospital Course|11191,11202|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Hospital Course|11191,11202|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11191,11202|false|false|false|C0087111|Therapeutic procedure|therapeutic
Disorder|Disease or Syndrome|Hospital Course|11220,11226|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|11220,11226|false|false|false|||stroke
Finding|Finding|Hospital Course|11220,11226|false|false|false|C5977286|Stroke (heart beat)|stroke
Event|Event|Hospital Course|11227,11236|false|false|false|||neurology
Event|Event|Hospital Course|11243,11252|false|false|false|||discharge
Finding|Body Substance|Hospital Course|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11243,11252|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11243,11252|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|11258,11264|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Hospital Course|11258,11264|false|false|false|||stroke
Finding|Finding|Hospital Course|11258,11264|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|Hospital Course|11258,11269|false|false|false|C1277291|Stroke risk|stroke risk
Finding|Idea or Concept|Hospital Course|11265,11269|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|Hospital Course|11265,11277|false|false|false|C1830376||risk factors
Finding|Finding|Hospital Course|11265,11277|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|Hospital Course|11265,11277|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|Hospital Course|11270,11277|false|false|false|||factors
Event|Event|Hospital Course|11308,11311|false|false|false|||A1c
Finding|Classification|Hospital Course|11308,11311|false|false|false|C4521595|United States Military enlisted E3 (qualifier value)|A1c
Procedure|Laboratory Procedure|Hospital Course|11308,11311|false|false|false|C0474680|Hemoglobin A1c measurement|A1c
Finding|Finding|Hospital Course|11320,11326|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Hospital Course|11320,11326|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Event|Event|Hospital Course|11327,11334|false|false|false|||chronic
Finding|Intellectual Product|Hospital Course|11327,11334|false|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|Hospital Course|11327,11334|false|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Functional Concept|Hospital Course|11345,11349|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11345,11366|false|false|false|C0226231|Structure of left vertebral artery|left vertebral artery
Finding|Pathologic Function|Hospital Course|11345,11376|false|false|false|C4536452|Occlusion of left vertebral artery (disorder)|left vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11350,11359|false|false|false|C0549207|Bone structure of spine|vertebral
Anatomy|Body Location or Region|Hospital Course|11350,11366|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11350,11366|false|false|false|C0042559;C4695118|Head+Neck>Vertebral artery;Structure of vertebral artery|vertebral artery
Finding|Pathologic Function|Hospital Course|11350,11376|false|false|false|C0265104|Vertebral artery obstruction (disorder)|vertebral artery occlusion
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|11360,11366|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|11360,11366|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Finding|Pathologic Function|Hospital Course|11360,11376|false|false|false|C0264995|Occlusion of artery (disorder)|artery occlusion
Disorder|Acquired Abnormality|Hospital Course|11367,11376|false|false|false|C0001168|Complete obstruction|occlusion
Event|Event|Hospital Course|11367,11376|false|false|false|||occlusion
Finding|Finding|Hospital Course|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Functional Concept|Hospital Course|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Organ or Tissue Function|Hospital Course|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Pathologic Function|Hospital Course|11367,11376|false|false|false|C0011382;C0028778;C0441597;C1110554;C1947917|Cardiovascular occlusion;Dental Occlusion;Obstruction;Occluded|occlusion
Finding|Finding|Hospital Course|11382,11390|false|false|false|C2984079|Somewhat|somewhat
Event|Activity|Hospital Course|11405,11415|false|false|false|C0599946|Attenuation|attenuated
Finding|Functional Concept|Hospital Course|11416,11420|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Social Behavior|Hospital Course|11424,11432|false|false|false|C0678975|inferiority|inferior
Drug|Chemical Viewed Structurally|Hospital Course|11433,11439|false|false|false|C1881507|Macromolecular Branch|branch
Event|Event|Hospital Course|11433,11439|false|false|false|||branch
Disorder|Disease or Syndrome|Hospital Course|11443,11457|false|false|false|C0020473;C0020476|Hyperlipidemia;Hyperlipoproteinemias|Hyperlipidemia
Event|Event|Hospital Course|11443,11457|false|false|false|||Hyperlipidemia
Finding|Finding|Hospital Course|11443,11457|false|false|false|C0428465|Serum lipids high (finding)|Hyperlipidemia
Drug|Biologically Active Substance|Hospital Course|11459,11462|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Hospital Course|11459,11462|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Hospital Course|11459,11462|false|false|false|||LDL
Procedure|Laboratory Procedure|Hospital Course|11459,11462|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Disorder|Disease or Syndrome|Hospital Course|11470,11477|false|false|false|C0028754|Obesity|Obesity
Event|Event|Hospital Course|11470,11477|false|false|false|||Obesity
Finding|Finding|Hospital Course|11470,11477|false|false|false|C4759928|BODY MASS INDEX QUANTITATIVE TRAIT LOCUS 20|Obesity
Event|Event|Hospital Course|11484,11491|false|false|false|||concern
Finding|Idea or Concept|Hospital Course|11484,11491|true|false|false|C2699424|Concern|concern
Event|Event|Hospital Course|11492,11497|false|false|false|||noted
Drug|Organic Chemical|Hospital Course|11502,11507|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Drug|Pharmacologic Substance|Hospital Course|11502,11507|false|false|false|C0723362|Sleep brand of diphenhydramine hydrochloride|sleep
Finding|Organism Function|Hospital Course|11502,11507|false|false|false|C0037313|Sleep|sleep
Disorder|Disease or Syndrome|Hospital Course|11502,11513|false|false|false|C0037315|Sleep Apnea Syndromes|sleep apnea
Event|Event|Hospital Course|11508,11513|false|false|false|||apnea
Finding|Sign or Symptom|Hospital Course|11508,11513|false|false|false|C0003578|Apnea|apnea
Event|Event|Hospital Course|11529,11534|false|false|false|||carry
Event|Event|Diagnosis|11553,11567|false|false|false|||echocardiogram
Procedure|Diagnostic Procedure|Diagnosis|11553,11567|false|false|false|C0013516|Echocardiography|echocardiogram
Event|Event|Diagnosis|11576,11580|false|false|false|||show
Event|Event|Diagnosis|11583,11586|false|false|false|||PFO
Event|Event|Diagnosis|11597,11602|false|false|false|||study
Finding|Intellectual Product|Diagnosis|11597,11602|false|false|false|C1705923|Study Object|study
Procedure|Research Activity|Diagnosis|11597,11602|false|false|false|C0008972;C0947630;C2603343|Clinical Research;Scientific Study;Study|study
Disorder|Disease or Syndrome|Diagnosis|11605,11608|false|false|false|C0002880;C0272325|Autoimmune hemolytic anemia;Factor 8 deficiency, acquired|AHA
Drug|Organic Chemical|Diagnosis|11605,11608|false|false|false|C0050451|acetohydroxamic acid|AHA
Drug|Pharmacologic Substance|Diagnosis|11605,11608|false|false|false|C0050451|acetohydroxamic acid|AHA
Event|Event|Diagnosis|11605,11608|false|false|false|||AHA
Drug|Amino Acid, Peptide, or Protein|Diagnosis|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Diagnosis|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Diagnosis|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Diagnosis|11609,11612|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Event|Event|Diagnosis|11609,11612|false|false|false|||ASA
Finding|Gene or Genome|Diagnosis|11609,11612|false|false|false|C1412553|ARSA gene|ASA
Anatomy|Cell Component|Diagnosis|11613,11617|false|false|false|C1167518|viral nucleocapsid location|Core
Finding|Body Substance|Diagnosis|11613,11617|false|false|false|C3274653|Core Specimen|Core
Event|Event|Diagnosis|11618,11626|false|false|false|||Measures
Finding|Functional Concept|Diagnosis|11618,11626|false|false|false|C1879489|Measures (attribute)|Measures
Finding|Functional Concept|Diagnosis|11631,11639|false|false|false|C0475224|Ischemic|Ischemic
Disorder|Disease or Syndrome|Diagnosis|11631,11646|false|false|false|C0948008|Ischemic stroke|Ischemic Stroke
Disorder|Disease or Syndrome|Diagnosis|11640,11646|false|false|false|C0038454|Cerebrovascular accident|Stroke
Event|Event|Diagnosis|11640,11646|false|false|false|||Stroke
Finding|Finding|Diagnosis|11640,11646|false|false|false|C5977286|Stroke (heart beat)|Stroke
Finding|Finding|Diagnosis|11651,11660|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|Transient
Finding|Functional Concept|Diagnosis|11661,11669|false|true|false|C0475224|Ischemic|Ischemic
Finding|Finding|Diagnosis|11671,11677|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|Attack
Finding|Social Behavior|Diagnosis|11671,11677|false|false|false|C1261512;C1304680|Attack (finding);Attack behavior|Attack
Disorder|Disease or Syndrome|Diagnosis|11681,11690|false|false|false|C0011168|Deglutition Disorders|Dysphagia
Procedure|Health Care Activity|Diagnosis|11681,11700|false|false|false|C0500456|Screening for dysphagia|Dysphagia screening
Event|Event|Diagnosis|11691,11700|false|false|false|||screening
Finding|Finding|Diagnosis|11691,11700|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|Diagnosis|11691,11700|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|Diagnosis|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|Diagnosis|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|Diagnosis|11691,11700|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Event|Event|Diagnosis|11715,11721|false|false|false|||intake
Finding|Functional Concept|Diagnosis|11715,11721|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|Diagnosis|11715,11721|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Finding|Diagnosis|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|11727,11730|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Diagnosis|11732,11741|false|false|false|||confirmed
Event|Event|Diagnosis|11757,11766|false|false|false|||confirmed
Anatomy|Body Location or Region|Diagnosis|11776,11779|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Diagnosis|11776,11779|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Diagnosis|11776,11779|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Event|Event|Diagnosis|11776,11779|false|false|false|||DVT
Procedure|Therapeutic or Preventive Procedure|Diagnosis|11776,11791|false|false|false|C0853245|DVT prophylaxis|DVT Prophylaxis
Event|Event|Diagnosis|11780,11791|false|false|false|||Prophylaxis
Procedure|Therapeutic or Preventive Procedure|Diagnosis|11780,11791|false|false|false|C0199176|Prophylactic treatment|Prophylaxis
Event|Event|Diagnosis|11792,11804|false|false|false|||administered
Finding|Finding|Diagnosis|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|11810,11813|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Diagnosis|11840,11847|false|false|false|||therapy
Finding|Finding|Diagnosis|11840,11847|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Diagnosis|11840,11847|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Diagnosis|11840,11847|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Diagnosis|11848,11860|false|false|false|||administered
Drug|Amino Acid, Peptide, or Protein|Diagnosis|11864,11867|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Diagnosis|11864,11867|false|false|false|C0082420|Endoglin, human|end
Event|Event|Diagnosis|11864,11867|false|false|false|||end
Finding|Functional Concept|Diagnosis|11864,11867|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Diagnosis|11864,11867|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Idea or Concept|Diagnosis|11871,11879|false|false|false|C1547192|Organization unit type - Hospital|hospital
Finding|Idea or Concept|Diagnosis|11880,11883|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|Diagnosis|11880,11883|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Finding|Diagnosis|11880,11885|false|false|false|C3842676|Day 2|day 2
Finding|Finding|Diagnosis|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|11892,11895|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|Diagnosis|11907,11910|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|11907,11910|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|11907,11910|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|11907,11910|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Event|Event|Diagnosis|11911,11921|false|false|false|||documented
Finding|Finding|Diagnosis|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|11927,11930|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|Diagnosis|11932,11935|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|11932,11935|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|11932,11935|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|11932,11935|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Drug|Organic Chemical|Diagnosis|11964,11970|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Diagnosis|11964,11970|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|Diagnosis|11964,11970|false|false|false|C1414273|EEF1A2 gene|statin
Procedure|Therapeutic or Preventive Procedure|Diagnosis|11964,11978|false|false|false|C1278454|Administration of prophylactic statin|statin therapy
Event|Event|Diagnosis|11971,11978|false|false|false|||therapy
Finding|Finding|Diagnosis|11971,11978|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Diagnosis|11971,11978|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Diagnosis|11971,11978|false|false|false|C0087111|Therapeutic procedure|therapy
Event|Event|Diagnosis|11979,11991|false|false|false|||administered
Drug|Organic Chemical|Diagnosis|11994,12005|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Diagnosis|11994,12005|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|Diagnosis|12013,12024|false|false|false|C0074554|simvastatin|simvastatin
Drug|Pharmacologic Substance|Diagnosis|12013,12024|false|false|false|C0074554|simvastatin|simvastatin
Drug|Organic Chemical|Diagnosis|12046,12058|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Diagnosis|12046,12058|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Diagnosis|12059,12063|false|false|false|||40mg
Drug|Organic Chemical|Diagnosis|12075,12087|false|false|false|C0965129|rosuvastatin|rosuvastatin
Drug|Pharmacologic Substance|Diagnosis|12075,12087|false|false|false|C0965129|rosuvastatin|rosuvastatin
Event|Event|Diagnosis|12088,12092|false|false|false|||20mg
Drug|Biologically Active Substance|Diagnosis|12106,12109|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12106,12109|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12106,12109|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12106,12109|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Finding|Diagnosis|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|12121,12124|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|Diagnosis|12138,12141|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12138,12141|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12138,12141|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12138,12141|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Drug|Biologically Active Substance|Diagnosis|12145,12148|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12145,12148|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12145,12148|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12145,12148|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Event|Event|Diagnosis|12154,12160|false|false|false|||reason
Finding|Idea or Concept|Diagnosis|12154,12160|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Event|Event|Diagnosis|12165,12170|false|false|false|||given
Drug|Organic Chemical|Diagnosis|12176,12182|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|Diagnosis|12176,12182|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Finding|Gene or Genome|Diagnosis|12176,12182|false|false|false|C1414273|EEF1A2 gene|Statin
Drug|Pharmacologic Substance|Diagnosis|12183,12193|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Diagnosis|12183,12193|false|false|false|||medication
Finding|Intellectual Product|Diagnosis|12183,12193|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Pathologic Function|Diagnosis|12183,12201|false|false|false|C0013182|Drug Allergy|medication allergy
Event|Event|Diagnosis|12194,12201|false|false|false|||allergy
Finding|Finding|Diagnosis|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|Diagnosis|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|Diagnosis|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|Diagnosis|12194,12201|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Event|Event|Diagnosis|12212,12219|false|false|false|||reasons
Finding|Idea or Concept|Diagnosis|12212,12219|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Event|Event|Diagnosis|12220,12230|false|false|false|||documented
Attribute|Clinical Attribute|Diagnosis|12234,12243|false|false|false|C0804815||physician
Event|Event|Diagnosis|12253,12261|false|false|false|||practice
Finding|Intellectual Product|Diagnosis|12253,12261|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Finding|Mental Process|Diagnosis|12253,12261|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Attribute|Clinical Attribute|Diagnosis|12269,12278|false|false|false|C0804815||physician
Attribute|Clinical Attribute|Diagnosis|12284,12293|false|false|false|C0804815||physician
Event|Event|Diagnosis|12294,12297|false|false|false|||APN
Finding|Gene or Genome|Diagnosis|12294,12297|false|false|false|C2986617|ANPEP wt Allele|APN
Event|Event|Diagnosis|12305,12315|false|false|false|||pharmacist
Finding|Idea or Concept|Diagnosis|12305,12315|false|false|false|C1546966|Primary Observer's Qualification - Pharmacist|pharmacist
Drug|Biologically Active Substance|Diagnosis|12320,12323|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12320,12323|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12320,12323|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12320,12323|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Individual Behavior|Diagnosis|12349,12356|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Intellectual Product|Diagnosis|12349,12356|false|false|false|C0037369;C0453996;C1548578|Location characteristic ID - Smoking;Smoking;Tobacco smoking behavior|Smoking
Finding|Individual Behavior|Diagnosis|12349,12366|false|false|false|C0085134|Cessation of smoking|Smoking cessation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12349,12366|false|false|false|C1095963|Smoking cessation therapy|Smoking cessation
Event|Activity|Diagnosis|12357,12366|false|false|false|C1880019|Cessation|cessation
Event|Event|Diagnosis|12357,12366|false|false|false|||cessation
Event|Event|Diagnosis|12367,12377|false|false|false|||counseling
Finding|Finding|Diagnosis|12367,12377|false|false|false|C0740209;C2148587|Encounter due to counseling;duration of counseling|counseling
Procedure|Health Care Activity|Diagnosis|12367,12377|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12367,12377|false|false|false|C0010210;C0542296|Counseling;Counselling service|counseling
Finding|Finding|Diagnosis|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|12388,12391|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Diagnosis|12402,12408|false|false|false|||reason
Finding|Idea or Concept|Diagnosis|12402,12408|true|false|false|C0392360|Indication of (contextual qualifier)|reason
Event|Event|Diagnosis|12430,12436|false|false|false|||unable
Finding|Finding|Diagnosis|12430,12436|false|false|false|C1299582|Unable|unable
Event|Event|Diagnosis|12440,12451|false|false|false|||participate
Disorder|Disease or Syndrome|Diagnosis|12456,12462|false|false|false|C0038454|Cerebrovascular accident|Stroke
Event|Event|Diagnosis|12456,12462|false|false|false|||Stroke
Finding|Finding|Diagnosis|12456,12462|false|false|false|C5977286|Stroke (heart beat)|Stroke
Procedure|Educational Activity|Diagnosis|12456,12472|false|false|false|C4303794|Education about stroke|Stroke education
Event|Event|Diagnosis|12463,12472|false|false|false|||education
Finding|Classification|Diagnosis|12463,12472|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Finding|Finding|Diagnosis|12463,12472|false|false|false|C0013622;C0013658;C0424927|Details of education;Educational Status;Educational aspects|education
Procedure|Educational Activity|Diagnosis|12463,12472|false|false|false|C0013621;C0039401|Education (procedure);Knowledge acquisition|education
Finding|Idea or Concept|Diagnosis|12494,12498|false|false|false|C0035647|Risk|risk
Attribute|Clinical Attribute|Diagnosis|12494,12506|false|false|false|C1830376||risk factors
Finding|Finding|Diagnosis|12494,12506|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Finding|Intellectual Product|Diagnosis|12494,12506|false|false|false|C0035648;C0455624;C1553898|History of - risk factor;risk factors;risk factors - observation list|risk factors
Event|Event|Diagnosis|12499,12506|false|false|false|||factors
Event|Activity|Diagnosis|12516,12524|false|false|false|C1879547|activation [action]|activate
Finding|Functional Concept|Diagnosis|12516,12524|false|false|false|C1515877;C3853838|activate - Data Operation;activate biological process|activate
Drug|Hazardous or Poisonous Substance|Diagnosis|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Organic Chemical|Diagnosis|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Drug|Pharmacologic Substance|Diagnosis|12525,12528|false|false|false|C0015063|Ethyl Methanesulfonate|EMS
Event|Event|Diagnosis|12525,12528|false|false|false|||EMS
Finding|Gene or Genome|Diagnosis|12525,12528|false|false|false|C5203240|EMSLR gene|EMS
Procedure|Health Care Activity|Diagnosis|12525,12528|false|false|false|C0013961|Emergency Medical Services|EMS
Disorder|Disease or Syndrome|Diagnosis|12533,12539|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Diagnosis|12533,12539|false|false|false|||stroke
Finding|Finding|Diagnosis|12533,12539|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Diagnosis|12541,12547|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Diagnosis|12541,12547|false|false|false|||stroke
Finding|Finding|Diagnosis|12541,12547|false|false|false|C5977286|Stroke (heart beat)|stroke
Finding|Conceptual Entity|Diagnosis|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Finding|Idea or Concept|Diagnosis|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Finding|Intellectual Product|Diagnosis|12548,12555|false|false|false|C0871599;C1549021;C1578603;C1578605;C4553014|Cautionary Warning;System Alert;Warning - AcknowledgementDetailType;Warning - EquipmentAlertLevel;Warning - Error severity|warning
Event|Governmental or Regulatory Activity|Diagnosis|12548,12561|false|false|false|C0871598|warning signs|warning signs
Event|Event|Diagnosis|12556,12561|false|false|false|||signs
Finding|Finding|Diagnosis|12556,12561|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Diagnosis|12556,12561|false|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Sign or Symptom|Diagnosis|12556,12574|false|false|false|C0037088|Signs and Symptoms|signs and symptoms
Event|Event|Diagnosis|12566,12574|false|false|false|||symptoms
Finding|Functional Concept|Diagnosis|12566,12574|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Diagnosis|12566,12574|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Attribute|Clinical Attribute|Diagnosis|12588,12599|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Diagnosis|12588,12599|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Diagnosis|12588,12599|false|false|false|||medications
Finding|Intellectual Product|Diagnosis|12588,12599|false|false|false|C4284232|Medications|medications
Event|Event|Diagnosis|12601,12605|false|false|false|||need
Finding|Functional Concept|Diagnosis|12601,12605|false|false|false|C0686904|Patient need for (contextual qualifier)|need
Finding|Functional Concept|Diagnosis|12601,12609|false|false|false|C0686904|Patient need for (contextual qualifier)|need for
Event|Event|Diagnosis|12610,12618|false|false|false|||followup
Procedure|Health Care Activity|Diagnosis|12610,12618|false|false|false|C1522577|follow-up|followup
Finding|Finding|Diagnosis|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|12654,12657|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Activity|Diagnosis|12669,12679|false|false|false|C1516048|Assessed|Assessment
Event|Event|Diagnosis|12669,12679|false|false|false|||Assessment
Finding|Intellectual Product|Diagnosis|12669,12679|false|false|false|C0679207|Knowledge acquisition using a method of assessment|Assessment
Procedure|Diagnostic Procedure|Diagnosis|12669,12679|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|Assessment
Procedure|Health Care Activity|Diagnosis|12669,12679|false|false|false|C0028708;C0031809;C0220825;C0542573;C0549068;C0549070;C0549071;C0549072;C0549073;C0549074;C0549075;C0549076;C0549078;C0549079;C0549080;C1161151;C1261322;C2237115|Evaluation;Evaluation procedure;Nutrition Assessment;Personal care assessment;Physical Examination;assessment of cognitive functions|Assessment
Procedure|Diagnostic Procedure|Diagnosis|12669,12698|false|false|false|C0431070|Assessment for rehabilitation|Assessment for rehabilitation
Event|Event|Diagnosis|12684,12698|false|false|false|||rehabilitation
Finding|Finding|Diagnosis|12684,12698|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Finding|Functional Concept|Diagnosis|12684,12698|false|false|false|C0007237;C0034992|Encounter due to care involving use of rehabilitation procedures;Rehabilitation aspects|rehabilitation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12684,12698|false|false|false|C0034991|Rehabilitation therapy|rehabilitation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12702,12707|false|false|false|C0034991|Rehabilitation therapy|rehab
Event|Event|Diagnosis|12708,12716|false|false|false|||services
Event|Occupational Activity|Diagnosis|12708,12716|false|false|false|C0557854|Services|services
Procedure|Health Care Activity|Diagnosis|12708,12716|false|false|false|C1704289|Clinical Service|services
Event|Event|Diagnosis|12717,12727|false|false|false|||considered
Finding|Finding|Diagnosis|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|12734,12737|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Diagnosis|12749,12759|false|false|false|||Discharged
Drug|Organic Chemical|Diagnosis|12763,12769|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Diagnosis|12763,12769|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|Diagnosis|12763,12769|false|false|false|C1414273|EEF1A2 gene|statin
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12763,12777|false|false|false|C1278454|Administration of prophylactic statin|statin therapy
Event|Event|Diagnosis|12770,12777|false|false|false|||therapy
Finding|Finding|Diagnosis|12770,12777|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Diagnosis|12770,12777|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Diagnosis|12770,12777|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Diagnosis|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|12783,12786|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Drug|Biologically Active Substance|Diagnosis|12799,12802|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12799,12802|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12799,12802|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12799,12802|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Finding|Idea or Concept|Diagnosis|12809,12815|false|false|false|C0392360|Indication of (contextual qualifier)|reason
Drug|Organic Chemical|Diagnosis|12831,12837|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Drug|Pharmacologic Substance|Diagnosis|12831,12837|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|Statin
Finding|Gene or Genome|Diagnosis|12831,12837|false|false|false|C1414273|EEF1A2 gene|Statin
Drug|Pharmacologic Substance|Diagnosis|12838,12848|false|false|false|C0013227|Pharmaceutical Preparations|medication
Event|Event|Diagnosis|12838,12848|false|false|false|||medication
Finding|Intellectual Product|Diagnosis|12838,12848|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Finding|Pathologic Function|Diagnosis|12838,12856|false|false|false|C0013182|Drug Allergy|medication allergy
Event|Event|Diagnosis|12849,12856|false|false|false|||allergy
Finding|Finding|Diagnosis|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Idea or Concept|Diagnosis|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Pathologic Function|Diagnosis|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Finding|Physiologic Function|Diagnosis|12849,12856|false|false|false|C0020517;C0489531;C1314973;C1527304;C1547542;C3539909|Allergic Reaction;Allergic disposition;Allergy - Charge Type Reason;History of allergies;Hypersensitivity;Response to antigens|allergy
Event|Event|Diagnosis|12867,12874|false|false|false|||reasons
Finding|Idea or Concept|Diagnosis|12867,12874|false|false|false|C0392360|Indication of (contextual qualifier)|reasons
Event|Event|Diagnosis|12875,12885|false|false|false|||documented
Attribute|Clinical Attribute|Diagnosis|12889,12898|false|false|false|C0804815||physician
Event|Event|Diagnosis|12908,12916|false|false|false|||practice
Finding|Intellectual Product|Diagnosis|12908,12916|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Finding|Mental Process|Diagnosis|12908,12916|false|false|false|C0237607;C3245512|Experience (Practice);HL7PublishingSubSection - practice|practice
Attribute|Clinical Attribute|Diagnosis|12924,12933|false|false|false|C0804815||physician
Attribute|Clinical Attribute|Diagnosis|12939,12948|false|false|false|C0804815||physician
Event|Event|Diagnosis|12949,12952|false|false|false|||APN
Finding|Gene or Genome|Diagnosis|12949,12952|false|false|false|C2986617|ANPEP wt Allele|APN
Event|Event|Diagnosis|12960,12970|false|false|false|||pharmacist
Finding|Idea or Concept|Diagnosis|12960,12970|false|false|false|C1546966|Primary Observer's Qualification - Pharmacist|pharmacist
Drug|Biologically Active Substance|Diagnosis|12975,12978|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Drug|Organic Chemical|Diagnosis|12975,12978|false|false|false|C0023823|Low-Density Lipoproteins|LDL
Event|Event|Diagnosis|12975,12978|false|false|false|||LDL
Procedure|Laboratory Procedure|Diagnosis|12975,12978|false|false|false|C0202117|Low density lipoprotein cholesterol measurement|LDL
Event|Event|Diagnosis|13004,13014|false|false|false|||Discharged
Event|Event|Diagnosis|13033,13040|false|false|false|||therapy
Finding|Finding|Diagnosis|13033,13040|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Finding|Functional Concept|Diagnosis|13033,13040|false|false|false|C0039798;C1363945|Therapy Object (animal model);therapeutic aspects|therapy
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13033,13040|false|false|false|C0087111|Therapeutic procedure|therapy
Finding|Finding|Diagnosis|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|13046,13049|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|13051,13055|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Finding|Intellectual Product|Diagnosis|13051,13055|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|Type
Drug|Pharmacologic Substance|Diagnosis|13061,13073|false|false|false|C5214487|Antiplatelet|Antiplatelet
Event|Event|Diagnosis|13080,13095|false|false|false|||Anticoagulation
Finding|Finding|Diagnosis|13080,13095|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Finding|Physiologic Function|Diagnosis|13080,13095|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|Anticoagulation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13080,13095|false|false|false|C0003281|Anticoagulation Therapy|Anticoagulation
Event|Event|Diagnosis|13109,13119|false|false|false|||Discharged
Anatomy|Body Space or Junction|Diagnosis|13123,13127|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Diagnosis|13123,13127|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Diagnosis|13123,13127|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Diagnosis|13123,13127|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Diagnosis|13128,13143|false|false|false|||anticoagulation
Finding|Finding|Diagnosis|13128,13143|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Diagnosis|13128,13143|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13128,13143|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Event|Diagnosis|13148,13156|false|false|false|||patients
Anatomy|Body Part, Organ, or Organ Component|Diagnosis|13162,13168|false|false|false|C0018792|Heart Atrium|atrial
Disorder|Disease or Syndrome|Diagnosis|13170,13182|false|false|false|C0232197|Fibrillation|fibrillation
Event|Event|Diagnosis|13170,13182|false|false|false|||fibrillation
Event|Event|Diagnosis|13183,13190|false|false|false|||flutter
Finding|Pathologic Function|Diagnosis|13183,13190|false|false|false|C0016385|Cardiac Flutter|flutter
Finding|Finding|Diagnosis|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Gene or Genome|Diagnosis|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Idea or Concept|Diagnosis|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Finding|Intellectual Product|Diagnosis|13196,13199|false|false|false|C0919479;C1298907;C1546947;C1546969;C1548171;C1549060;C1549065;C1549443;C1549445;C1705108;C1710701;C5202962;C5399964|YES Portal;YES1 gene;YES1 wt Allele;Yes;Yes (indicator);Yes (qualifier value);Yes - Assignment of Benefits;Yes - Event Expected;Yes - Expanded yes/no indicator;Yes - Identity May Be Divulged;Yes - Notify Clergy Code;Yes - Release Information;Yes - Yes/no indicator|Yes
Event|Event|Diagnosis|13213,13214|false|false|false|||N
Finding|Functional Concept|Diagnosis|13219,13228|false|false|false|C1516691|Cognitive|Cognitive
Event|Event|Diagnosis|13229,13239|false|false|false|||complaints
Finding|Finding|Diagnosis|13229,13239|false|false|false|C5441521|Complaint (finding)|complaints
Event|Event|Diagnosis|13242,13245|false|false|false|||B12
Finding|Gene or Genome|Diagnosis|13242,13245|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Finding|Intellectual Product|Diagnosis|13252,13260|false|false|false|C3241998|one time|one time
Finding|Finding|Diagnosis|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Diagnosis|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Diagnosis|13256,13260|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Event|Event|Diagnosis|13264,13279|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13264,13279|false|false|false|C0242297|Dietary Supplementation|supplementation
Finding|Intellectual Product|Diagnosis|13281,13285|false|false|false|C1720594|Then - dosing instruction fragment|then
Event|Event|Diagnosis|13286,13291|false|false|false|||start
Anatomy|Body Space or Junction|Diagnosis|13292,13296|false|false|false|C0226896|Oral cavity|oral
Drug|Biomedical or Dental Material|Diagnosis|13292,13296|false|false|false|C1272919|Oral Dosage Form|oral
Finding|Finding|Diagnosis|13292,13296|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Finding|Functional Concept|Diagnosis|13292,13296|false|false|false|C1527415;C4521986|Oral (intended site);Oral Route of Administration|oral
Event|Event|Diagnosis|13297,13300|false|false|false|||B12
Finding|Gene or Genome|Diagnosis|13297,13300|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Event|Event|Diagnosis|13302,13317|false|false|false|||supplementation
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13302,13317|false|false|false|C0242297|Dietary Supplementation|supplementation
Finding|Functional Concept|Diagnosis|13320,13330|false|false|false|C0521023|treponemal|Treponemal
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Immunologic Factor|Diagnosis|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Drug|Pharmacologic Substance|Diagnosis|13331,13341|false|false|false|C0003241;C3495458|Antibodies;antibodies (medication)|antibodies
Event|Event|Diagnosis|13331,13341|false|false|false|||antibodies
Lab|Laboratory or Test Result|Diagnosis|13331,13350|false|false|false|C0855852|Antibody NOS negative|antibodies negative
Event|Event|Diagnosis|13342,13350|false|false|false|||negative
Finding|Classification|Diagnosis|13342,13350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Diagnosis|13342,13350|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Diagnosis|13342,13350|false|false|false|C5237010|Expression Negative|negative
Event|Event|Diagnosis|13353,13361|false|false|false|||consider
Finding|Idea or Concept|Diagnosis|13353,13361|false|false|false|C0750591|consider|consider
Finding|Functional Concept|Diagnosis|13362,13371|false|false|false|C1516691|Cognitive|cognitive
Event|Event|Diagnosis|13382,13390|false|false|false|||referral
Procedure|Health Care Activity|Diagnosis|13382,13390|false|false|false|C0034927|Patient referral|referral
Event|Event|Diagnosis|13394,13404|false|false|false|||outpatient
Finding|Classification|Diagnosis|13394,13404|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Diagnosis|13394,13404|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|Diagnosis|13409,13415|false|false|false|||memory
Finding|Finding|Diagnosis|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|Diagnosis|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|Diagnosis|13409,13415|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Event|Event|Diagnosis|13417,13429|false|false|false|||difficulties
Finding|Finding|Diagnosis|13417,13429|true|false|false|C1299586|Has difficulty doing (qualifier value)|difficulties
Event|Event|Diagnosis|13434,13445|false|false|false|||appreciated
Event|Activity|Diagnosis|13453,13464|false|false|false|C4321457|Examination|examination
Event|Event|Diagnosis|13453,13464|false|false|false|||examination
Procedure|Health Care Activity|Diagnosis|13453,13464|false|false|false|C0031809;C0582103|Medical Examination;Physical Examination|examination
Disorder|Disease or Syndrome|Diagnosis|13467,13471|false|false|false|C0004238|Atrial Fibrillation|Afib
Lab|Laboratory or Test Result|Diagnosis|13467,13471|false|false|false|C0344434|Atrial Fibrillation by ECG Finding|Afib
Anatomy|Body Space or Junction|Diagnosis|13482,13487|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|Diagnosis|13482,13487|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|Diagnosis|13482,13487|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|Diagnosis|13482,13487|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Attribute|Clinical Attribute|Diagnosis|13488,13494|false|false|false|C0488347||pauses
Event|Event|Diagnosis|13488,13494|false|false|false|||pauses
Drug|Organic Chemical|Diagnosis|13505,13512|false|false|false|C0012265|digoxin|digoxin
Drug|Pharmacologic Substance|Diagnosis|13505,13512|false|false|false|C0012265|digoxin|digoxin
Event|Event|Diagnosis|13505,13512|false|false|false|||digoxin
Procedure|Laboratory Procedure|Diagnosis|13505,13512|false|false|false|C0337449|Digoxin measurement|digoxin
Disorder|Disease or Syndrome|Diagnosis|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Diagnosis|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Diagnosis|13559,13562|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Diagnosis|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Diagnosis|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Diagnosis|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Diagnosis|13559,13562|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Diagnosis|13559,13562|false|false|false|||PCP
Finding|Gene or Genome|Diagnosis|13559,13562|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Diagnosis|13559,13562|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Event|Event|Diagnosis|13566,13575|false|false|false|||increased
Drug|Organic Chemical|Diagnosis|13591,13602|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Diagnosis|13591,13602|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Diagnosis|13591,13602|false|false|false|||therapeutic
Finding|Functional Concept|Diagnosis|13591,13602|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Diagnosis|13591,13602|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Diagnosis|13591,13602|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|Diagnosis|13603,13609|false|false|false|||dosing
Drug|Organic Chemical|Diagnosis|13613,13620|false|false|false|C3530466|Eliquis|Eliquis
Drug|Pharmacologic Substance|Diagnosis|13613,13620|false|false|false|C3530466|Eliquis|Eliquis
Disorder|Mental or Behavioral Dysfunction|Diagnosis|13629,13632|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13629,13632|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Diagnosis|13629,13632|false|false|false|C1530795|BID protein, human|BID
Event|Event|Diagnosis|13629,13632|false|false|false|||BID
Finding|Gene or Genome|Diagnosis|13629,13632|false|false|false|C1332410|BID gene|BID
Event|Event|Diagnosis|13642,13646|false|false|false|||dose
Attribute|Clinical Attribute|Diagnosis|13653,13656|false|false|false|C1114365||age
Drug|Biologically Active Substance|Diagnosis|13653,13656|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Diagnosis|13653,13656|false|false|false|C0162574|Glycation End Products, Advanced|age
Event|Event|Diagnosis|13653,13656|false|false|false|||age
Attribute|Clinical Attribute|Diagnosis|13661,13667|false|false|false|C0944911||weight
Event|Event|Diagnosis|13661,13667|false|false|false|||weight
Finding|Finding|Diagnosis|13661,13667|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Finding|Sign or Symptom|Diagnosis|13661,13667|false|false|false|C0424653;C2053618|Weight symptom (finding);infant weight for previous delivery (history)|weight
Procedure|Health Care Activity|Diagnosis|13661,13667|false|false|false|C1305866|Weighing patient|weight
Event|Event|Diagnosis|13684,13691|false|false|false|||started
Drug|Organic Chemical|Diagnosis|13692,13704|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Diagnosis|13692,13704|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Diagnosis|13692,13704|false|false|false|||atorvastatin
Disorder|Disease or Syndrome|Diagnosis|13707,13710|false|false|false|C0020538|Hypertensive disease|HTN
Event|Event|Diagnosis|13707,13710|false|false|false|||HTN
Event|Event|Diagnosis|13713,13721|false|false|false|||continue
Finding|Idea or Concept|Diagnosis|13713,13721|false|false|false|C0549178|Continuous|continue
Finding|Idea or Concept|Diagnosis|13722,13726|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Diagnosis|13722,13726|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Diagnosis|13722,13726|false|false|false|C1553498|home health encounter|home
Drug|Pharmacologic Substance|Diagnosis|13727,13744|false|false|false|C0003364|Antihypertensive Agents|antihypertensives
Event|Event|Diagnosis|13727,13744|false|false|false|||antihypertensives
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13756,13764|false|false|false|C0041199|Troponin|troponin
Drug|Biologically Active Substance|Diagnosis|13756,13764|false|false|false|C0041199|Troponin|troponin
Event|Event|Diagnosis|13756,13764|false|false|false|||troponin
Procedure|Laboratory Procedure|Diagnosis|13756,13764|false|false|false|C0523952|Troponin measurement|troponin
Finding|Conceptual Entity|Diagnosis|13766,13774|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|RESOLVED
Finding|Pathologic Function|Diagnosis|13766,13774|false|false|false|C1514893;C2699488|Resolution;physiologic resolution|RESOLVED
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13778,13786|false|false|false|C0041199|Troponin|Troponin
Drug|Biologically Active Substance|Diagnosis|13778,13786|false|false|false|C0041199|Troponin|Troponin
Event|Event|Diagnosis|13778,13786|false|false|false|||Troponin
Procedure|Laboratory Procedure|Diagnosis|13778,13786|false|false|false|C0523952|Troponin measurement|Troponin
Event|Event|Diagnosis|13787,13795|false|false|false|||elevated
Event|Event|Diagnosis|13804,13812|false|false|false|||negative
Finding|Classification|Diagnosis|13804,13812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Diagnosis|13804,13812|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Diagnosis|13804,13812|false|false|false|C5237010|Expression Negative|negative
Event|Event|Diagnosis|13816,13825|false|false|false|||admission
Procedure|Health Care Activity|Diagnosis|13816,13825|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|Diagnosis|13828,13840|false|false|false|C0586553|Raised TSH level|elevated TSH
Attribute|Clinical Attribute|Diagnosis|13837,13840|false|false|false|C2708739||TSH
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Drug|Hormone|Diagnosis|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Drug|Pharmacologic Substance|Diagnosis|13837,13840|false|false|false|C0040160|thyrotropin|TSH
Event|Event|Diagnosis|13837,13840|false|false|false|||TSH
Procedure|Laboratory Procedure|Diagnosis|13837,13840|false|false|false|C0202230|Thyroid stimulating hormone measurement|TSH
Event|Event|Diagnosis|13850,13857|false|false|false|||recheck
Disorder|Disease or Syndrome|Diagnosis|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Mental or Behavioral Dysfunction|Diagnosis|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Disorder|Neoplastic Process|Diagnosis|13869,13872|false|false|false|C0431128;C1535939;C2919094|PCP - Hallucinogen-Related Disorder;Papillary craniopharyngioma;Pneumocystis jiroveci pneumonia|PCP
Drug|Amino Acid, Peptide, or Protein|Diagnosis|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Enzyme|Diagnosis|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Hazardous or Poisonous Substance|Diagnosis|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Organic Chemical|Diagnosis|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Drug|Pharmacologic Substance|Diagnosis|13869,13872|false|false|false|C0030855;C0031381;C1700512|BMP1 protein, human;Pentachlorophenol;Phencyclidine|PCP
Event|Event|Diagnosis|13869,13872|false|false|false|||PCP
Finding|Gene or Genome|Diagnosis|13869,13872|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Finding|Molecular Function|Diagnosis|13869,13872|false|false|false|C1418873;C1422070;C1744653;C3896095;C5551061|BMP1 wt Allele;PGPEP1 gene;PRCP gene;obsolete serine-type Pro-X carboxypeptidase activity;peptidyl carrier protein activity|PCP
Attribute|Clinical Attribute|Diagnosis|13879,13890|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Diagnosis|13879,13890|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Diagnosis|13879,13890|false|false|false|||Medications
Finding|Intellectual Product|Diagnosis|13879,13890|false|false|false|C4284232|Medications|Medications
Finding|Finding|Diagnosis|13879,13903|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|Diagnosis|13894,13903|false|false|false|||Admission
Procedure|Health Care Activity|Diagnosis|13894,13903|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Diagnosis|13922,13932|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Diagnosis|13922,13932|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Diagnosis|13922,13937|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|Diagnosis|13933,13937|false|false|false|||list
Finding|Intellectual Product|Diagnosis|13933,13937|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|Diagnosis|13941,13949|false|false|false|||accurate
Drug|Organic Chemical|Diagnosis|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Diagnosis|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Diagnosis|13954,13962|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Diagnosis|13954,13962|false|false|false|||complete
Finding|Functional Concept|Diagnosis|13954,13962|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Diagnosis|13954,13962|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|Diagnosis|13967,13975|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|Diagnosis|13967,13975|false|false|false|C0004147|atenolol|Atenolol
Drug|Organic Chemical|Diagnosis|13995,14003|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Diagnosis|13995,14003|false|false|false|C1831808|apixaban|Apixaban
Drug|Organic Chemical|Diagnosis|14024,14032|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Diagnosis|14024,14032|false|false|false|C0126174|losartan|Losartan
Event|Event|Diagnosis|14024,14032|false|false|false|||Losartan
Drug|Organic Chemical|Diagnosis|14024,14042|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Diagnosis|14024,14042|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Diagnosis|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Diagnosis|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Diagnosis|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Diagnosis|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Diagnosis|14033,14042|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Diagnosis|14033,14042|false|false|false|||Potassium
Finding|Physiologic Function|Diagnosis|14033,14042|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Diagnosis|14033,14042|false|false|false|C0202194|Potassium measurement|Potassium
Drug|Organic Chemical|Diagnosis|14062,14069|false|false|false|C0012265|digoxin|Digoxin
Drug|Pharmacologic Substance|Diagnosis|14062,14069|false|false|false|C0012265|digoxin|Digoxin
Procedure|Laboratory Procedure|Diagnosis|14062,14069|false|false|false|C0337449|Digoxin measurement|Digoxin
Drug|Antibiotic|Diagnosis|14092,14104|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|Diagnosis|14092,14104|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Event|Event|Diagnosis|14124,14133|false|false|false|||Discharge
Finding|Body Substance|Diagnosis|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Diagnosis|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Diagnosis|14124,14133|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Diagnosis|14124,14133|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Diagnosis|14124,14145|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Diagnosis|14134,14145|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Diagnosis|14134,14145|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|Diagnosis|14134,14145|false|false|false|||Medications
Finding|Intellectual Product|Diagnosis|14134,14145|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Diagnosis|14151,14163|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Diagnosis|14151,14163|false|false|false|C0286651|atorvastatin|Atorvastatin
Event|Event|Diagnosis|14173,14176|false|false|false|||QPM
Event|Event|Diagnosis|14178,14180|false|false|false|||RX
Drug|Organic Chemical|Diagnosis|14182,14194|false|false|false|C0286651|atorvastatin|atorvastatin
Drug|Pharmacologic Substance|Diagnosis|14182,14194|false|false|false|C0286651|atorvastatin|atorvastatin
Event|Event|Diagnosis|14182,14194|false|false|false|||atorvastatin
Drug|Biomedical or Dental Material|Diagnosis|14203,14209|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Diagnosis|14213,14221|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Diagnosis|14216,14221|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Diagnosis|14216,14221|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Diagnosis|14222,14226|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|Diagnosis|14255,14261|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Diagnosis|14262,14269|false|false|false|||Refills
Finding|Idea or Concept|Diagnosis|14262,14269|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Diagnosis|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Pharmacologic Substance|Diagnosis|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Drug|Vitamin|Diagnosis|14278,14292|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|Cyanocobalamin
Event|Event|Diagnosis|14278,14292|false|false|false|||Cyanocobalamin
Event|Event|Diagnosis|14297,14300|false|false|false|||mcg
Drug|Organic Chemical|Diagnosis|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Pharmacologic Substance|Diagnosis|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Drug|Vitamin|Diagnosis|14315,14329|false|false|false|C0042845;C3714801|Cyanocobalamin Drug Class;vitamin B12|cyanocobalamin
Event|Event|Diagnosis|14315,14329|false|false|false|||cyanocobalamin
Procedure|Laboratory Procedure|Diagnosis|14315,14344|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|cyanocobalamin (vitamin B-12)
Drug|Organic Chemical|Diagnosis|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Drug|Pharmacologic Substance|Diagnosis|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Drug|Vitamin|Diagnosis|14331,14338|false|false|false|C0042890|Vitamins|vitamin
Event|Event|Diagnosis|14331,14338|false|false|false|||vitamin
Drug|Organic Chemical|Diagnosis|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Pharmacologic Substance|Diagnosis|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Vitamin|Diagnosis|14331,14340|false|false|false|C0042849;C1704763;C5442122|B Vitamin Family;VITAMIN B;vitamin B complex|vitamin B
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Diagnosis|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Organic Chemical|Diagnosis|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Pharmacologic Substance|Diagnosis|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Drug|Vitamin|Diagnosis|14331,14343|false|false|false|C0042845;C0086024|cobalamins;vitamin B12|vitamin B-12
Procedure|Laboratory Procedure|Diagnosis|14331,14343|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|vitamin B-12
Drug|Biomedical or Dental Material|Diagnosis|14355,14361|false|false|false|C0039225|Tablet Dosage Form|tablet
Finding|Functional Concept|Diagnosis|14365,14373|false|false|false|C1527415|Oral Route of Administration|by mouth
Anatomy|Body Location or Region|Diagnosis|14368,14373|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Diagnosis|14368,14373|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Finding|Intellectual Product|Diagnosis|14375,14379|false|false|false|C1720092|Once - dosing instruction fragment|once
Drug|Biomedical or Dental Material|Diagnosis|14396,14402|false|false|false|C0039225|Tablet Dosage Form|Tablet
Event|Event|Diagnosis|14403,14410|false|false|false|||Refills
Finding|Idea or Concept|Diagnosis|14403,14410|false|false|false|C0807726|refill|Refills
Drug|Organic Chemical|Diagnosis|14419,14427|false|false|false|C1831808|apixaban|Apixaban
Drug|Pharmacologic Substance|Diagnosis|14419,14427|false|false|false|C1831808|apixaban|Apixaban
Disorder|Mental or Behavioral Dysfunction|Diagnosis|14438,14441|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Diagnosis|14438,14441|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Diagnosis|14438,14441|false|false|false|C1530795|BID protein, human|BID
Event|Event|Diagnosis|14438,14441|false|false|false|||BID
Finding|Gene or Genome|Diagnosis|14438,14441|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Diagnosis|14448,14456|false|false|false|C0004147|atenolol|Atenolol
Drug|Pharmacologic Substance|Diagnosis|14448,14456|false|false|false|C0004147|atenolol|Atenolol
Drug|Antibiotic|Diagnosis|14478,14490|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|Diagnosis|14478,14490|false|false|false|C0282386|levofloxacin|LevoFLOXacin
Drug|Organic Chemical|Diagnosis|14512,14520|false|false|false|C0126174|losartan|Losartan
Drug|Pharmacologic Substance|Diagnosis|14512,14520|false|false|false|C0126174|losartan|Losartan
Event|Event|Diagnosis|14512,14520|false|false|false|||Losartan
Drug|Organic Chemical|Diagnosis|14512,14530|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Pharmacologic Substance|Diagnosis|14512,14530|false|false|false|C0700492|losartan potassium|Losartan Potassium
Drug|Biologically Active Substance|Diagnosis|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Element, Ion, or Isotope|Diagnosis|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Food|Diagnosis|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Inorganic Chemical|Diagnosis|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Drug|Pharmacologic Substance|Diagnosis|14521,14530|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|Potassium
Event|Event|Diagnosis|14521,14530|false|false|false|||Potassium
Finding|Physiologic Function|Diagnosis|14521,14530|false|false|false|C4553027|Potassium metabolic function|Potassium
Procedure|Laboratory Procedure|Diagnosis|14521,14530|false|false|false|C0202194|Potassium measurement|Potassium
Event|Event|Diagnosis|14551,14560|false|false|false|||Discharge
Finding|Body Substance|Diagnosis|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Diagnosis|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Diagnosis|14551,14560|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Diagnosis|14551,14560|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Diagnosis|14551,14572|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Diagnosis|14551,14572|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Diagnosis|14561,14572|false|false|false|C2926604||Disposition
Event|Event|Diagnosis|14561,14572|false|false|false|||Disposition
Procedure|Health Care Activity|Diagnosis|14561,14572|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|Diagnosis|14574,14578|false|false|false|||Home
Finding|Idea or Concept|Diagnosis|14574,14578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Diagnosis|14574,14578|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Diagnosis|14574,14578|false|false|false|C1553498|home health encounter|Home
Event|Occupational Activity|Diagnosis|14584,14591|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|Diagnosis|14584,14591|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Event|Event|Diagnosis|14594,14602|false|false|false|||Facility
Finding|Intellectual Product|Diagnosis|14594,14602|false|false|false|C4695111|ADMIN.FACILITY|Facility
Event|Event|Diagnosis|14610,14619|false|false|false|||Discharge
Finding|Body Substance|Diagnosis|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Diagnosis|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Diagnosis|14610,14619|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Diagnosis|14610,14619|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Diagnosis|14610,14629|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Diagnosis|14620,14629|false|false|false|C0945731||Diagnosis
Event|Event|Diagnosis|14620,14629|false|false|false|||Diagnosis
Finding|Classification|Diagnosis|14620,14629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Diagnosis|14620,14629|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Diagnosis|14620,14629|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|Diagnosis|14631,14640|false|false|false|C0687129;C1550450|Encounter due to vagabond status;Living Arrangement - Transient|transient
Disorder|Mental or Behavioral Dysfunction|Diagnosis|14641,14651|false|false|false|C0013362|Dysarthria|dysarthria
Event|Event|Diagnosis|14641,14651|false|false|false|||dysarthria
Disorder|Neoplastic Process|Diagnosis|14656,14665|true|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|Diagnosis|14656,14665|false|false|false|||secondary
Finding|Functional Concept|Diagnosis|14656,14665|true|false|false|C1522484|metastatic qualifier|secondary
Disorder|Disease or Syndrome|Diagnosis|14669,14672|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|Diagnosis|14669,14672|false|false|false|||TIA
Disorder|Disease or Syndrome|Diagnosis|14676,14682|false|true|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Diagnosis|14676,14682|false|false|false|||stroke
Finding|Finding|Diagnosis|14676,14682|false|true|false|C5977286|Stroke (heart beat)|stroke
Finding|Intellectual Product|Diagnosis|14683,14687|false|false|false|C1547225|Mild Severity of Illness Code|Mild
Drug|Organic Chemical|Diagnosis|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Diagnosis|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Diagnosis|14688,14695|false|false|false|C0042890|Vitamins|Vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Diagnosis|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Organic Chemical|Diagnosis|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Pharmacologic Substance|Diagnosis|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Vitamin|Diagnosis|14688,14699|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Procedure|Laboratory Procedure|Diagnosis|14688,14699|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|Vitamin B12
Disorder|Disease or Syndrome|Diagnosis|14688,14710|false|false|false|C0042847|Vitamin B 12 Deficiency|Vitamin B12 deficiency
Finding|Finding|Diagnosis|14688,14710|false|false|false|C5886863|Decreased circulating vitamin B12 concentration|Vitamin B12 deficiency
Finding|Gene or Genome|Diagnosis|14696,14699|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Disorder|Disease or Syndrome|Diagnosis|14700,14710|false|false|false|C0162429|Malnutrition|deficiency
Event|Event|Diagnosis|14700,14710|false|false|false|||deficiency
Finding|Functional Concept|Diagnosis|14700,14710|false|false|false|C0011155|Deficiency|deficiency
Finding|Mental Process|Discharge Condition|14734,14740|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|14734,14747|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|14734,14747|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|14741,14747|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|14741,14747|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|14749,14754|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|14749,14754|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|14759,14767|false|false|false|||coherent
Finding|Finding|Discharge Condition|14759,14767|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|14769,14774|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|14769,14791|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|14769,14791|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|14778,14791|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|14778,14791|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|14778,14791|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|14793,14798|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|14793,14798|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|14793,14798|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|14793,14798|false|false|false|||Alert
Finding|Finding|Discharge Condition|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|14793,14798|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|14803,14814|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|14803,14814|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|14816,14824|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|14816,14824|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|14816,14824|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|14825,14831|false|false|false|C5889824||Status
Event|Event|Discharge Condition|14825,14831|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|14825,14831|false|false|false|C1546481|What subject filter - Status|Status
Finding|Functional Concept|Discharge Condition|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|14833,14843|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|14833,14843|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|14846,14854|false|false|false|||requires
Event|Event|Discharge Condition|14855,14865|false|false|false|||assistance
Finding|Social Behavior|Discharge Condition|14855,14865|false|false|false|C0018896|Helping Behavior|assistance
Drug|Amino Acid, Peptide, or Protein|Discharge Condition|14869,14872|false|false|false|C1454018|AICDA protein, human|aid
Drug|Enzyme|Discharge Condition|14869,14872|false|false|false|C1454018|AICDA protein, human|aid
Event|Event|Discharge Condition|14869,14872|false|false|false|||aid
Finding|Gene or Genome|Discharge Condition|14869,14872|false|false|false|C1421876;C3540469|AICDA gene;AICDA wt Allele|aid
Procedure|Therapeutic or Preventive Procedure|Discharge Condition|14869,14872|false|false|false|C0021588;C0280108|AID - Artificial insemination by donor;dacarbazine/doxorubicin/ifosfamide protocol|aid
Event|Event|Discharge Condition|14874,14880|false|false|false|||walker
Finding|Gene or Genome|Discharge Instructions|14918,14922|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|14942,14954|false|false|false|||hospitalized
Event|Event|Discharge Instructions|14962,14970|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|14962,14970|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|14962,14970|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|14982,14988|false|false|false|||speech
Finding|Organism Function|Discharge Instructions|14982,14988|false|false|false|C0037817|Speech|speech
Procedure|Diagnostic Procedure|Discharge Instructions|14982,14988|false|false|false|C0846595|Speech assessment|speech
Event|Event|Discharge Instructions|14997,15004|false|false|false|||concern
Finding|Idea or Concept|Discharge Instructions|14997,15004|false|false|false|C2699424|Concern|concern
Finding|Intellectual Product|Discharge Instructions|15012,15017|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|ACUTE
Disorder|Disease or Syndrome|Discharge Instructions|15012,15033|false|false|false|C5392833|Acute Ischemic Stroke|ACUTE ISCHEMIC STROKE
Finding|Functional Concept|Discharge Instructions|15018,15026|false|false|false|C0475224|Ischemic|ISCHEMIC
Disorder|Disease or Syndrome|Discharge Instructions|15018,15033|false|false|false|C0948008|Ischemic stroke|ISCHEMIC STROKE
Disorder|Disease or Syndrome|Discharge Instructions|15027,15033|false|false|false|C0038454|Cerebrovascular accident|STROKE
Event|Event|Discharge Instructions|15027,15033|false|false|false|||STROKE
Finding|Finding|Discharge Instructions|15027,15033|false|false|false|C5977286|Stroke (heart beat)|STROKE
Attribute|Clinical Attribute|Discharge Instructions|15037,15046|false|false|false|C3864998||condition
Disorder|Disease or Syndrome|Discharge Instructions|15037,15046|false|false|false|C0012634|Disease|condition
Event|Event|Discharge Instructions|15037,15046|false|false|false|||condition
Finding|Conceptual Entity|Discharge Instructions|15037,15046|false|false|false|C1705253|Logical Condition|condition
Disorder|Disease or Syndrome|Discharge Instructions|15055,15060|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|15055,15060|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|15055,15060|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Anatomy|Body Location or Region|Discharge Instructions|15062,15068|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15062,15068|false|false|false|C0005847;C0042591|Blood Vessel;Vessel Positions|vessel
Event|Event|Discharge Instructions|15069,15078|false|false|false|||providing
Drug|Biologically Active Substance|Discharge Instructions|15079,15085|false|false|false|C0030054|oxygen|oxygen
Drug|Element, Ion, or Isotope|Discharge Instructions|15079,15085|false|false|false|C0030054|oxygen|oxygen
Drug|Pharmacologic Substance|Discharge Instructions|15079,15085|false|false|false|C0030054|oxygen|oxygen
Event|Event|Discharge Instructions|15079,15085|false|false|false|||oxygen
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|15079,15085|false|false|false|C0184633|Oxygen Therapy Care|oxygen
Drug|Food|Discharge Instructions|15090,15099|false|false|false|C0678695|Nutrients|nutrients
Event|Event|Discharge Instructions|15090,15099|false|false|false|||nutrients
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15107,15112|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|15107,15112|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|15116,15123|false|false|false|||blocked
Drug|Organic Chemical|Discharge Instructions|15130,15134|false|false|false|C0009074|clotrimazole|clot
Drug|Pharmacologic Substance|Discharge Instructions|15130,15134|false|false|false|C0009074|clotrimazole|clot
Event|Event|Discharge Instructions|15130,15134|false|false|false|||clot
Finding|Pathologic Function|Discharge Instructions|15130,15134|false|false|false|C0302148|Blood Clot|clot
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15140,15145|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|15140,15145|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|15153,15157|false|false|false|||part
Finding|Idea or Concept|Discharge Instructions|15153,15157|false|false|false|C1552020|Role Class - part|part
Anatomy|Anatomical Structure|Discharge Instructions|15166,15170|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15166,15170|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Discharge Instructions|15166,15170|false|false|false|C1551342|Document Body|body
Event|Event|Discharge Instructions|15190,15197|false|false|false|||directs
Event|Event|Discharge Instructions|15212,15217|false|false|false|||parts
Anatomy|Anatomical Structure|Discharge Instructions|15226,15230|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15226,15230|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Discharge Instructions|15226,15230|false|false|false|C1551342|Document Body|body
Disorder|Injury or Poisoning|Discharge Instructions|15235,15241|false|false|false|C0010957|Tissue damage|damage
Event|Event|Discharge Instructions|15235,15241|false|false|false|||damage
Finding|Functional Concept|Discharge Instructions|15235,15241|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Finding|Gene or Genome|Discharge Instructions|15235,15241|false|false|false|C1883709;C2681922|Damage;MAGEE1 gene|damage
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15249,15254|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|15249,15254|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|15267,15275|false|false|false|||deprived
Disorder|Disease or Syndrome|Discharge Instructions|15283,15288|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|15283,15288|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|15283,15288|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Organ or Tissue Function|Discharge Instructions|15283,15295|false|false|false|C0678861;C0920762|Arterial blood supply;Vascular blood supply|blood supply
Finding|Physiologic Function|Discharge Instructions|15283,15295|false|false|false|C0678861;C0920762|Arterial blood supply;Vascular blood supply|blood supply
Event|Activity|Discharge Instructions|15289,15295|false|false|false|C1999230|Providing (action)|supply
Event|Event|Discharge Instructions|15289,15295|false|false|false|||supply
Finding|Functional Concept|Discharge Instructions|15289,15295|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Finding|Idea or Concept|Discharge Instructions|15289,15295|false|false|false|C0243163;C1561604;C4760136|Supply (process);Supply (system);supply aspects|supply
Event|Event|Discharge Instructions|15300,15306|false|false|false|||result
Event|Event|Discharge Instructions|15312,15319|false|false|false|||variety
Finding|Conceptual Entity|Discharge Instructions|15312,15319|false|false|false|C1883525;C2346866|Assortment;Variety (taxon)|variety
Event|Event|Discharge Instructions|15324,15332|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|15324,15332|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|15324,15332|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|15347,15350|false|false|false|||MRI
Finding|Gene or Genome|Discharge Instructions|15347,15350|false|false|false|C1824234|CYREN gene|MRI
Procedure|Diagnostic Procedure|Discharge Instructions|15347,15350|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Procedure|Health Care Activity|Discharge Instructions|15347,15350|false|false|false|C0024485;C0587658|Magnetic Resonance Imaging;Magnetic resonance imaging service|MRI
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15359,15364|false|false|false|C0006104;C4266577|Brain;Head>Brain|brain
Disorder|Disease or Syndrome|Discharge Instructions|15359,15364|false|false|false|C0006111|Brain Diseases|brain
Event|Event|Discharge Instructions|15373,15377|false|false|false|||show
Event|Event|Discharge Instructions|15379,15387|false|false|false|||evidence
Finding|Idea or Concept|Discharge Instructions|15379,15387|false|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Discharge Instructions|15379,15390|false|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Disorder|Disease or Syndrome|Discharge Instructions|15391,15397|false|false|false|C0038454|Cerebrovascular accident|stroke
Event|Event|Discharge Instructions|15391,15397|false|false|false|||stroke
Finding|Finding|Discharge Instructions|15391,15397|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Discharge Instructions|15401,15404|false|false|false|C0007787;C0917805|Transient Cerebral Ischemia;Transient Ischemic Attack|TIA
Event|Event|Discharge Instructions|15401,15404|false|false|false|||TIA
Event|Event|Discharge Instructions|15411,15419|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|15411,15419|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|15411,15419|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Drug|Organic Chemical|Discharge Instructions|15436,15443|false|false|false|C0163712|Relate - vinyl resin|related
Event|Event|Discharge Instructions|15436,15443|false|false|false|||related
Finding|Finding|Discharge Instructions|15436,15443|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Discharge Instructions|15436,15443|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|Discharge Instructions|15448,15453|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|15448,15453|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|15448,15453|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|15448,15462|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|15448,15462|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|15448,15462|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Discharge Instructions|15454,15462|false|false|false|||pressure
Finding|Finding|Discharge Instructions|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|15454,15462|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|15454,15462|false|false|false|C0033095||pressure
Disorder|Disease or Syndrome|Discharge Instructions|15464,15475|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Disorder|Injury or Poisoning|Discharge Instructions|15464,15475|false|false|false|C0011175;C2062903|Dehydration;dehydration (Na, H2O)|dehydration
Event|Event|Discharge Instructions|15464,15475|false|false|false|||dehydration
Procedure|Laboratory Procedure|Discharge Instructions|15464,15475|false|false|false|C4284399|Dehydration procedure|dehydration
Drug|Organic Chemical|Discharge Instructions|15477,15484|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Drug|Pharmacologic Substance|Discharge Instructions|15477,15484|false|false|false|C0001962;C0001975|Alcohols;ethanol|alcohol
Finding|Intellectual Product|Discharge Instructions|15477,15484|false|false|false|C1547288|Alcohol - Recreational Drug Use Code|alcohol
Finding|Finding|Discharge Instructions|15477,15488|false|false|false|C0001948;C0552479|Alcohol consumption;history of alcohol use|alcohol use
Finding|Individual Behavior|Discharge Instructions|15477,15488|false|false|false|C0001948;C0552479|Alcohol consumption;history of alcohol use|alcohol use
Event|Event|Discharge Instructions|15485,15488|false|false|false|||use
Finding|Functional Concept|Discharge Instructions|15485,15488|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Finding|Intellectual Product|Discharge Instructions|15485,15488|false|false|false|C0042153;C0457083;C1947944|Usage;Use - dosing instruction imperative;utilization qualifier|use
Event|Event|Discharge Instructions|15495,15506|false|false|false|||combination
Finding|Finding|Discharge Instructions|15495,15506|false|false|false|C3811910|combination - answer to question|combination
Event|Event|Discharge Instructions|15517,15524|false|false|false|||factors
Event|Event|Discharge Instructions|15534,15542|false|false|false|||changing
Attribute|Clinical Attribute|Discharge Instructions|15548,15559|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|15548,15559|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|15548,15559|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|15548,15559|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|Discharge Instructions|15581,15589|false|false|false|C1831808|apixaban|apixaban
Drug|Pharmacologic Substance|Discharge Instructions|15581,15589|false|false|false|C1831808|apixaban|apixaban
Event|Event|Discharge Instructions|15581,15589|false|false|false|||apixaban
Drug|Organic Chemical|Discharge Instructions|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Discharge Instructions|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Discharge Instructions|15617,15624|false|false|false|C0042890|Vitamins|Vitamin
Drug|Nucleic Acid, Nucleoside, or Nucleotide|Discharge Instructions|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Organic Chemical|Discharge Instructions|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Pharmacologic Substance|Discharge Instructions|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Drug|Vitamin|Discharge Instructions|15617,15628|false|false|false|C0042845;C0086024;C2936883|Vitamin B12 [EPC];cobalamins;vitamin B12|Vitamin B12
Procedure|Laboratory Procedure|Discharge Instructions|15617,15628|false|false|false|C0202252|VITAMIN B12 MEASUREMENT|Vitamin B12
Event|Event|Discharge Instructions|15625,15628|false|false|false|||B12
Finding|Gene or Genome|Discharge Instructions|15625,15628|false|false|false|C1417635;C1420797;C3538796|NDUFB3 gene;TNFAIP1 gene;TNFAIP1 wt Allele|B12
Drug|Food|Discharge Instructions|15635,15645|false|false|false|C0242295|Dietary Supplements|supplement
Event|Event|Discharge Instructions|15635,15645|false|false|false|||supplement
Finding|Functional Concept|Discharge Instructions|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Idea or Concept|Discharge Instructions|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Finding|Intellectual Product|Discharge Instructions|15635,15645|false|false|false|C1549514;C1947943;C2348609|Supplement;Supplement (document);Supplement - Diet Code Specification Type|supplement
Event|Event|Discharge Instructions|15654,15658|false|false|false|||take
Attribute|Clinical Attribute|Discharge Instructions|15670,15681|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|15670,15681|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|Discharge Instructions|15670,15681|false|false|false|||medications
Finding|Intellectual Product|Discharge Instructions|15670,15681|false|false|false|C4284232|Medications|medications
Event|Event|Discharge Instructions|15685,15695|false|false|false|||prescribed
Event|Event|Discharge Instructions|15705,15711|false|false|false|||follow
Finding|Intellectual Product|Discharge Instructions|15725,15737|false|false|false|C1547426|Location Service Code - Primary Care|primary care
Procedure|Health Care Activity|Discharge Instructions|15725,15737|false|false|false|C0033137|Primary Health Care|primary care
Event|Activity|Discharge Instructions|15733,15737|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|15733,15737|false|false|false|||care
Finding|Finding|Discharge Instructions|15733,15737|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|15733,15737|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Attribute|Clinical Attribute|Discharge Instructions|15738,15747|false|false|false|C0804815||physician
Event|Event|Discharge Instructions|15751,15757|false|false|false|||listed
Event|Event|Discharge Instructions|15782,15788|false|false|false|||follow
Event|Event|Discharge Instructions|15802,15814|false|false|false|||cardiologist
Event|Event|Discharge Instructions|15828,15833|false|false|false|||noted
Attribute|Clinical Attribute|Discharge Instructions|15853,15859|false|false|false|C0488347||pauses
Event|Event|Discharge Instructions|15853,15859|false|false|false|||pauses
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|15863,15870|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Discharge Instructions|15863,15870|false|false|false|C1314974|Cardiac attachment|cardiac
Procedure|Diagnostic Procedure|Discharge Instructions|15863,15881|false|false|false|C0150496|Cardiac monitoring|cardiac monitoring
Event|Activity|Discharge Instructions|15871,15881|false|false|false|C1283169||monitoring
Event|Event|Discharge Instructions|15871,15881|false|false|false|||monitoring
Procedure|Health Care Activity|Discharge Instructions|15871,15881|false|false|false|C0150369|Preventive monitoring|monitoring
Event|Event|Discharge Instructions|15891,15901|false|false|false|||experience
Event|Event|Discharge Instructions|15913,15921|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|15913,15921|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|15913,15921|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|15936,15940|false|false|false|||seek
Event|Event|Discharge Instructions|15942,15951|false|false|false|||emergency
Finding|Finding|Discharge Instructions|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Idea or Concept|Discharge Instructions|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Intellectual Product|Discharge Instructions|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Finding|Pathologic Function|Discharge Instructions|15942,15951|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|15942,15951|false|false|false|C0013956|Emergency Situation|emergency
Procedure|Health Care Activity|Discharge Instructions|15942,15951|false|false|false|C1553500|emergency encounter|emergency
Finding|Functional Concept|Discharge Instructions|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Idea or Concept|Discharge Instructions|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Finding|Intellectual Product|Discharge Instructions|15952,15959|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|medical
Procedure|Health Care Activity|Discharge Instructions|15952,15959|false|false|false|C0199168|Medical service|medical
Event|Event|Discharge Instructions|15960,15969|false|false|false|||attention
Finding|Intellectual Product|Discharge Instructions|15960,15969|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Discharge Instructions|15960,15969|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Event|Event|Discharge Instructions|15981,15990|false|false|false|||Emergency
Finding|Finding|Discharge Instructions|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Idea or Concept|Discharge Instructions|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Intellectual Product|Discharge Instructions|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Finding|Pathologic Function|Discharge Instructions|15981,15990|false|false|false|C1546399;C1546844;C1561583;C1561584;C1561585;C1561586;C1561587;C1561588;C1561589;C2745965|Admission Type - Emergency;Certification patient type - Emergency;Consent Bypass Reason - Emergency;Consent Non-Disclosure Reason - Emergency;Emergencies [Disease/Finding];Encounter Admission Source - emergency;Level of Care - Emergency;Patient Class - Emergency;Referral category - Emergency;Visit Priority Code - Emergency|Emergency
Phenomenon|Phenomenon or Process|Discharge Instructions|15981,15990|false|false|false|C0013956|Emergency Situation|Emergency
Procedure|Health Care Activity|Discharge Instructions|15981,15990|false|false|false|C1553500|emergency encounter|Emergency
Finding|Functional Concept|Discharge Instructions|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Idea or Concept|Discharge Instructions|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Finding|Intellectual Product|Discharge Instructions|15991,15998|false|false|false|C0205476;C1547184;C1561579|Medical;Medical referral type;Medical school type|Medical
Procedure|Health Care Activity|Discharge Instructions|15991,15998|false|false|false|C0199168|Medical service|Medical
Event|Event|Discharge Instructions|16000,16008|false|false|false|||Services
Event|Occupational Activity|Discharge Instructions|16000,16008|false|false|false|C0557854|Services|Services
Procedure|Health Care Activity|Discharge Instructions|16000,16008|false|false|false|C1704289|Clinical Service|Services
Event|Event|Discharge Instructions|16050,16059|false|false|false|||attention
Finding|Intellectual Product|Discharge Instructions|16050,16059|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Mental Process|Discharge Instructions|16050,16059|false|false|false|C0004268;C4281780|Attention;Attention - G-code|attention
Finding|Intellectual Product|Discharge Instructions|16068,16080|false|false|false|C1272517|Sudden onset (contextual qualifier) (qualifier value)|sudden onset
Event|Event|Discharge Instructions|16075,16080|false|false|false|||onset
Event|Event|Discharge Instructions|16085,16096|false|false|false|||persistence
Finding|Mental Process|Discharge Instructions|16085,16096|false|false|false|C0546816|Persistence|persistence
Event|Event|Discharge Instructions|16106,16114|false|false|false|||symptoms
Finding|Functional Concept|Discharge Instructions|16106,16114|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Finding|Sign or Symptom|Discharge Instructions|16106,16114|false|false|false|C0683368;C1457887|Symptoms;Symptoms aspect|symptoms
Event|Event|Discharge Instructions|16125,16132|false|false|false|||partial
Finding|Idea or Concept|Discharge Instructions|16125,16132|false|false|false|C1550516|Target Awareness - partial|partial
Drug|Organic Chemical|Discharge Instructions|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Discharge Instructions|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Discharge Instructions|16136,16144|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|Discharge Instructions|16136,16144|false|false|false|||complete
Finding|Functional Concept|Discharge Instructions|16136,16144|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Discharge Instructions|16136,16144|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Event|Event|Discharge Instructions|16145,16149|false|false|false|||loss
Finding|Finding|Discharge Instructions|16145,16149|false|false|false|C5890125|Loss (adaptation)|loss
Disorder|Disease or Syndrome|Discharge Instructions|16145,16159|false|false|false|C0042798;C0456909|Blindness;Low Vision|loss of vision
Finding|Finding|Discharge Instructions|16145,16159|false|false|false|C3665346;C3665386|Abnormal vision;Unspecified visual loss|loss of vision
Finding|Sign or Symptom|Discharge Instructions|16145,16159|false|false|false|C3665346;C3665386|Abnormal vision;Unspecified visual loss|loss of vision
Attribute|Clinical Attribute|Discharge Instructions|16153,16159|false|false|false|C2707266||vision
Event|Event|Discharge Instructions|16153,16159|false|false|false|||vision
Finding|Organism Function|Discharge Instructions|16153,16159|false|false|false|C0042789|Vision|vision
Event|Event|Discharge Instructions|16169,16173|false|false|false|||loss
Finding|Finding|Discharge Instructions|16169,16173|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|Discharge Instructions|16181,16188|false|false|false|||ability
Finding|Functional Concept|Discharge Instructions|16181,16188|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|Discharge Instructions|16181,16191|false|false|false|C5420000|Ability Question|ability to
Event|Event|Discharge Instructions|16198,16203|false|false|false|||words
Anatomy|Body Location or Region|Discharge Instructions|16214,16219|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Anatomy|Body Space or Junction|Discharge Instructions|16214,16219|false|false|false|C0226896;C0230028|Oral cavity;Oral region|mouth
Event|Event|Discharge Instructions|16229,16233|false|false|false|||loss
Finding|Finding|Discharge Instructions|16229,16233|false|false|false|C5890125|Loss (adaptation)|loss
Event|Event|Discharge Instructions|16241,16248|false|false|false|||ability
Finding|Functional Concept|Discharge Instructions|16241,16248|false|false|false|C5891046|Oral Intake Ability|ability
Finding|Intellectual Product|Discharge Instructions|16241,16251|false|false|false|C5420000|Ability Question|ability to
Event|Event|Discharge Instructions|16252,16262|false|false|false|||understand
Event|Event|Discharge Instructions|16270,16278|false|false|false|||speaking
Event|Event|Discharge Instructions|16296,16304|false|false|false|||weakness
Finding|Sign or Symptom|Discharge Instructions|16296,16304|false|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Anatomy|Anatomical Structure|Discharge Instructions|16324,16328|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16324,16328|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Discharge Instructions|16324,16328|false|false|false|C1551342|Document Body|body
Event|Event|Discharge Instructions|16338,16346|false|false|false|||drooping
Anatomy|Body Location or Region|Discharge Instructions|16366,16370|false|false|false|C0015450;C4266571|Face;Head>Face|face
Disorder|Disease or Syndrome|Discharge Instructions|16366,16370|false|false|false|C3160739|FANCONI ANEMIA, COMPLEMENTATION GROUP E|face
Event|Event|Discharge Instructions|16366,16370|false|false|false|||face
Finding|Gene or Genome|Discharge Instructions|16366,16370|false|false|false|C1414531;C1423759;C2828055|ELOVL6 gene;FANCE gene;FANCE wt Allele|face
Event|Event|Discharge Instructions|16380,16384|false|false|false|||loss
Finding|Finding|Discharge Instructions|16380,16384|false|false|false|C5890125|Loss (adaptation)|loss
Finding|Sign or Symptom|Discharge Instructions|16380,16397|false|false|false|C0028643|Numbness|loss of sensation
Event|Event|Discharge Instructions|16388,16397|false|false|false|||sensation
Finding|Finding|Discharge Instructions|16388,16397|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|Discharge Instructions|16388,16397|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|Discharge Instructions|16388,16397|false|false|false|C2229507|sensory exam|sensation
Anatomy|Anatomical Structure|Discharge Instructions|16417,16421|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|16417,16421|false|false|false|C0152338;C0444584;C0460148;C1268086;C4082212|Adult human body;Body structure;Human body structure;Structure of body of caudate nucleus;Whole body|body
Finding|Intellectual Product|Discharge Instructions|16417,16421|false|false|false|C1551342|Document Body|body
Procedure|Health Care Activity|Discharge Instructions|16460,16468|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|16469,16481|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|16469,16481|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|16469,16481|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

