CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Pharmaceutical Preparations|Drug|false|false||MEDICINEnull|Medicine|Title|false|false||MEDICINEnull|lisinopril|Drug|false|false||lisinopril
null|lisinopril|Drug|false|false||lisinoprilnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Diabetic foot ulcer|Disorder|false|false|C4299097;C0016504|diabetic foot ulcernull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false||diabeticnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C1456868;C0206172;C0041582;C1547940;C1550672;C0085119|foot
null|Foot|Anatomy|false|false|C0555980;C1456868;C0206172;C0041582;C1547940;C1550672;C0085119|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C4299097;C0016504|ulcer
null|null|Finding|false|false|C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C4299097;C0016504|ulcernull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Hallux structure|Anatomy|false|false|C0332840;C0002688;C1546539|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|Poorly controlled|Finding|false|false||poorly controllednull|Bad|Modifier|false|false||poorlynull|Disease Controlled|Finding|false|false||controlled
null|Control function|Finding|false|false||controlled
null|Controlled mark|Finding|false|false||controllednull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Retinal Diseases|Disorder|false|false||retinopathynull|Neuropathy|Disorder|false|false||neuropathynull|Pad Dosage Form|Drug|false|false|C3669270|PADnull|Pad Mass|Disorder|false|false|C3669270|PAD
null|Peripheral Arterial Diseases|Disorder|false|false|C3669270|PADnull|PADI4 wt Allele|Finding|false|false|C3669270|PAD
null|PADI4 gene|Finding|false|false|C3669270|PAD
null|DHX40 gene|Finding|false|false|C3669270|PADnull|PAD Regimen|Procedure|false|false|C3669270|PADnull|Strucure of thick cushion of skin|Anatomy|false|false|C2347441;C0332568;C1704436;C3540603;C1425478;C1425244;C0555980;C0085119;C0041582;C1547940;C1550672;C3814046|PADnull|Pad Device|Device|false|false||PAD
null|Pads|Device|false|false||PADnull|Pad (unit of presentation)|LabModifier|false|false||PAD
null|Pad Dosing Unit|LabModifier|false|false||PADnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504;C3669270|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504;C3669270|footnull|Lower extremity>Foot|Anatomy|false|false|C1956346;C0010068;C0175816;C0085119;C0555980;C4284121;C3813548;C1428349;C1413983;C2239547;C1413078;C0280573;C0170509;C0011905;C1707433;C0041582;C1547940;C1550672|foot
null|Foot|Anatomy|false|false|C1956346;C0010068;C0175816;C0085119;C0555980;C4284121;C3813548;C1428349;C1413983;C2239547;C1413078;C0280573;C0170509;C0011905;C1707433;C0041582;C1547940;C1550672|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C3669270;C4299097;C0016504|ulcer
null|null|Finding|false|false|C3669270;C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C3669270;C4299097;C0016504|ulcernull|Hallux structure|Anatomy|false|false|C0280573;C0170509;C0011905;C1707433;C1956346;C0010068;C0175816|halluxnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false|C4299097;C0016504;C0018534|CAD
null|Coronary heart disease|Disorder|false|false|C4299097;C0016504;C0018534|CAD
null|Coronary Artery Disease|Disorder|false|false|C4299097;C0016504;C0018534|CADnull|CAD gene|Finding|false|false|C4299097;C0016504|CAD
null|CALD1 wt Allele|Finding|false|false|C4299097;C0016504|CAD
null|B4GALNT2 gene|Finding|false|false|C4299097;C0016504|CAD
null|DFFB wt Allele|Finding|false|false|C4299097;C0016504|CAD
null|ACOD1 gene|Finding|false|false|C4299097;C0016504|CAD
null|DFFB gene|Finding|false|false|C4299097;C0016504|CADnull|cytarabine/daunorubicin protocol|Procedure|false|false|C4299097;C0016504;C0018534|CAD
null|Computer Assisted Diagnosis|Procedure|false|false|C4299097;C0016504;C0018534|CAD
null|Collision-Induced Dissociation|Procedure|false|false|C4299097;C0016504;C0018534|CAD
null|CyADIC regimen|Procedure|false|false|C4299097;C0016504;C0018534|CADnull|Caddo language|Entity|false|false||CADnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|Agreement (document)|Finding|false|false||agreement
null|Agreement|Finding|false|false||agreementnull|null|Attribute|false|false||agreementnull|3 Days|Time|false|false||3 daysnull|day|Time|false|false||daysnull|subjective (symptom)|Finding|false|false||subjectivenull|null|Attribute|false|false||subjectivenull|Subjective observation (qualifier value)|Modifier|false|false||subjectivenull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Chills|Finding|false|false||chillsnull|Administration Method - Pain|Finding|false|false|C0018534|pain
null|Pain|Finding|false|false|C0018534|painnull|null|Attribute|false|false||painnull|Hallux structure|Anatomy|false|false|C1424898;C1549543;C0030193|great toenull|RXFP2 gene|Finding|false|false|C0040357;C4299090;C0018534|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C1424898|toe
null|Toes|Anatomy|false|false|C1424898|toenull|Recent|Time|false|false||recentlynull|Specimen Type - Ulcer|Finding|false|false||ulcer
null|null|Finding|false|false||ulcer
null|Ulcer|Finding|false|false||ulcernull|Podiatry (discipline)|Title|false|false||podiatrynull|Specimen Type - Ulcer|Finding|false|false||ulcer
null|null|Finding|false|false||ulcer
null|Ulcer|Finding|false|false||ulcernull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Prostatic Intraepithelial Neoplasias|Disorder|false|false||pinnull|DYNLL1 gene|Finding|false|false||pinnull|Pin Device Component|Device|false|false||pin
null|Medical pins|Device|false|false||pin
null|Pins - Internal fixators|Device|false|false||pinnull|span - body measurement finding|Finding|false|false||span
null|Span - parameter|Finding|false|false||spannull|Span Distance|LabModifier|false|false||spannull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Tennis (activity)|Finding|false|false||tennisnull|Ball Device|Device|false|false||ballnull|Presentation|Finding|false|false||Presentednull|Urgent Care|Device|false|false||urgent carenull|Urgent Care|Entity|false|false||urgent carenull|Certification patient type - Urgent|Finding|false|false||urgent
null|Admission Type - Urgent|Finding|false|false||urgent
null|Triage Code - Urgent|Finding|false|false||urgent
null|Visit Priority Code - Urgent|Finding|false|false||urgentnull|Act Priority - urgent|Time|false|false||urgentnull|Urgent|Modifier|false|false||urgentnull|urgent - premium|LabModifier|false|false||urgentnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Fever|Finding|false|false||febrilenull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|Apyrexial|Finding|false|false||afebrilenull|arrival - ActRelationshipType|Finding|false|false||arrivalnull|null|Event|false|false||arrivalnull|Sustained|Finding|false|false||sustainednull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Podiatry (discipline)|Title|false|false||Podiatrynull|Traumatic Wound|Disorder|false|false|C0018534|wound
null|Wounds and Injuries|Disorder|false|false|C0018534|wound
null|Traumatic injury|Disorder|false|false|C0018534|woundnull|Route of Administration - Wound|Finding|false|false|C0018534|wound
null|null|Finding|false|false|C0018534|wound
null|Specimen Type - Wound|Finding|false|false|C0018534|woundnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Medial|Modifier|false|false||medialnull|Hallux structure|Anatomy|false|false|C1549529;C1547965;C1550680;C3263723;C0043251;C0043250|halluxnull|Probes|Device|false|false||probesnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|bone
null|null|Finding|false|false|C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|Message Waiting Priority - High|Finding|false|false||high
null|high - ActExposureLevelCode|Finding|false|false||high
null|IPSS Risk Category High|Finding|false|false||high
null|IPSS-R Risk Category High|Finding|false|false||high
null|High (finding)|Finding|false|false||highnull|Observation Value - High|Modifier|false|false||high
null|High|Modifier|false|false||high
null|Abnormally high|Modifier|false|false||highnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|X-rays, Homeopathic Preparations|Drug|false|false||X-raysnull|Plain x-ray|Procedure|false|false||X-rays
null|Diagnostic radiologic examination|Procedure|false|false||X-raysnull|Roentgen Rays|Phenomenon|false|false||X-raysnull|Bony|Finding|false|false||bonynull|Superficial ulcer|Disorder|false|false||erosionnull|Erosion lesion|Finding|false|false||erosionnull|Subcutaneous Route of Administration|Finding|true|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Gas - SpecimenType|Drug|true|false||gas
null|Gases|Drug|true|false||gas
null|Gas Dosage Form|Drug|true|false||gasnull|Gas - Specimen Source Codes|Finding|true|false||gas
null|gastrointestinal gas|Finding|true|false||gas
null|PAGR1 wt Allele|Finding|true|false||gas
null|GALNS wt Allele|Finding|true|false||gas
null|GALNS gene|Finding|true|false||gas
null|GAST wt Allele|Finding|true|false||gas
null|GAST gene|Finding|true|false||gas
null|germacrene-A synthase activity|Finding|true|false||gas
null|PAGR1 gene|Finding|true|false||gasnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||Plannull|Treatment Plan|Finding|false|false||Plan
null|Planned|Finding|false|false||Plan
null|null|Finding|false|false||Plannull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Target Awareness - partial|Finding|false|false|C0040357;C4299090;C0018534|partialnull|Partial|LabModifier|false|false||partialnull|Amputation of left great toe|Procedure|false|false|C0040357;C4299090;C0018534|amputation of left great toenull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0040357;C4299090;C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0040357;C4299090;C0018534|amputationnull|Amputation|Procedure|false|false|C0018534;C0040357;C4299090|amputationnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C4316611;C0002688;C1550516;C0332840;C1552822;C1424898;C1546539|great toenull|RXFP2 gene|Finding|false|false|C0018534|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C0332840;C1550516;C4316611;C1546539;C0002688|toe
null|Toes|Anatomy|false|false|C0332840;C1550516;C4316611;C1546539;C0002688|toenull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|abdnull|ABD (body structure)|Anatomy|false|false|C3811055;C1549543;C0030193|abd
null|Abdomen|Anatomy|false|false|C3811055;C1549543;C0030193|abdnull|Administration Method - Pain|Finding|false|false|C0449202;C0000726|pain
null|Pain|Finding|false|false|C0449202;C0000726|painnull|null|Attribute|false|false||painnull|rectal discharge diarrhea (physical finding)|Finding|false|false||diarrhea
null|Diarrhea|Finding|false|false||diarrheanull|excessive urination|Finding|false|false||excessive urinationnull|Excessive (qualifier value)|Modifier|false|false||excessivenull|Urination|Finding|false|false||urinationnull|Orthostasis|Finding|false|false||orthostasis
null|Orthostatic intolerance|Finding|false|false||orthostasisnull|null|Finding|false|false||dyspnea
null|Dyspnea|Finding|false|false||dyspneanull|Chest Pain|Finding|false|false|C1527391;C0817096|chest painnull|null|Attribute|false|false|C1527391;C0817096|chest painnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C1549543;C0030193;C0008031;C2926613|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C1549543;C0030193;C0008031;C2926613|chestnull|Administration Method - Pain|Finding|false|false|C1527391;C0817096|pain
null|Pain|Finding|false|false|C1527391;C0817096|painnull|null|Attribute|false|false||painnull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Taking vital signs|Procedure|false|false||vital signsnull|null|Attribute|false|false||vital signs
null|Vital signs|Attribute|false|false||vital signsnull|Vital High Nitrogen Enteral Nutrition|Drug|false|false||vitalnull|Vital (qualifier value)|Modifier|false|false||vitalnull|Aspects of signs|Finding|false|false||signs
null|Physical findings|Finding|false|false||signsnull|Manufactured sign|Device|false|false||signsnull|Apyrexial|Finding|false|false||afebrilenull|Tachycardia by ECG Finding|Finding|false|false||tachycardia
null|Tachycardia|Finding|false|false||tachycardianull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Feels warm|Finding|false|false||warmnull|warming process|Phenomenon|false|false||warmnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Diaphoretic|Modifier|false|false||diaphoreticnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false|C0024109|Respnull|Respiratory rate|Attribute|false|false||Respnull|Lung|Anatomy|false|false|C0851355;C1550016|lungsnull|Remote control command - Clear|Finding|false|false|C0024109|clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Medullary sponge kidney|Disorder|false|false||MSK
null|Medullary sponge kidney|Disorder|false|false||MSKnull|SIK1 gene|Finding|false|false||MSKnull|Erythema|Disorder|false|false|C0040357;C4299090;C2987514;C0018534|erythemanull|Hallux structure|Anatomy|false|false|C0041834|big toenull|Large|LabModifier|false|false||bignull|Lower extremity>Toes|Anatomy|false|false|C0041834|toe
null|Toes|Anatomy|false|false|C0041834|toenull|Tracking|Modifier|false|false||trackingnull|inferiority|Finding|false|false|C2987514|inferiornull|Inferior|Modifier|false|false||inferiornull|nitrogenous base|Drug|false|false|C2987514|base
null|Base|Drug|false|false|C2987514|base
null|Dental Base|Drug|false|false|C2987514|base
null|base - RoleClass|Drug|false|false|C2987514|basenull|Base - General Qualifier|Finding|false|false|C2987514|base
null|BPIFA4P gene|Finding|false|false|C2987514|base
null|Base - RX Component Type|Finding|false|false|C2987514|basenull|Anatomical base|Anatomy|false|false|C0041834;C1549548;C1705938;C1843354;C0678975;C1704464;C0178499;C1550601;C1880279|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Emotional tenderness|Finding|false|false|C0230445;C1305418;C0489800|Tenderness
null|Sore to touch|Finding|false|false|C0230445;C1305418;C0489800|Tendernessnull|Tracking|Modifier|false|false||trackingnull|Pathname|Finding|false|false|C0230445;C1305418;C0489800|pathnull|Pathology procedure|Procedure|false|false|C0489800;C0230445;C1305418|pathnull|RXFP2 gene|Finding|false|false|C0489800;C0230445;C1305418|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Posterior part of left leg|Anatomy|false|false|C0684239;C0234233;C0919386;C1424898;C1705483|L calfnull|Structure of calf of leg|Anatomy|false|false|C0684239;C0234233;C1424898;C0919386;C1705483|calf
null|null|Anatomy|false|false|C0684239;C0234233;C1424898;C0919386;C1705483|calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Limited component (foundation metadata concept)|Finding|false|false||Limited
null|Limited (extensiveness)|Finding|false|false||Limitednull|Plantar flexion|Finding|false|false|C0442036;C0230463|plantar flexionnull|Plantar (qualifier value)|Anatomy|false|false|C0231452;C0231784|plantar
null|Sole of Foot|Anatomy|false|false|C0231452;C0231784|plantarnull|null|Finding|false|false|C0442036;C0230463|flexionnull|W flexion|Attribute|false|false||flexionnull|Limited component (foundation metadata concept)|Finding|false|false||Limited
null|Limited (extensiveness)|Finding|false|false||Limitednull|Rupture of Membranes|Finding|false|false|C0003086;C0003087;C4284979|ROM
null|ROM1 gene|Finding|false|false|C0003086;C0003087;C4284979|ROMnull|Range of motion technique (procedure)|Procedure|false|false|C0003086;C0003087;C4284979|ROMnull|Read Only Memory Device|Device|false|false||ROMnull|Romani Language|Entity|false|false||ROMnull|Lower extremity>Ankle|Anatomy|false|false|C1419600;C0948106;C1562926|ankle
null|Ankle|Anatomy|false|false|C1419600;C0948106;C1562926|ankle
null|Ankle joint structure|Anatomy|false|false|C1419600;C0948106;C1562926|anklenull|Lower extremity>Toes|Anatomy|false|false||toe
null|Toes|Anatomy|false|false||toenull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Long Interspersed Elements|Drug|false|false||Lines
null|Long Interspersed Elements|Drug|false|false||Linesnull|Lines Quantity Limit Request|Finding|false|false||Linesnull|Lines - QueryQuantityUnit|Modifier|false|false||Lines
null|Linear|Modifier|false|false||Linesnull|Drain device|Device|false|false||Drainsnull|20 gauge|LabModifier|false|false||20g
null|20 grams|LabModifier|false|false||20gnull|Structure of left hand|Anatomy|false|false|C0741992|L handnull|Hand problem|Finding|false|false|C4285005;C0018563;C0230371|handnull|Upper extremity>Hand|Anatomy|false|false|C0741992|hand
null|Hand|Anatomy|false|false|C0741992|handnull|Laboratory test finding|Lab|false|false||Labsnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|White (population group)|Subject|false|false||Whites
null|Caucasian|Subject|false|false||Whites
null|Caucasians|Subject|false|false||Whitesnull|Neut brand of sodium bicarbonate|Drug|false|false||neut
null|Neut brand of sodium bicarbonate|Drug|false|false||neutnull|Neutralization Tests|Procedure|false|false||neutnull|Scientific Study|Procedure|false|false||Studiesnull|Diagnostic radiologic examination|Procedure|false|false|C4299097;C0016504|Xraynull|Roentgen Rays|Phenomenon|false|false|C4299097;C0016504|Xraynull|Foot problem|Finding|false|false|C4299097;C0016504|Footnull|Lower extremity>Foot|Anatomy|false|false|C0043299;C0043309;C0555980|Foot
null|Foot|Anatomy|false|false|C0043299;C0043309;C0555980|Footnull|Foot Unit of Length|LabModifier|false|false||Footnull|LAT protein, human|Drug|false|false||Lat
null|L-Type Amino Acid Transporter|Drug|false|false||Lat
null|L-Type Amino Acid Transporter|Drug|false|false||Lat
null|ORC3 protein, human|Drug|false|false||Lat
null|ORC3 protein, human|Drug|false|false||Lat
null|LAT protein, human|Drug|false|false||Latnull|LAT gene|Finding|false|false||Lat
null|ORC3 wt Allele|Finding|false|false||Lat
null|ORC3 gene|Finding|false|false||Lat
null|SPNS1 gene|Finding|false|false||Latnull|Latin Language|Entity|false|false||Latnull|Table Cell Horizontal Align - left|Finding|false|false||Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Reading (datum presentation)|Finding|false|false||read
null|Do Reading Question|Finding|false|false||read
null|Reading (activity)|Finding|false|false||readnull|Nucleotide Sequence Read|Procedure|false|false||readnull|Ulceration|Finding|false|false|C0040357;C4299090;C0018534|ulceration
null|Ulcer|Finding|false|false|C0040357;C4299090;C0018534|ulcerationnull|Medial|Modifier|false|false||medialnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Aspect (characteristic)|Modifier|false|false||aspectnull|Aspect - Kind of quantity|LabModifier|false|false||aspectnull|Hallux structure|Anatomy|false|false|C1424898;C3887532;C0041582|great toenull|RXFP2 gene|Finding|false|false|C0018534;C0040357;C4299090|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C3887532;C0041582;C1424898|toe
null|Toes|Anatomy|false|false|C3887532;C0041582;C1424898|toenull|Superficial ulcer|Disorder|false|false|C0576464;C3669027;C0223792;C0222682;C2987514|erosionnull|Erosion lesion|Finding|false|false|C0576464;C3669027;C2987514;C0223792;C0222682|erosionnull|Medial|Modifier|false|false||medialnull|nitrogenous base|Drug|false|false|C0223792;C0222682;C0576464;C3669027;C2987514|base
null|Base|Drug|false|false|C0223792;C0222682;C0576464;C3669027;C2987514|base
null|Dental Base|Drug|false|false|C0223792;C0222682;C0576464;C3669027;C2987514|base
null|base - RoleClass|Drug|false|false|C0223792;C0222682;C0576464;C3669027;C2987514|basenull|Base - General Qualifier|Finding|false|false|C0576464;C3669027;C0223792;C0222682;C2987514|base
null|BPIFA4P gene|Finding|false|false|C0576464;C3669027;C0223792;C0222682;C2987514|base
null|Base - RX Component Type|Finding|false|false|C0576464;C3669027;C0223792;C0222682;C2987514|basenull|Anatomical base|Anatomy|false|false|C1959609;C1549548;C1705938;C1843354;C0333307;C1704464;C0178499;C1550601;C1880279|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Bone structure of distal phalanx|Anatomy|false|false|C1959609;C1424898;C1549548;C1705938;C1843354;C0333307;C1704464;C0178499;C1550601;C1880279;C4522154|distal phalanx
null|null|Anatomy|false|false|C1959609;C1424898;C1549548;C1705938;C1843354;C0333307;C1704464;C0178499;C1550601;C1880279;C4522154|distal phalanxnull|Distal Resection Margin|Attribute|false|false|C0576464;C3669027;C0223792;C0222682|distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Phalanx of hand|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C1424898;C0333307;C1549548;C1705938;C1843354;C1959609;C4522154|phalanx
null|Phalanx structure|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C1424898;C0333307;C1549548;C1705938;C1843354;C1959609;C4522154|phalanxnull|RXFP2 gene|Finding|false|false|C0576464;C3669027;C0223792;C0222682|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C1552654|toe
null|Toes|Anatomy|false|false|C1552654|toenull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Parameterized Data Type - Interval|Finding|false|false|C0040357;C4299090|intervalnull|Interval|Time|false|false||intervalnull|findings aspects|Finding|false|false||Findingsnull|null|Attribute|false|false||Findingsnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|MRI with contrast|Procedure|false|false||MRI with contrastnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Further|Modifier|false|false||furthernull|Knowledge acquisition using a method of assessment|Finding|false|false||assessmentnull|assessment of cognitive functions|Procedure|false|false||assessment
null|Physical Examination|Procedure|false|false||assessment
null|Nutrition Assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Personal care assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Evaluation procedure|Procedure|false|false||assessment
null|Evaluation|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessmentnull|Assessed|Event|false|false||assessmentnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|piperacillin-tazobactam combination|Drug|false|false||Piperacillin-Tazobactamnull|piperacillin|Drug|false|false||Piperacillin
null|piperacillin|Drug|false|false||Piperacillinnull|tazobactam|Drug|false|false||Tazobactam
null|tazobactam|Drug|false|false||Tazobactamnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Consultation|Procedure|false|false||Consultsnull|Podiatry (discipline)|Title|false|false||Podiatrynull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|arrival - ActRelationshipType|Finding|false|false|C3714591|arrivalnull|null|Event|false|false||arrivalnull|Floor (anatomic)|Anatomy|false|false|C1578483;C1550655;C1578481;C1578486;C1578484;C1578485;C1555577|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false|C3714591|patient
null|Specimen Type - Patient|Finding|false|false|C3714591|patient
null|Mail Claim Party - Patient|Finding|false|false|C3714591|patient
null|Report source - Patient|Finding|false|false|C3714591|patient
null|null|Finding|false|false|C3714591|patient
null|Disabled Person Code - Patient|Finding|false|false|C3714591|patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|Chills|Finding|false|false||chillsnull|Blanket|Device|false|false||blanketsnull|Structure of left foot|Anatomy|false|false|C1552822;C0555980|Left footnull|Table Cell Horizontal Align - left|Finding|false|false|C4299097;C0016504;C0230461|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C1552822;C0555980|foot
null|Foot|Anatomy|false|false|C1552822;C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Gauze dressing|Device|false|false||gauze dressingnull|Gauzes|Device|false|false||gauzenull|Dressing Dosage Form|Drug|false|false||dressingnull|Ability to dress|Finding|false|false||dressing
null|null|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Very|Modifier|false|false||verynull|Tender|Modifier|false|false||tendernull|Review of systems (procedure)|Procedure|false|false||REVIEW OF SYSTEMSnull|null|Attribute|false|false||REVIEW OF SYSTEMS
null|null|Attribute|false|false||REVIEW OF SYSTEMSnull|Review of|Finding|false|false||REVIEW OFnull|Review (Publication Type)|Finding|false|false||REVIEW
null|Act Class - review|Finding|false|false||REVIEWnull|System|Finding|false|false||SYSTEMSnull|Complete, Multiple Vitamins with Iron|Drug|false|false||Complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||Complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||Completenull|Completion Status for valid values - Complete|Finding|false|false|C0262327|Complete
null|Data operation - complete|Finding|false|false|C0262327|Complete
null|Finish - dosing instruction imperative|Finding|false|false|C0262327|Completenull|Complete|Modifier|false|false||Completenull|Reactive Oxygen Species|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|rosiglitazone|Drug|false|false|C0262327|ROS
null|Reactive Oxygen Species|Drug|false|false|C0262327|ROSnull|ROS1 wt Allele|Finding|false|false|C0262327|ROS
null|ROS1 gene|Finding|false|false|C0262327|ROSnull|Review of systems (procedure)|Procedure|false|false|C0262327|ROSnull|rostral sulcus|Anatomy|false|false|C1548561;C3853530;C1706059;C0289313;C0162772;C0812281;C1709820;C0489633|ROSnull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|COPD pharmacologic substance|Drug|false|false||COPDnull|Chronic obstructive pulmonary disease of horses|Disorder|false|false||COPD
null|Chronic Obstructive Airway Disease|Disorder|false|false||COPDnull|ARCN1 gene|Finding|false|false||COPDnull|DFFB protein, human|Drug|false|false||CAD
null|DFFB protein, human|Drug|false|false||CADnull|Cold Hemagglutinin Disease|Disorder|false|false||CAD
null|Coronary heart disease|Disorder|false|false||CAD
null|Coronary Artery Disease|Disorder|false|false||CADnull|CAD gene|Finding|false|false||CAD
null|CALD1 wt Allele|Finding|false|false||CAD
null|B4GALNT2 gene|Finding|false|false||CAD
null|DFFB wt Allele|Finding|false|false||CAD
null|ACOD1 gene|Finding|false|false||CAD
null|DFFB gene|Finding|false|false||CADnull|cytarabine/daunorubicin protocol|Procedure|false|false||CAD
null|Computer Assisted Diagnosis|Procedure|false|false||CAD
null|Collision-Induced Dissociation|Procedure|false|false||CAD
null|CyADIC regimen|Procedure|false|false||CADnull|Caddo language|Entity|false|false||CADnull|Burning Mouth Syndrome|Disorder|false|false|C0226032|BMSnull|Proximal Resection Margin|Attribute|false|false||proximalnull|Proximal|Modifier|false|false||proximalnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738;C1413980;C4551552;C0006430|LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false|C0226032;C0226032|DESnull|DES gene|Finding|false|false|C0226032;C0226032|DESnull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1413980;C5550999;C0398738;C4551552;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Graph Edge|Finding|false|false||edgenull|Along edge (qualifier value)|Modifier|false|false||edgenull|integrated stress response signaling|Finding|false|false|C0226032|ISRnull|Middle|Modifier|false|false||midnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738;C5445058;C4551552;C1413980|LADnull|Ladino Language|Entity|false|false||LADnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false|C0226032|DESnull|DES gene|Finding|false|false|C0226032|DESnull|Stenosis|Finding|false|false||stenosisnull|Stenosis <Pimeliinae>|Entity|false|false||stenosisnull|Stenosis Morphology|Modifier|false|false||stenosisnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|null|Device|false|false||stentnull|DES protein, human|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|Desmosine|Drug|false|false||DES
null|DES protein, human|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DES
null|diethylstilbestrol|Drug|false|false||DESnull|CEREBELLAR ATAXIA, IMPAIRED INTELLECTUAL DEVELOPMENT, AND DYSEQUILIBRIUM SYNDROME 1|Disorder|false|false||DESnull|DES gene|Finding|false|false||DESnull|Coronary Artery Bypass Surgery|Procedure|false|false||CABGnull|Lima|Entity|false|false||LIMAnull|Leukocyte adhesion deficiency type 1|Disorder|false|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|false|false|C0226032|LADnull|ITGB2 wt Allele|Finding|false|false|C0226032|LAD
null|DLD gene|Finding|false|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C5550999;C0398738;C1414063;C1706333|LADnull|Ladino Language|Entity|false|false||LADnull|Scalable Vector Graphics|Entity|false|false||SVGnull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Migraine Disorders|Disorder|false|false||Migrainesnull|shoulder pain chronic|Disorder|false|false|C0037004;C4299050|Chronic shoulder painnull|Chronic - Admission Level of Care Code|Finding|false|false|C0037004;C4299050|Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false|C0037004;C4299050|Chronicnull|chronic|Time|false|false||Chronicnull|Shoulder Pain|Finding|false|false|C0037004;C4299050|shoulder painnull|Procedures on Shoulder|Procedure|false|false|C0037004;C4299050|shoulder
null|Examination of shoulder(s)|Procedure|false|false|C0037004;C4299050|shouldernull|Upper extremity>Shoulder|Anatomy|false|false|C1547296;C0037011;C0869975;C0221590;C2598155;C0748678;C1555457;C1549543;C0030193|shoulder
null|Shoulder|Anatomy|false|false|C1547296;C0037011;C0869975;C0221590;C2598155;C0748678;C1555457;C1549543;C0030193|shouldernull|Administration Method - Pain|Finding|false|false|C0037004;C4299050|pain
null|Pain|Finding|false|false|C0037004;C4299050|painnull|null|Attribute|false|false|C0037004;C4299050|painnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|OSA protein, Drosophila|Drug|false|false||OSA
null|OSA protein, Drosophila|Drug|false|false||OSAnull|Sleep Apnea, Obstructive|Disorder|false|false||OSAnull|Osa <eudicots>|Entity|false|false||OSA
null|Osage language|Entity|false|false||OSA
null|Osa|Entity|false|false||OSAnull|Peripheral Neuropathy|Disorder|false|false||Peripheral neuropathy
null|Peripheral Nervous System Diseases|Disorder|false|false||Peripheral neuropathynull|Peripheral|Modifier|false|false||Peripheralnull|Neuropathy|Disorder|false|false||neuropathynull|Restless Legs Syndrome|Disorder|false|false|C1140621;C0023216|Restless legnull|Restlessness|Finding|false|false|C1140621;C0023216|Restless
null|Agitation|Finding|false|false|C1140621;C0023216|Restlessnull|Leg|Anatomy|false|false|C0085631;C3887611;C0035258|leg
null|Lower Extremity|Anatomy|false|false|C0085631;C3887611;C0035258|legnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Ward (environment)|Device|false|false||wardnull|Ward (person)|Subject|false|false||wardnull|Ward (environment)|Entity|false|false||wardnull|Full|Modifier|false|false||fullnull|Details|Modifier|false|false||detailsnull|Relationship - Mother|Finding|false|false||Mothernull|Mother (person)|Subject|false|false||Mothernull|Possible|Finding|false|false||possiblenull|Possible diagnosis|Modifier|false|false||possible
null|Possibly Related to Intervention|Modifier|false|false||possiblenull|Alcohol abuse|Disorder|false|false||alcohol abusenull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Drug abuse|Disorder|false|false||abusenull|Victim of abuse (finding)|Finding|false|false||abusenull|Abuse|Event|false|false||abusenull|Indirect exposure mechanism - Father|Finding|false|false||Father
null|Relationship - Father|Finding|false|false||Father
null|Father - courtesy title|Finding|false|false||Fathernull|Father (person)|Subject|false|false||Fathernull|Deceased - ActIneligibilityReason|Finding|false|false||deceased
null|Deceased - Military Status|Finding|false|false||deceased
null|Cessation of life|Finding|false|false||deceasednull|Hodgkin Disease|Disorder|false|false||Hodgkin's Diseasenull|Hodgkin Disease|Disorder|false|false||Hodgkinnull|Disease|Disorder|false|false||Diseasenull|Old|Time|false|false||oldnull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||GENERALnull|General medical service|Procedure|false|false||GENERALnull|Generalized|Modifier|false|false||GENERALnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|patient appears in no acute distress (physical finding)|Finding|false|false||In no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|HEENT|Anatomy|false|false||HEENTnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Cardiac attachment|Finding|false|false|C0018787|CARDIACnull|Heart|Anatomy|false|false|C1314974|CARDIACnull|Cardiac - anatomy qualifier|Modifier|false|false||CARDIACnull|MAS1L gene|Finding|true|false||MRGnull|Lung|Anatomy|false|false||LUNGSnull|Cancer/Testis Antigen|Drug|false|false||CTAnull|PCYT1A wt Allele|Finding|false|false||CTA
null|CERNA3 gene|Finding|false|false||CTAnull|Cardiac Computerized Tomographic Angiography|Procedure|false|false||CTAnull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|ABDOMENnull|Abdomen problem|Finding|false|false|C0230168;C0000726|ABDOMENnull|Abdomen|Anatomy|false|false|C0941288;C0153662|ABDOMEN
null|Abdominal Cavity|Anatomy|false|false|C0941288;C0153662|ABDOMENnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Deep palpation|Procedure|false|false||deep palpationnull|Deep Resection Margin|Attribute|false|false||deepnull|Deep (qualifier value)|Modifier|false|false||deepnull|Palpation|Procedure|false|false||palpationnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|All extremities|Anatomy|false|false||EXTREMITIES
null|Limb structure|Anatomy|false|false||EXTREMITIESnull|Structure of left foot|Anatomy|false|false|C0555980;C1552822|left footnull|Table Cell Horizontal Align - left|Finding|false|false|C4299097;C0016504;C0230461|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C0230461;C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C1552822;C0555980|foot
null|Foot|Anatomy|false|false|C1552822;C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Gauze dressing|Device|false|false||gauze dressingnull|Gauzes|Device|false|false||gauzenull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing patient (procedure)|Procedure|false|false||dressing
null|Dressing of skin or wound|Procedure|false|false||dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|MILDLY|Modifier|false|false||mildly
null|Mild (qualifier value)|Modifier|false|false||mildlynull|erythematous|Finding|false|false||erythematousnull|Very|Modifier|false|false||verynull|Tender|Modifier|false|false||tendernull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Edema|Finding|true|false||edemanull|null|Attribute|true|false||edemanull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurologic (qualifier value)|Modifier|false|false||NEUROLOGICnull|Sensory (qualifier value)|Modifier|false|false||Sensorynull|Motor function (finding)|Finding|false|false||motor functionnull|Motor function (observable entity)|Phenomenon|false|false||motor functionnull|motor movement|Finding|false|false||motornull|Motor Device|Device|false|false||motornull|Function (attribute)|Finding|false|false||function
null|physiological aspects|Finding|false|false||function
null|Mathematical Operator|Finding|false|false||function
null|Functional Status|Finding|false|false||functionnull|Function Axis|Subject|false|false||functionnull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|general appearance (physical finding)|Finding|false|false||General Appearancenull|null|Attribute|false|false||General Appearancenull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Generalnull|General medical service|Procedure|false|false||Generalnull|Generalized|Modifier|false|false||Generalnull|patient appearance regarding mental status exam|Procedure|false|false||Appearancenull|null|Attribute|false|false||Appearancenull|Personal appearance|Subject|false|false||Appearancenull|Appearance|Modifier|false|false||Appearancenull|Kind of quantity - Appearance|LabModifier|false|false||Appearancenull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|HEENT|Anatomy|false|false||HEENTnull|Scleral Diseases|Disorder|false|false|C0036410|Scleranull|examination of sclera|Procedure|false|false|C0036410|Scleranull|Sclera|Anatomy|false|false|C0205180;C0036412;C2228481|Scleranull|Anicteric|Finding|false|false|C0036410|anictericnull|Myelofibrosis|Disorder|false|false|C0694605|MMMnull|Medial part of medial mammillary nucleus|Anatomy|false|false|C0026987|MMMnull|Disorder of oropharynx|Disorder|false|false|C0521367|oropharyngealnull|Oropharyngeal Route of Administration|Finding|false|false|C0521367|oropharyngealnull|Oropharyngeal|Anatomy|false|false|C0221198;C0553694;C1522409|oropharyngealnull|Lesion|Finding|false|false|C0521367|lesionsnull|Leukocyte adhesion deficiency type 1|Disorder|true|false|C0226032|LAD
null|Leukocyte adhesion deficiency|Disorder|true|false|C0226032|LADnull|ITGB2 wt Allele|Finding|true|false|C0226032|LAD
null|DLD gene|Finding|true|false|C0226032|LADnull|Anterior descending branch of left coronary artery|Anatomy|false|false|C1414063;C1706333;C5550999;C0398738|LADnull|Ladino Language|Entity|true|false||LADnull|Lung|Anatomy|false|false||Lungsnull|Relational Operator - Equal|Finding|false|false||Equalnull|Equal|Modifier|false|false||Equalnull|Chest rise|Finding|false|false|C1527391;C0817096|chest risenull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C4321377;C5570649|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C4321377;C5570649|chestnull|risedronate|Drug|false|false||rise
null|risedronate|Drug|false|false||risenull|Relational and Item-Specific Encoding Task|Finding|false|false|C1527391;C0817096|risenull|Language Ability Proficiency - Good|Finding|false|false||Good
null|Language Proficiency - Good|Finding|false|false||Goodnull|Specimen Quality - Good|Modifier|false|false||Good
null|Good|Modifier|false|false||Goodnull|Air Movements|Phenomenon|false|false||air movementnull|Air (substance)|Drug|false|false||air
null|air|Drug|false|false||air
null|air|Drug|false|false||airnull|ACUTE INSULIN RESPONSE|Finding|false|false||air
null|AIRN gene|Finding|false|false||air
null|AI/RHEUM|Finding|false|false||airnull|Movement|Finding|false|false||movementnull|Increased (finding)|Finding|true|false||increased
null|Increase|Finding|true|false||increasednull|Increased|LabModifier|false|false||increasednull|Work|Event|true|false||worknull|outcomes otolaryngology breathing|Finding|false|false||breathing
null|Inspiration (function)|Finding|false|false||breathing
null|Respiration|Finding|false|false||breathingnull|null|Attribute|false|false||breathingnull|respiratory system process|Phenomenon|false|false||breathingnull|Decreased breath sounds|Finding|false|false|C1261077|Decreased breath soundsnull|null|Attribute|false|false|C1261077|breath sounds
null|Respiratory Sounds|Attribute|false|false|C1261077|breath soundsnull|Breath|Finding|false|false|C1261077|breathnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false|C1261077|soundsnull|Structure of left lower lobe of lung|Anatomy|false|false|C0037709;C0225386;C0035234;C3484186;C0238844|LLLnull|Basilar Rales|Finding|false|false|C2987514|Rales
null|Rales|Finding|false|false|C2987514|Ralesnull|Table Cell Horizontal Align - left|Finding|false|false|C2987514|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|nitrogenous base|Drug|false|false|C2987514|base
null|Base|Drug|false|false|C2987514|base
null|Dental Base|Drug|false|false|C2987514|base
null|base - RoleClass|Drug|false|false|C2987514|basenull|Base - General Qualifier|Finding|false|false|C2987514|base
null|BPIFA4P gene|Finding|false|false|C2987514|base
null|Base - RX Component Type|Finding|false|false|C2987514|basenull|Anatomical base|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C0240859;C0034642;C1552822;C1549548;C1705938;C1843354|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Wheezing|Finding|false|false||wheezesnull|Rhonchi|Finding|false|false||rhonchinull|Heart murmur|Finding|true|false||murmursnull|Pericardial friction rub|Finding|true|false||rubsnull|Carotid Arteries|Anatomy|false|false||carotidnull|Bruit|Finding|false|false||bruitsnull|Carotid Arteries|Anatomy|false|false|C0034107|carotidnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false|C0007272|pulsesnull|Radial|Finding|false|false||radial
null|Circumpennate|Finding|false|false||radialnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Dorsalis pedis pulse|Finding|false|false||dorsalis pedis pulsenull|Physiologic pulse|Finding|false|false||pulsenull|Pulse taking|Procedure|false|false||pulsenull|Pulse Rate|Attribute|false|false||pulsenull|Pulse phenomenon|Phenomenon|false|false||pulsenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Unable|Finding|false|false||unablenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Bandage Dosage Form|Drug|false|false||bandagenull|Bandage|Device|false|false||bandagenull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Bowel sounds|Finding|false|false|C0021853|Bowel soundsnull|Intestines|Anatomy|false|false|C0232693;C0037709;C0150312;C0449450|Bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false|C0021853|soundsnull|Present|Finding|false|false|C0021853|present
null|Presentation|Finding|false|false|C0021853|presentnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Palpation|Procedure|false|false||palpationnull|All extremities|Anatomy|false|false||Extremities
null|Limb structure|Anatomy|false|false||Extremitiesnull|Clubbing|Disorder|true|false||clubbingnull|Cyanosis|Finding|true|false||cyanosisnull|Structure of left foot|Anatomy|false|false|C1305428;C0518459;C1552822;C0152053;C0278286;C1705365;C0555980|Left footnull|Table Cell Horizontal Align - left|Finding|false|false|C0230461|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C0152053;C0278286;C1305428;C0518459;C0555980|foot
null|Foot|Anatomy|false|false|C0152053;C0278286;C1305428;C0518459;C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Dressing Dosage Form|Drug|false|false|C0230461|dressingnull|null|Finding|false|false|C4299097;C0016504;C0230461|dressing
null|Ability to dress|Finding|false|false|C4299097;C0016504;C0230461|dressingnull|Dressing patient (procedure)|Procedure|false|false|C4299097;C0016504;C0230461|dressing
null|Dressing of skin or wound|Procedure|false|false|C4299097;C0016504;C0230461|dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Cleaning (activity)|Event|false|false||cleannull|Erythema|Disorder|false|false|C1515974|Erythemanull|Edema|Finding|false|false|C1515974|edemanull|null|Attribute|false|false||edemanull|null|Finding|false|false|C1515974|marginnull|Marginal|Modifier|false|false||marginnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0543467;C0587668;C0013604;C0041834;C4761388;C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Suture Dosage Form|Drug|false|false|C0502420;C1515974|Suturenull|null|Finding|false|false|C1515974;C0502420|Suturenull|Closure by suture|Procedure|false|false|C0502420;C1515974|Suturenull|Suture Joint|Anatomy|false|false|C1706068;C0009068;C1546778;C1546803|Suturenull|Suture Device|Device|false|false||Suture
null|Surgical sutures|Device|false|false||Suturenull|null|Finding|false|false|C1515974;C0502420|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C1706068;C0034161;C1546758;C1546803;C0009068;C1947930|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Cleaning (activity)|Event|false|false|C1515974|cleannull|Pus specimen|Drug|true|false||pusnull|Pus Specimen Code|Finding|true|false|C1515974|pus
null|Pus|Finding|true|false|C1515974|pusnull|Pashtu language|Entity|true|false||pusnull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|Skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|Skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|Skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|Skinnull|Skin rash|Finding|true|false|C1515974|rashes
null|Exanthema|Finding|true|false|C1515974|rashesnull|Lesion|Finding|true|false|C1515974|lesionsnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0221198;C5779628;C0015230;C0543467;C0587668|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services|Finding|false|false||time
null|Time (foundation metadata concept)|Finding|false|false||time
null|Value type - Time|Finding|false|false||time
null|Instructions for Use of the CPT Codebook - Time|Finding|false|false||time
null|Data types - Time|Finding|false|false||time
null|null|Finding|false|false||timenull|Time|Time|false|false||timenull|Gender Status - Intact|Finding|false|false||intactnull|Intact|Modifier|false|false||intactnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0005768;C0229664;C0005767;C0851353|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|C-Reactive Protein, human|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-Reactive Protein, human|Drug|false|false||CRPnull|CRP wt Allele|Finding|false|false||CRP
null|CRP gene|Finding|false|false||CRP
null|CSRP1 gene|Finding|false|false||CRP
null|PPIAP10 gene|Finding|false|false||CRPnull|Pidgin and Creole language|Entity|false|false||CRPnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Partial pressure of Oxygen|Finding|false|false||pO2
null|US Military enlisted E5|Finding|false|false||pO2null|PO2 measurement|Procedure|false|false||pO2null|Carbon dioxide measurement, partial pressure|Procedure|false|false||pCO2null|Carbon dioxide, partial pressure|Lab|false|false||pCO2null|nitrogenous base|Drug|false|false|C2987514|Base
null|Base|Drug|false|false|C2987514|Base
null|Dental Base|Drug|false|false|C2987514|Base
null|base - RoleClass|Drug|false|false|C2987514|Basenull|Base - General Qualifier|Finding|false|false|C2987514|Base
null|BPIFA4P gene|Finding|false|false|C2987514|Base
null|Base - RX Component Type|Finding|false|false|C2987514|Basenull|Anatomical base|Anatomy|false|false|C1549548;C1705938;C1843354;C1704464;C0178499;C1550601;C1880279|Basenull|Base - unit of product usage|LabModifier|false|false||Basenull|lactate in blood (lab test)|Procedure|false|false||BLOOD Lactatenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|lactate|Drug|false|false||Lactate
null|lactate|Drug|false|false||Lactate
null|Lactates|Drug|false|false||Lactatenull|Lactic acid measurement|Procedure|false|false||Lactatenull|Color of urine|Finding|false|false||URINE Colornull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|color additive|Drug|false|false||Color
null|Coloring Excipient|Drug|false|false||Colornull|color - solid dosage form|Modifier|false|false||Color
null|Color|Modifier|false|false||Colornull|Color quantity|LabModifier|false|false||Colornull|Cereal plant straw|Drug|false|false||Strawnull|Straw package type|Device|false|false||Strawnull|Straw Color|Modifier|false|false||Strawnull|Straw (unit of presentation)|LabModifier|false|false||Strawnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Hematuria|Disorder|false|false||URINE Bloodnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|nitrite ion|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|Nitrites|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitrite
null|nitrite ion|Drug|false|false||Nitritenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Proteins|Drug|false|false||Protein
null|Proteins|Drug|false|false||Proteinnull|Protein Info|Finding|false|false||Proteinnull|Protein measurement|Procedure|false|false||Proteinnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Ketones|Drug|false|false||Ketonenull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|Neg - answer|Finding|false|false||NEGnull|Negative - qualifier|Modifier|false|false||NEGnull|null|Lab|false|false|C0014792|URINE RBC
null|Red blood cells urine positive|Lab|false|false|C0014792|URINE RBCnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0221752;C2188659;C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Leukocytes|Anatomy|false|false||WBCnull|Yeast, Dried|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeast
null|Candida albicans allergenic extract|Drug|false|false||Yeastnull|Saccharomyces cerevisiae|Entity|false|false||Yeast
null|Yeasts|Entity|false|false||Yeastnull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|Mucus in urine (finding)|Finding|false|false||URINE Mucousnull|Portion of urine|Finding|false|false||URINE
null|null|Finding|false|false||URINE
null|Urine|Finding|false|false||URINE
null|In Urine|Finding|false|false||URINE
null|Urine specimen|Finding|false|false||URINEnull|Mucus (substance)|Finding|false|false||Mucous
null|mucus layer|Finding|false|false||Mucousnull|Mucous appearance|Modifier|false|false||Mucousnull|Retinoic Acid Response Element|Finding|false|false||RAREnull|Infrequent|Time|false|false||RAREnull|Rare|Modifier|false|false||RAREnull|Parameterized Data Type - Interval|Finding|false|false||INTERVALnull|Interval|Time|false|false||INTERVALnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C0004002;C0242192;C1121182;C2257651;C1415274;C1140170;C4553172;C0202113;C0851148;C4522245;C1266129;C1370889;C1415181;C1420113;C5960784|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Lactate Dehydrogenase|Drug|false|false||LDH
null|Lactate Dehydrogenase|Drug|false|false||LDHnull|Lifetime Drinking History|Finding|false|false|C1185650|LDHnull|Lactate dehydrogenase measurement|Procedure|false|false|C1185650|LDHnull|Alkaline Phosphatase|Drug|false|false||AlkPhos
null|Alkaline Phosphatase|Drug|false|false||AlkPhosnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Mandibular left third molar abutment mesial hemisection|Device|false|false||17AMnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|C-Reactive Protein, human|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-Reactive Protein, human|Drug|false|false||CRPnull|CRP wt Allele|Finding|false|false||CRP
null|CRP gene|Finding|false|false||CRP
null|CSRP1 gene|Finding|false|false||CRP
null|PPIAP10 gene|Finding|false|false||CRPnull|Pidgin and Creole language|Entity|false|false||CRPnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Structure of left foot|Anatomy|false|false|C0043299;C1552822;C0043309;C0555980|LEFT FOOTnull|Table Cell Horizontal Align - left|Finding|false|false|C4299097;C0016504;C0230461|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|FOOTnull|Lower extremity>Foot|Anatomy|false|false|C1552822;C0555980;C0043309;C0043299|FOOT
null|Foot|Anatomy|false|false|C1552822;C0555980;C0043309;C0043299|FOOTnull|Foot Unit of Length|LabModifier|false|false||FOOTnull|Diagnostic radiologic examination|Procedure|false|false|C0230461;C4299097;C0016504|XRAYnull|Roentgen Rays|Phenomenon|false|false|C4299097;C0016504;C0230461|XRAYnull|Ulceration|Finding|false|false||ulceration
null|Ulcer|Finding|false|false||ulcerationnull|Medial|Modifier|false|false||medialnull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Aspect (characteristic)|Modifier|false|false||aspectnull|Aspect - Kind of quantity|LabModifier|false|false||aspectnull|Hallux structure|Anatomy|false|false|C1424898|great toenull|RXFP2 gene|Finding|false|false|C0018534;C0040357;C4299090|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C1424898|toe
null|Toes|Anatomy|false|false|C1424898|toenull|Superficial ulcer|Disorder|false|false|C0576464;C3669027;C0223792;C0222682;C2987514|erosionnull|Erosion lesion|Finding|false|false|C0223792;C0222682;C2987514;C0576464;C3669027|erosionnull|Medial|Modifier|false|false||medialnull|nitrogenous base|Drug|false|false|C2987514|base
null|Base|Drug|false|false|C2987514|base
null|Dental Base|Drug|false|false|C2987514|base
null|base - RoleClass|Drug|false|false|C2987514|basenull|Base - General Qualifier|Finding|false|false|C2987514;C0576464;C3669027;C0223792;C0222682|base
null|BPIFA4P gene|Finding|false|false|C2987514;C0576464;C3669027;C0223792;C0222682|base
null|Base - RX Component Type|Finding|false|false|C2987514;C0576464;C3669027;C0223792;C0222682|basenull|Anatomical base|Anatomy|false|false|C1704464;C0178499;C1550601;C1880279;C1549548;C1705938;C1843354;C1959609;C0333307|basenull|Base - unit of product usage|LabModifier|false|false||basenull|Bone structure of distal phalanx|Anatomy|false|false|C0333307;C1549548;C1705938;C1843354;C1959609|distal phalanx
null|null|Anatomy|false|false|C0333307;C1549548;C1705938;C1843354;C1959609|distal phalanxnull|Distal Resection Margin|Attribute|false|false|C0223792;C0222682|distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Phalanx of hand|Anatomy|false|false|C1959609;C1549548;C1705938;C1843354;C4522154;C0333307|phalanx
null|Phalanx structure|Anatomy|false|false|C1959609;C1549548;C1705938;C1843354;C4522154;C0333307|phalanxnull|Hallux structure|Anatomy|false|false|C1424898|great toenull|RXFP2 gene|Finding|false|false|C0040357;C4299090;C0018534|greatnull|Greater|LabModifier|false|false||great
null|Large|LabModifier|false|false||greatnull|Lower extremity>Toes|Anatomy|false|false|C1424898|toe
null|Toes|Anatomy|false|false|C1424898|toenull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Parameterized Data Type - Interval|Finding|false|false||intervalnull|Interval|Time|false|false||intervalnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|MRI with contrast|Procedure|false|false||MRI with contrastnull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Contrast Media|Drug|false|false||contrastnull|Contrast|Modifier|false|false||contrastnull|Further|Modifier|false|false||furthernull|Knowledge acquisition using a method of assessment|Finding|false|false||assessmentnull|assessment of cognitive functions|Procedure|false|false||assessment
null|Physical Examination|Procedure|false|false||assessment
null|Nutrition Assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Personal care assessment|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|Evaluation procedure|Procedure|false|false||assessment
null|Evaluation|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessment
null|null|Procedure|false|false||assessmentnull|Assessed|Event|false|false||assessmentnull|Nias Language|Entity|false|false||NIASnull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|Triphasic|Time|false|false||triphasicnull|Doppler studies|Procedure|false|false||Dopplernull|Waveforms|Phenomenon|false|false||waveformsnull|Table Cell Horizontal Align - right|Finding|false|false|C0015811|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Femur|Anatomy|false|false|C1552823|femoralnull|popliteal|Anatomy|false|false|C0397581|poplitealnull|Procedure on artery|Procedure|false|false|C0442037;C0226004;C0003842|arteriesnull|Arteries|Anatomy|false|false|C0397581|arteries
null|Arterial system|Anatomy|false|false|C0397581|arteriesnull|Absent|Finding|false|false||Absentnull|Expression Negative|Lab|false|false||Absentnull|Waveforms|Phenomenon|false|false||waveformnull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Tibial Arteries|Anatomy|false|false||tibial arterynull|Bone structure of tibia|Anatomy|false|false||tibialnull|Arterial system|Anatomy|false|false||artery
null|Arteries|Anatomy|false|false||arterynull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|null|Attribute|false|false||ABI
null|Ankle brachial pressure index (observable entity)|Attribute|false|false||ABInull|Blood Vessel|Anatomy|false|false||vesselsnull|LEFT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE LEFT SIDE OF THE BODY)|Modifier|false|false||left side
null|Left|Modifier|false|false||left sidenull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Side|Modifier|false|false||sidenull|Triphasic|Time|false|false||triphasicnull|Doppler studies|Procedure|false|false||Dopplernull|Waveforms|Phenomenon|false|false||waveformsnull|Table Cell Horizontal Align - left|Finding|false|false|C0015811|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Femur|Anatomy|false|false|C1552822|femoralnull|Structure of popliteal artery|Anatomy|false|false|C0397581|popliteal arteriesnull|popliteal|Anatomy|false|false|C0397581|poplitealnull|Procedure on artery|Procedure|false|false|C0442037;C0226004;C0003842;C0032649|arteriesnull|Arteries|Anatomy|false|false|C0397581|arteries
null|Arterial system|Anatomy|false|false|C0397581|arteriesnull|Monophasic|Time|false|false||Monophasicnull|Waveforms|Phenomenon|false|false||waveformsnull|Posterior pituitary disease|Disorder|false|false|C0040184|posteriornull|Dorsal|Modifier|false|false||posteriornull|Bone structure of tibia|Anatomy|false|false|C0751438|tibialnull|Procedure on artery|Procedure|false|false|C0226004;C0003842|arteriesnull|Arteries|Anatomy|false|false|C0397581|arteries
null|Arterial system|Anatomy|false|false|C0397581|arteriesnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|null|Attribute|false|false||ABI
null|Ankle brachial pressure index (observable entity)|Attribute|false|false||ABInull|Pulse volume|Finding|false|false||Pulse volumenull|Physiologic pulse|Finding|false|false||Pulsenull|Pulse taking|Procedure|false|false||Pulsenull|Pulse Rate|Attribute|false|false||Pulsenull|Pulse phenomenon|Phenomenon|false|false||Pulsenull|Volume (publication)|Finding|false|false||volumenull|Volume|LabModifier|false|false||volumenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Structure of calf of leg|Anatomy|false|false||calf
null|null|Anatomy|false|false||calfnull|Cattle calf (organism)|Entity|false|false||calfnull|Lower extremity>Ankle|Anatomy|false|false||ankle
null|Ankle|Anatomy|false|false||ankle
null|Ankle joint structure|Anatomy|false|false||anklenull|Metatarsal bone structure|Anatomy|false|false||metatarsalnull|Significant|Finding|false|false||Significantnull|Event Seriousness - Significant|Modifier|false|false||Significantnull|Bilateral|Modifier|false|false||bilateralnull|Bone structure of tibia|Anatomy|false|false|C0003834|tibialnull|Arterial insufficiency|Disorder|false|false|C0003842;C0040184|arterial insufficiencynull|Arteries|Anatomy|false|false|C0003834|arterialnull|Arterial|Modifier|false|false||arterialnull|Insufficiency|Finding|false|false||insufficiencynull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|At rest (qualifier value)|Finding|false|false||at restnull|REST protein, human|Drug|false|false||rest
null|REST protein, human|Drug|false|false||restnull|REST gene|Finding|false|false||rest
null|site-specific telomere resolvase activity|Finding|false|false||rest
null|Rest|Finding|false|false||restnull|More|LabModifier|false|false||morenull|Significant|Finding|false|false||significantnull|Event Seriousness - Significant|Modifier|false|false||significantnull|RIGHT SIDE (USED TO IDENTIFY PROCEDURES PERFORMED ON THE RIGHT SIDE OF THE BODY)|Modifier|false|false||right side
null|Right|Modifier|false|false||right sidenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Side|Modifier|false|false||sidenull|Plain chest X-ray|Procedure|false|false||CXRnull|Comparison|Event|false|false||Comparisonnull|Relevance|Modifier|false|false||relevantnull|Changing|Finding|true|false||changenull|Change - procedure|Procedure|true|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Alignment|Modifier|false|false||Alignmentnull|Wiring of sternum|Procedure|false|false|C0038293|sternal wiresnull|Sternum|Anatomy|false|false|C0407260|sternalnull|Bone Wires|Device|false|false||wiresnull|null|Modifier|false|false||unremarkablenull|Mild Severity of Illness Code|Finding|false|false||Mildnull|Mild (qualifier value)|Modifier|false|false||Mild
null|Mild Allergy Severity|Modifier|false|false||Mildnull|Descending aorta|Anatomy|false|false|C1547177;C0869784|descending aorta
null|null|Anatomy|false|false|C1547177;C0869784|descending aortanull|Sequencing - Descending|Finding|false|false|C4037978;C0003483;C1305624;C0011666|descendingnull|Descending|Modifier|false|false||descendingnull|Procedure on aorta|Procedure|false|false|C4037978;C0003483;C1305624;C0011666|aortanull|Chest+Abdomen>Aorta|Anatomy|false|false|C1547177;C0869784|aorta
null|Aorta|Anatomy|false|false|C1547177;C0869784|aortanull|Borderline|Modifier|false|false||Borderlinenull|size|Modifier|false|false||sizenull|size - solid dosage form|LabModifier|false|false||sizenull|Malignant neoplasm of heart|Disorder|false|false|C4037974;C0018787|heart
null|benign neoplasm of heart|Disorder|false|false|C4037974;C0018787|heartnull|HEART PROBLEM|Finding|false|false|C4037974;C0018787|heartnull|Chest>Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heart
null|Heart|Anatomy|false|false|C0795691;C0153957;C0153500|heartnull|Pleural effusion (disorder)|Finding|true|false|C0032225|pleural effusionsnull|Pleural Diseases|Disorder|false|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0032226;C0032227;C0013687|pleuralnull|Pleural|Modifier|false|false||pleuralnull|effusion|Finding|true|false|C0032225|effusionsnull|Pneumonia|Disorder|false|false||pneumonianull|Pulmonary Edema|Finding|false|false|C0024109|pulmonary edemanull|Pulmonary (intended site)|Finding|false|false|C0024109|pulmonarynull|Lung|Anatomy|false|false|C2707265;C0013604;C4522268;C0034063|pulmonarynull|null|Attribute|false|false|C0024109|pulmonarynull|Pulmonary (qualifier value)|Modifier|false|false||pulmonarynull|Edema|Finding|false|false|C0024109|edemanull|null|Attribute|false|false||edemanull|CYREN gene|Finding|false|false|C0230461|MRInull|Magnetic resonance imaging service|Procedure|false|false|C0230461|MRI
null|Magnetic Resonance Imaging|Procedure|false|false|C0230461|MRInull|Maori Language|Entity|false|false||MRInull|Structure of left foot|Anatomy|false|false|C1824234;C0024485;C0587658;C0555980;C1552822|LEFT FOOTnull|Table Cell Horizontal Align - left|Finding|false|false|C0230461|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Foot problem|Finding|false|false|C0230461;C4299097;C0016504|FOOTnull|Lower extremity>Foot|Anatomy|false|false|C0555980|FOOT
null|Foot|Anatomy|false|false|C0555980|FOOTnull|Foot Unit of Length|LabModifier|false|false||FOOTnull|Prostate Stromal Proliferation of Uncertain Malignant Potential|Disorder|false|false|C0225317;C4532079|stump
null|Atypical Spitz Nevus|Disorder|false|false|C0225317;C4532079|stump
null|Amputation Stumps|Disorder|false|false|C0225317;C4532079|stump
null|Neoplasm of uncertain behavior of smooth muscle|Disorder|false|false|C0225317;C4532079|stumpnull|Neck+Chest>Soft tissue|Anatomy|false|false|C3542022;C1547928;C4522245;C0002690;C5848682;C1514517|soft tissue
null|soft tissue|Anatomy|false|false|C3542022;C1547928;C4522245;C0002690;C5848682;C1514517|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0225317;C4532079|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0040300;C0225317;C4532079|tissuenull|Body tissue|Anatomy|false|false|C1547928|tissuenull|Plantar (qualifier value)|Anatomy|false|false|C0332568;C1704436;C3887682;C0812278;C1705088;C1708004;C1366645;C0279453|plantar
null|Sole of Foot|Anatomy|false|false|C0332568;C1704436;C3887682;C0812278;C1705088;C1708004;C1366645;C0279453|plantarnull|Fat pad|Anatomy|false|false|C3540603;C1425478;C1425244;C1435181;C0015677;C3887682;C3887682;C0812278;C1705088;C1708004;C1366645;C3814046;C0332568;C1704436;C0279453|fat padnull|Platelet Glycoprotein 4, human|Drug|false|false|C0935625;C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0935625;C0001527|fat
null|FAT1 protein, human|Drug|false|false|C0935625;C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0935625;C0001527|fat
null|Fatty acid glycerol esters|Drug|false|false|C0935625;C0001527|fatnull|Platelet Glycoprotein 4, human|Finding|false|false|C3669270;C0935625;C0001527;C0442036;C0230463|fat
null|CD36 gene|Finding|false|false|C3669270;C0935625;C0001527;C0442036;C0230463|fat
null|FAT1 gene|Finding|false|false|C3669270;C0935625;C0001527;C0442036;C0230463|fat
null|CD36 wt Allele|Finding|false|false|C3669270;C0935625;C0001527;C0442036;C0230463|fat
null|FAT1 wt Allele|Finding|false|false|C3669270;C0935625;C0001527;C0442036;C0230463|fatnull|doxorubicin/fluorouracil/triazinate protocol|Procedure|false|false|C0001527;C0935625;C0442036;C0230463;C3669270|fatnull|Adipose tissue|Anatomy|false|false|C3814046;C3540603;C1425478;C1425244;C3887682;C0812278;C1705088;C1708004;C1366645;C0332568;C1704436;C1435181;C0015677;C3887682;C0279453|fatnull|Obese build|Subject|false|false||fatnull|Fantse Language|Entity|false|false||fatnull|Pad Dosage Form|Drug|false|false|C3669270|padnull|Pad Mass|Disorder|false|false|C0442036;C0230463;C0935625;C0001527;C3669270|pad
null|Peripheral Arterial Diseases|Disorder|false|false|C0442036;C0230463;C0935625;C0001527;C3669270|padnull|PADI4 wt Allele|Finding|false|false|C0935625;C3669270;C0001527|pad
null|PADI4 gene|Finding|false|false|C0935625;C3669270;C0001527|pad
null|DHX40 gene|Finding|false|false|C0935625;C3669270;C0001527|padnull|PAD Regimen|Procedure|false|false|C0001527;C0935625;C3669270|padnull|Strucure of thick cushion of skin|Anatomy|false|false|C3887682;C0812278;C1705088;C1708004;C1366645;C3540603;C1425478;C1425244;C3814046;C0332568;C1704436;C2347441;C0279453|padnull|Pad Device|Device|false|false||pad
null|Pads|Device|false|false||padnull|Pad (unit of presentation)|LabModifier|false|false||pad
null|Pad Dosing Unit|LabModifier|false|false||padnull|Table Cell Vertical Align - middle|Finding|false|false||middlenull|Middle|Modifier|false|false||middle
null|Midline (qualifier value)|Modifier|false|false||middlenull|Phalanx structure|Anatomy|false|false|C1547928|phalanges
null|Phalanx of hand|Anatomy|false|false|C1547928|phalangesnull|Tissue Specimen Code|Finding|false|false|C0040300;C0223792;C0222682|tissuenull|Body tissue|Anatomy|false|false|C1547928|tissuenull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Abscess|Disorder|false|false||abscessnull|null|Finding|false|false||abscessnull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Signal|Phenomenon|false|false||signalnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Distal Resection Margin|Attribute|false|false||distalnull|Distal (qualifier value)|Modifier|false|false||distalnull|Adrenal Cortex Diseases|Disorder|false|false|C1176472;C0007776|cortex
null|cortex bone disorders|Disorder|false|false|C1176472;C0007776|cortexnull|Cortex of Organ|Anatomy|false|false|C0001614;C0595905|cortex
null|Cerebral cortex|Anatomy|false|false|C0001614;C0595905|cortexnull|Bark - plant part|Entity|false|false||cortexnull|First metatarsal structure|Anatomy|false|false||first metatarsalnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Metatarsal bone structure|Anatomy|false|false||metatarsalnull|Comparison study|Procedure|false|false||comparison study
null|comparative study research|Procedure|false|false||comparison studynull|Comparison|Event|false|false||comparisonnull|Study Object|Finding|false|false||studynull|Scientific Study|Procedure|false|false||study
null|Study|Procedure|false|false||study
null|Clinical Research|Procedure|false|false||studynull|Room of building - Study|Device|false|false||studynull|Has focus|Finding|false|false||focusnull|Focal|Modifier|false|false||focusnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|Inflammatory fistula|Finding|false|false|C1185740;C1305231;C0030471;C0018670;C0152336;C0025584;C0459701|sinus tractsnull|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinus
null|Sinus brand of acetaminophen-pseudoephedrine|Drug|false|false|C1305231;C0030471|sinusnull|pathologic fistula|Disorder|false|false|C0025584;C1305231;C0030471;C0459701;C1185740|sinusnull|Sinus - general anatomical term|Anatomy|false|false|C0723346;C0544791;C0016169|sinus
null|Nasal sinus|Anatomy|false|false|C0723346;C0544791;C0016169|sinusnull|Tract|Anatomy|false|false|C0544791;C0016169|tractsnull|Medial|Modifier|false|false||medialnull|Problems with head|Disorder|false|false|C0018670;C0152336;C0025584;C0459701|headnull|Procedure on head|Procedure|false|false|C0025584;C0018670;C0152336;C0459701|headnull|Structure of head of caudate nucleus|Anatomy|false|false|C0362076;C0876917;C0544791|head
null|Head|Anatomy|false|false|C0362076;C0876917;C0544791|headnull|Head Device|Device|false|false||headnull|First metatarsal structure|Anatomy|false|false|C0876917;C0016169;C0544791;C0362076|first metatarsalnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Metatarsal bone structure|Anatomy|false|false|C0876917;C0016169;C0544791;C0362076|metatarsalnull|Status post|Time|false|false||status post
null|Post|Time|false|false||status postnull|What subject filter - Status|Finding|false|false||statusnull|null|Attribute|false|false||statusnull|Social status|Modifier|false|false||status
null|Status|Modifier|false|false||statusnull|SLC35G1 gene|Finding|false|false||post
null|DESI1 gene|Finding|false|false||postnull|Post Device|Device|false|false||postnull|Post|Time|false|false||postnull|Amputated structure (morphologic abnormality)|Disorder|false|false||amputationnull|Amputation Specimen Code|Finding|false|false||amputationnull|Amputation|Procedure|false|false||amputationnull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|maltose tetrapalmitate|Drug|false|false||MTP
null|maltose tetrapalmitate|Drug|false|false||MTPnull|MTTP wt Allele|Finding|false|false||MTP
null|MTTP gene|Finding|false|false||MTPnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Dorsal|Modifier|false|false||Dorsalnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Diffuse|Modifier|false|false||diffusenull|Edematous skin|Finding|false|false|C1123023;C4520765|skin edemanull|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0521464;C0013604;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0521464;C0013604;C0178298;C0496955|skinnull|Edema|Finding|false|false|C1123023;C4520765|edemanull|null|Attribute|false|false||edemanull|Plain chest X-ray|Procedure|false|false||CXRnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICC PLACEMENTnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|null|Procedure|false|false||PLACEMENT
null|Implantation procedure|Procedure|false|false||PLACEMENT
null|Clinical act of insertion|Procedure|false|false||PLACEMENTnull|Placement|Modifier|false|false||PLACEMENTnull|Query Status Code - new|Finding|false|false||New
null|Act Status - new|Finding|false|false||Newnull|Newar Language|Entity|false|false||Newnull|New|Modifier|false|false||Newnull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false||PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|KAT5 wt Allele|Finding|false|false||tip
null|ITFG1 gene|Finding|false|false||tip
null|METTL8 gene|Finding|false|false||tip
null|TIPRL gene|Finding|false|false||tipnull|TIP regimen|Procedure|false|false||tipnull|Device tip (physical object)|Device|false|false||tipnull|Tip|Modifier|false|false||tipnull|Junction Device|Device|false|false||junctionnull|Junctional|Modifier|false|false||junctionnull|Superior vena cava structure|Anatomy|false|false|C1413046|superior vena cava
null|Chest>Vena cava.superior|Anatomy|false|false|C1413046|superior vena cavanull|Upper|Modifier|false|false||superiornull|Chest+Abdomen>Vena cava.superior &or Vena cava.inferior|Anatomy|false|false|C1413046|vena cava
null|Vena caval structure|Anatomy|false|false|C1413046|vena cavanull|Structure of vein of trunk|Anatomy|false|false|C1413046|venanull|CA5A gene|Finding|false|false|C0447122;C0042459;C4266604;C4266402;C0042460|cavanull|Right atrial structure|Anatomy|false|false|C1552823|right atriumnull|Table Cell Horizontal Align - right|Finding|false|false|C0018792;C0225844|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Heart Atrium|Anatomy|false|false|C1552823|atriumnull|Pneumothorax|Disorder|true|false||pneumothoraxnull|Remote control command - Clear|Finding|false|false|C0024109|Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Lung|Anatomy|false|false|C1550016|lungsnull|Pathology processes|Finding|false|false||PATHOLOGY
null|Pathological aspects|Finding|false|false||PATHOLOGYnull|Pathology procedure|Procedure|false|false||PATHOLOGYnull|Pathology|Title|false|false||PATHOLOGYnull|Operative Surgical Procedures|Procedure|false|false|C0040300|SURGICAL
null|Surgical service|Procedure|false|false|C0040300|SURGICALnull|Tissue Specimen Code|Finding|false|false|C0040300|TISSUEnull|Body tissue|Anatomy|false|false|C0543467;C0587668;C1547928|TISSUEnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|Bone
null|null|Finding|false|false|C1442209;C0262950|Bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616;C1547296;C0332290;C0392747;C1555457;C0332290|Bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616;C1547296;C0332290;C0392747;C1555457;C0332290|Bonenull|Changing|Finding|false|false|C1442209;C0262950|changesnull|Changed status|LabModifier|false|false||changesnull|Consistent with|Finding|false|false|C1442209;C0262950|consistent withnull|Compatible|Modifier|false|false||consistent withnull|Consistent with|Finding|false|false|C1442209;C0262950|consistentnull|Chronic - Admission Level of Care Code|Finding|false|false|C1442209;C0262950|chronicnull|Provision of recurring care for chronic illness|Procedure|false|false|C1442209;C0262950|chronicnull|chronic|Time|false|false||chronicnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Acute osteomyelitis|Disorder|true|false||acute osteomyelitisnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Osteomyelitis|Disorder|true|false||osteomyelitisnull|Operative Surgical Procedures|Procedure|false|false|C0040300|SURGICAL
null|Surgical service|Procedure|false|false|C0040300|SURGICALnull|Tissue Specimen Code|Finding|false|false|C0040300|TISSUEnull|Body tissue|Anatomy|false|false|C1547928;C0543467;C0587668|TISSUEnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Hallux structure|Anatomy|false|false|C1552822;C0015252;C0728940;C1424898|GREAT TOEnull|RXFP2 gene|Finding|false|false|C0040357;C4299090;C0018534|GREATnull|Greater|LabModifier|false|false||GREAT
null|Large|LabModifier|false|false||GREATnull|Lower extremity>Toes|Anatomy|false|false|C0015252;C0728940;C1424898|TOE
null|Toes|Anatomy|false|false|C0015252;C0728940;C1424898|TOEnull|Excision|Procedure|false|false|C0040357;C4299090;C0018534|EXCISION
null|removal technique|Procedure|false|false|C0040357;C4299090;C0018534|EXCISIONnull|Acute osteomyelitis|Disorder|false|false||Acute osteomyelitisnull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|Focal|Modifier|false|false||focalnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|Bone
null|null|Finding|false|false|C1442209;C0262950|Bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bonenull|Changing|Finding|false|false|C1442209;C0262950|changesnull|Changed status|LabModifier|false|false||changesnull|Skin and subcutaneous tissue disorders|Disorder|false|false|C0222331;C0278403;C1123023;C4520765|Skin
null|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C0222331;C0278403;C1123023;C4520765|Skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765;C0222331;C0278403|Skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765;C0222331;C0278403|Skinnull|Skin, Human|Anatomy|false|false|C0333361;C3887532;C0041582;C0021368;C0178298;C0496955;C1546781;C0444099;C1547295;C1547229|Skin
null|Skin|Anatomy|false|false|C0333361;C3887532;C0041582;C0021368;C0178298;C0496955;C1546781;C0444099;C1547295;C1547229|Skinnull|Subcutaneous Tissue|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|subcutis
null|Subcutaneous Fat|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099|subcutisnull|Ulceration|Finding|false|false|C1123023;C4520765|ulceration
null|Ulcer|Finding|false|false|C1123023;C4520765|ulcerationnull|Acute inflammation|Finding|false|false|C1123023;C4520765|acute inflammationnull|Admission Level of Care Code - Acute|Finding|false|false|C1123023;C4520765|acute
null|Acute - Triage Code|Finding|false|false|C1123023;C4520765|acutenull|acute|Time|false|false||acutenull|Inflammation|Finding|false|false|C1123023;C4520765|inflammationnull|Atherosclerosis|Disorder|false|false||Atherosclerosis
null|Arteriosclerosis|Disorder|false|false||Atherosclerosisnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Bone structure of proximal phalanx|Anatomy|false|false|C1549548;C1705938;C1843354;C1552822;C4489236;C4761388|PROXIMAL PHALANX
null|null|Anatomy|false|false|C1549548;C1705938;C1843354;C1552822;C4489236;C4761388|PROXIMAL PHALANXnull|Proximal Resection Margin|Attribute|false|false|C0576462;C3669035|PROXIMALnull|Proximal|Modifier|false|false||PROXIMALnull|Phalanx structure|Anatomy|false|false|C4761388;C1549548;C1705938;C1843354|PHALANX
null|Phalanx of hand|Anatomy|false|false|C4761388;C1549548;C1705938;C1843354|PHALANXnull|nitrogenous base|Drug|false|false|C2987514|BASE
null|Base|Drug|false|false|C2987514|BASE
null|Dental Base|Drug|false|false|C2987514|BASE
null|base - RoleClass|Drug|false|false|C2987514|BASEnull|Base - General Qualifier|Finding|false|false|C0576462;C3669035;C2987514;C0223792;C0222682|BASE
null|BPIFA4P gene|Finding|false|false|C0576462;C3669035;C2987514;C0223792;C0222682|BASE
null|Base - RX Component Type|Finding|false|false|C0576462;C3669035;C2987514;C0223792;C0222682|BASEnull|Anatomical base|Anatomy|false|false|C1549548;C1705938;C1843354;C4761388;C1704464;C0178499;C1550601;C1880279|BASEnull|Base - unit of product usage|LabModifier|false|false||BASEnull|null|Finding|false|false|C0223792;C0222682;C0576462;C3669035;C2987514|MARGINnull|Marginal|Modifier|false|false||MARGINnull|Table Cell Horizontal Align - left|Finding|false|false|C0576462;C3669035|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Excision|Procedure|false|false||EXCISION
null|removal technique|Procedure|false|false||EXCISIONnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|Bone
null|null|Finding|false|false|C1442209;C0262950|Bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bonenull|Changing|Finding|false|false|C1442209;C0262950|changesnull|Changed status|LabModifier|false|false||changesnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Acute osteomyelitis|Disorder|true|false||acute osteomyelitisnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Osteomyelitis|Disorder|true|false||osteomyelitisnull|Bone structure of proximal phalanx|Anatomy|false|false|C1552822;C0015252;C0728940|PROXIMAL PHALANX
null|null|Anatomy|false|false|C1552822;C0015252;C0728940|PROXIMAL PHALANXnull|Proximal Resection Margin|Attribute|false|false||PROXIMALnull|Proximal|Modifier|false|false||PROXIMALnull|Phalanx structure|Anatomy|false|false||PHALANX
null|Phalanx of hand|Anatomy|false|false||PHALANXnull|Table Cell Horizontal Align - left|Finding|false|false|C0576462;C3669035|LEFTnull|Left sided|Modifier|false|false||LEFT
null|Left|Modifier|false|false||LEFTnull|Excision|Procedure|false|false|C0576462;C3669035|EXCISION
null|removal technique|Procedure|false|false|C0576462;C3669035|EXCISIONnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|Bone
null|null|Finding|false|false|C1442209;C0262950|Bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616;C0392747|Bonenull|Changing|Finding|false|false|C1442209;C0262950|changesnull|Changed status|LabModifier|false|false||changesnull|Evidence of (contextual qualifier)|Finding|true|false||evidence ofnull|Evidence|Finding|true|false||evidencenull|Acute osteomyelitis|Disorder|true|false||acute osteomyelitisnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Osteomyelitis|Disorder|true|false||osteomyelitisnull|Microbiology Diagnostic Service Section ID|Finding|false|false||MICROBIOLOGY
null|Microbiological|Finding|false|false||MICROBIOLOGY
null|Microbiology - Laboratory Class|Finding|false|false||MICROBIOLOGYnull|Microbiology procedure|Procedure|false|false||MICROBIOLOGYnull|Science of Microbiology|Title|false|false||MICROBIOLOGYnull|Tissue Specimen Code|Finding|false|false|C0040300|TISSUEnull|Body tissue|Anatomy|false|false|C1547928|TISSUEnull|Proximal Resection Margin|Attribute|false|false||PROXIMALnull|Proximal|Modifier|false|false||PROXIMALnull|Gram's stain|Drug|false|false||GRAM STAIN
null|Gram's stain|Drug|false|false||GRAM STAINnull|Bacterial stain, routine|Procedure|false|false||GRAM STAINnull|gram|LabModifier|false|false||GRAMnull|Stains|Drug|false|false||STAINnull|Staining method|Procedure|false|false||STAINnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Specimen Type - Leukocytes|Finding|false|false|C0023516|LEUKOCYTES
null|null|Finding|false|false|C0023516|LEUKOCYTESnull|Leukocytes|Anatomy|false|false|C1550647;C1547962|LEUKOCYTESnull|Knowledge Field|Finding|false|false||FIELD
null|Force Field|Finding|false|false||FIELD
null|Field|Finding|false|false||FIELDnull|field - patient encounter|Procedure|false|false||FIELDnull|Gram-Positive Cocci|Entity|false|false||GRAM POSITIVE COCCInull|gram|LabModifier|false|false||GRAMnull|BRAF Gene Rearrangement|Disorder|false|false||POSITIVEnull|Rh Positive Blood Group|Finding|false|false||POSITIVE
null|Positive Finding|Finding|false|false||POSITIVE
null|Positive|Finding|false|false||POSITIVEnull|Positive Charge|Modifier|false|false||POSITIVEnull|Positive Number|LabModifier|false|false||POSITIVEnull|Cocci bacteria|Entity|false|false||COCCInull|Mandibular left second premolar mesial prosthesis|Device|false|false||20PMnull|Tissue Specimen Code|Finding|false|false|C0040300|TISSUEnull|Body tissue|Anatomy|false|false|C1547928;C1546485|TISSUEnull|Diagnosis Type - Final|Finding|false|false|C0040300|Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Staphylococcus aureus|Entity|false|false||STAPH AUREUSnull|Staphylococcal Infections|Disorder|false|false||STAPHnull|Genus staphylococcus|Entity|false|false||STAPHnull|Blood coagulation tests|Procedure|false|false||COAGnull|Growth & development aspects|Finding|false|false||GROWTH
null|Tissue Growth|Finding|false|false||GROWTH
null|Growth|Finding|false|false||GROWTH
null|growth aspects|Finding|false|false||GROWTHnull|Growth action|Phenomenon|false|false||GROWTHnull|Microbial susceptibility tests|Procedure|false|false||Susceptibility testingnull|Susceptibility (property) (qualifier value)|Finding|false|false||Susceptibilitynull|Disease susceptibility|Attribute|false|false||Susceptibilitynull|null|Subject|false|false||Susceptibilitynull|Testing|Finding|false|false||testing
null|Tests (qualifier value)|Finding|false|false||testingnull|Culture Dose Form|Drug|false|false||culturenull|Culture (Anthropological)|Finding|false|false||culture
null|Cultural aspects|Finding|false|false||culturenull|Microbial culture (procedure)|Procedure|false|false||culture
null|Laboratory culture|Procedure|false|false||culturenull|Anaerobic microbial culture|Procedure|false|false||ANAEROBIC CULTUREnull|Anaerobic|Modifier|false|false||ANAEROBICnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Bacteria, Anaerobic|Entity|true|false||ANAEROBESnull|Acid fast stain|Drug|false|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|false|false||FAST
null|FASTK Gene|Finding|false|false||FAST
null|FOXD3-AS1 gene|Finding|false|false||FAST
null|FASTK wt Allele|Finding|false|false||FAST
null|Fasting|Finding|false|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Acid fast stain|Drug|true|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|true|false||FAST
null|FASTK Gene|Finding|true|false||FAST
null|FOXD3-AS1 gene|Finding|true|false||FAST
null|FASTK wt Allele|Finding|true|false||FAST
null|Fasting|Finding|true|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Bacilli <Bacillota>|Entity|true|false||BACILLI
null|Genus Bacillus|Entity|true|false||BACILLInull|Direct - PostalAddressUse|Finding|false|false||DIRECT
null|direct address|Finding|false|false||DIRECTnull|Direct type of relationship|Modifier|false|false||DIRECT
null|Direct (qualifier)|Modifier|false|false||DIRECTnull|Smearing technique|Finding|false|false||SMEARnull|Smear test|Procedure|false|false||SMEARnull|Smear - instruction imperative|Event|false|false||SMEARnull|Acid fast stain|Drug|false|false||ACID FASTnull|Fas-activated serine/threonine kinase activity|Finding|false|false||FAST
null|FASTK Gene|Finding|false|false||FAST
null|FOXD3-AS1 gene|Finding|false|false||FAST
null|FASTK wt Allele|Finding|false|false||FAST
null|Fasting|Finding|false|false||FASTnull|Rapid|Modifier|false|false||FASTnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Preliminary|Time|false|false||Preliminarynull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|Blood culture|Procedure|false|false||BLOOD CULTUREnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Culture Dose Form|Drug|false|false||CULTUREnull|Culture (Anthropological)|Finding|false|false||CULTURE
null|Cultural aspects|Finding|false|false||CULTUREnull|Microbial culture (procedure)|Procedure|false|false||CULTURE
null|Laboratory culture|Procedure|false|false||CULTUREnull|Final report|Finding|false|false||FINAL REPORTnull|Diagnosis Type - Final|Finding|false|false||FINALnull|Final|Time|false|false||FINALnull|End-stage|Modifier|false|false||FINALnull|Report (document)|Finding|false|false||REPORTnull|Reporting|Procedure|false|false||REPORTnull|null|Attribute|false|false||REPORTnull|Blood culture|Procedure|false|false||Blood Culturenull|Blood and lymphatic system disorders|Disorder|false|false||Bloodnull|peripheral blood|Finding|false|false||Blood
null|Blood|Finding|false|false||Blood
null|In Blood|Finding|false|false||Bloodnull|Culture Dose Form|Drug|false|false||Culturenull|Culture (Anthropological)|Finding|false|false||Culture
null|Cultural aspects|Finding|false|false||Culturenull|Microbial culture (procedure)|Procedure|false|false||Culture
null|Laboratory culture|Procedure|false|false||Culturenull|Extended Priority Codes - Routine|Finding|false|false||Routine
null|Report priority - Routine|Finding|false|false||Routine
null|Admission Type - Routine|Finding|false|false||Routine
null|Level of Care - Routine|Finding|false|false||Routine
null|Processing priority - Routine|Finding|false|false||Routine
null|Referral priority - Routine|Finding|false|false||Routinenull|Routine coag|Procedure|false|false||Routinenull|Priority - Routine|Time|false|false||Routinenull|Routine|Modifier|false|false||Routinenull|Diagnosis Type - Final|Finding|false|false||Finalnull|Final|Time|false|false||Finalnull|End-stage|Modifier|false|false||Finalnull|Growth & development aspects|Finding|true|false||GROWTH
null|Tissue Growth|Finding|true|false||GROWTH
null|Growth|Finding|true|false||GROWTH
null|growth aspects|Finding|true|false||GROWTHnull|Growth action|Phenomenon|true|false||GROWTHnull|summary - ActRelationshipSubset|Finding|false|false||SUMMARY
null|Summary (document)|Finding|false|false||SUMMARYnull|Hypertensive disease|Disorder|false|false||HTNnull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false||diabeticnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0206172;C0555980|foot
null|Foot|Anatomy|false|false|C0206172;C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false||ulcer
null|null|Finding|false|false||ulcer
null|Ulcer|Finding|false|false||ulcernull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C1552822;C0029443|halluxnull|Osteomyelitis|Disorder|false|false|C0018534|osteomyelitisnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Sterile maggot wound debridement|Procedure|false|false||debridement
null|Debridement|Procedure|false|false||debridementnull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Tissue Specimen Code|Finding|false|false|C0040300|tissuenull|Body tissue|Anatomy|false|false|C1547928|tissuenull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|bone
null|null|Finding|false|false|C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|removal technique|Procedure|false|false||removal
null|Excision|Procedure|false|false||removal
null|Extraction|Procedure|false|false||removalnull|Removing (action)|Event|false|false||removalnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C0332840;C0002688;C1546539|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|On IV|Finding|false|false||on IVnull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|Finding|false|false||MSSAnull|Methicillin susceptible Staphylococcus aureus|Entity|false|false||MSSAnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Continuous|Finding|false|false||continuenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Infusion procedures|Procedure|false|false||infusionsnull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Osteomyelitis|Disorder|false|false|C0018534|Osteomyelitisnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C0029443|halluxnull|Skin ulcer due to diabetes mellitus|Disorder|false|false||diabetic ulcernull|Diabetic|Finding|false|false||diabeticnull|Specimen Type - Ulcer|Finding|false|false||ulcer
null|null|Finding|false|false||ulcer
null|Ulcer|Finding|false|false||ulcernull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false||halluxnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Target Awareness - partial|Finding|false|false||partialnull|Partial|LabModifier|false|false||partialnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C0002688;C0332840;C1552822;C1546539|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|Podiatry (discipline)|Title|false|false||podiatrynull|Initially|Time|false|false||initiallynull|On IV|Finding|false|false||on IVnull|vancomycin|Drug|false|false||Vancomycin
null|vancomycin|Drug|false|false||Vancomycinnull|Vancomycin measurement|Procedure|false|false||Vancomycinnull|Flagyl|Drug|false|false||Flagyl
null|Flagyl|Drug|false|false||Flagylnull|cefepime|Drug|false|false||cefepime
null|cefepime|Drug|false|false||cefepimenull|Initial (abbreviation)|Finding|false|false||Initialnull|Initially|Time|false|false||Initialnull|Firstly|Modifier|false|false||Initialnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Culture (Anthropological)|Finding|false|false||culturesnull|Positive|Finding|false|false||positive fornull|BRAF Gene Rearrangement|Disorder|false|false||positivenull|Rh Positive Blood Group|Finding|false|false||positive
null|Positive Finding|Finding|false|false||positive
null|Positive|Finding|false|false||positivenull|Positive Charge|Modifier|false|false||positivenull|Positive Number|LabModifier|false|false||positivenull|Encounter due to being carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|Finding|false|false||MSSAnull|Methicillin susceptible Staphylococcus aureus|Entity|false|false||MSSAnull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Apyrexial|Finding|false|false||afebrilenull|Structure of left foot|Anatomy|false|false|C0555980;C0041834|left footnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C0230461;C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0041834;C0555980|foot
null|Foot|Anatomy|false|false|C0041834;C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Erythema|Disorder|false|false|C4299097;C0016504;C0230461|erythemanull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Specimen Type - Ulcer|Finding|false|false||ulcer
null|null|Finding|false|false||ulcer
null|Ulcer|Finding|false|false||ulcernull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Concern|Finding|false|false||concernnull|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|false|false||poor
null|Patient Condition Code - Poor|Finding|false|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Specimen Type - Blood arterial|Finding|false|false|C0003842;C2335890|arterial blood
null|Arterial blood|Finding|false|false|C0003842;C2335890|arterial bloodnull|Portion of arterial blood|Anatomy|false|false|C0005775;C0232338;C1550611;C0229665|arterial bloodnull|Arteries|Anatomy|false|false|C1550611;C0229665;C0005768;C0229664;C0005767;C0851353;C0005775;C0232338|arterialnull|Arterial|Modifier|false|false||arterialnull|Blood flow|Finding|false|false|C2335890;C0003842|blood flow
null|Blood Circulation|Finding|false|false|C2335890;C0003842|blood flownull|Blood and lymphatic system disorders|Disorder|false|false|C0003842|bloodnull|peripheral blood|Finding|false|false|C0003842|blood
null|Blood|Finding|false|false|C0003842|blood
null|In Blood|Finding|false|false|C0003842|bloodnull|Flow|Phenomenon|false|false||flownull|Arteries|Anatomy|false|false|C2003888;C0947630|arterialnull|Arterial|Modifier|false|false||arterialnull|Scientific Study|Procedure|false|false|C0278454;C0015385;C0023216;C0003842|studiesnull|Bilateral|Modifier|false|false||bilateralnull|Lower Extremity|Anatomy|false|false|C2003888;C0947630|lower extremitiesnull|Body Site Modifier - Lower|Anatomy|false|false|C2003888|lowernull|Lower (action)|Event|false|false|C0003842;C0023216;C0278454;C0015385;C1548802|lowernull|Lower - spatial qualifier|Modifier|false|false||lowernull|All extremities|Anatomy|false|false|C0947630;C2003888|extremities
null|Limb structure|Anatomy|false|false|C0947630;C2003888|extremitiesnull|Scientific Study|Procedure|false|false||studiesnull|Mild Severity of Illness Code|Finding|false|false||mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|atherosclerotic|Finding|false|false||atheroscleroticnull|Disease|Disorder|false|false||diseasenull|Structure of left lower leg|Anatomy|false|false||left leg
null|Left lower extremity|Anatomy|false|false||left legnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Leg|Anatomy|false|false||leg
null|Lower Extremity|Anatomy|false|false||legnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980|foot
null|Foot|Anatomy|false|false|C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|atherosclerotic|Finding|false|false||atheroscleroticnull|Disease|Disorder|false|false|C0230442;C0230415|diseasenull|Structure of right lower leg|Anatomy|false|false|C1552823;C0012634;C0555980|right leg
null|Right lower extremity|Anatomy|false|false|C1552823;C0012634;C0555980|right legnull|Table Cell Horizontal Align - right|Finding|false|false|C0230442;C0230415|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Leg|Anatomy|false|false|C0555980|leg
null|Lower Extremity|Anatomy|false|false|C0555980|legnull|Foot problem|Finding|false|false|C0230442;C0230415;C1140621;C0023216;C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980|foot
null|Foot|Anatomy|false|false|C0555980|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Vascular Surgical Procedures|Procedure|false|false|C0005847|Vascular surgerynull|Vascular surgery specialty|Title|false|false||Vascular surgerynull|Blood Vessel|Anatomy|false|false|C0038895;C1457907;C1547138;C0543467;C0042381|Vascularnull|Vascular|Modifier|false|false||Vascularnull|Level of Care - Surgery|Finding|false|false|C0005847|surgery
null|Surgical procedure finding|Finding|false|false|C0005847|surgery
null|Surgical aspects|Finding|false|false|C0005847|surgerynull|Operative Surgical Procedures|Procedure|false|false|C0005847|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Potential|Modifier|false|false||potentialnull|Intervention regimes|Procedure|false|false||intervention
null|Nursing interventions|Procedure|false|false||intervention
null|Interventional procedure|Procedure|false|false||interventionnull|Further|Modifier|false|false||furthernull|Blood Vessel|Anatomy|false|false|C0886296;C0184661;C1273869|vascularnull|Vascular|Modifier|false|false||vascularnull|Intervention regimes|Procedure|true|false|C0005847|intervention
null|Nursing interventions|Procedure|true|false|C0005847|intervention
null|Interventional procedure|Procedure|true|false|C0005847|interventionnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Podiatry (discipline)|Title|false|false||podiatrynull|Total|Modifier|false|false||totalnull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C0332840;C0002688;C1546539|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|Lacking|Modifier|false|false||lacknull|Clinical NEC (not elsewhere classified in LNC)|Finding|false|false||clinicalnull|Clinical|Modifier|false|false||clinicalnull|Improvement|Finding|false|false||improvementnull|Blood Cell Count|Procedure|false|false|C0007634;C0005773|blood cell count
null|Complete Blood Count|Procedure|false|false|C0007634;C0005773|blood cell countnull|Blood Cells|Anatomy|false|false|C0851353;C0005771;C0009555|blood cellnull|Blood and lymphatic system disorders|Disorder|false|false|C0007634;C0005773|bloodnull|peripheral blood|Finding|false|false|C0007634|blood
null|Blood|Finding|false|false|C0007634|blood
null|In Blood|Finding|false|false|C0007634|bloodnull|Cell Count|Procedure|false|false|C0007634|cell countnull|CELP gene|Finding|false|false|C0007634|cell
null|CEL gene|Finding|false|false|C0007634|cellnull|Cells|Anatomy|false|false|C1413336;C1413337;C0007584;C0005768;C0229664;C0005767;C0851353;C0005771;C0009555|cellnull|Cell Device|Device|false|false||cell
null|Cellular Phone|Device|false|false||cellnull|Cell (compartment)|Modifier|false|false||cellnull|Count Dosing Unit|LabModifier|false|false||count
null|Count|LabModifier|false|false||countnull|Pathology report|Finding|false|false||pathology reportnull|Pathology processes|Finding|false|false||pathology
null|Pathological aspects|Finding|false|false||pathologynull|Pathology procedure|Procedure|false|false||pathologynull|Pathology|Title|false|false||pathologynull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Cleaning (activity)|Event|false|false||cleannull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Have Pain|Finding|false|false||have painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Erythema|Disorder|false|false|C1515974|erythemanull|Swelling|Finding|false|false|C1515974|swelling
null|Edema|Finding|false|false|C1515974|swellingnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgical
null|Surgical service|Procedure|false|false|C1515974|surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C0013604;C0038999;C1546778;C0041834;C0543467;C0587668|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|CYREN gene|Finding|false|false||MRInull|Magnetic resonance imaging service|Procedure|false|false||MRI
null|Magnetic Resonance Imaging|Procedure|false|false||MRInull|Maori Language|Entity|false|false||MRInull|Structure of left foot|Anatomy|false|false|C0555980;C1552822|left footnull|Table Cell Horizontal Align - left|Finding|false|false|C0230461;C4299097;C0016504|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C1552822|foot
null|Foot|Anatomy|false|false|C0555980;C1552822|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Surgical Flaps|Anatomy|false|false|C1717255;C0543467;C0587668;C1705203;C1427618;C0013604;C1412362|surgical flapnull|Operative Surgical Procedures|Procedure|false|false|C0038925;C0038925|surgical
null|Surgical service|Procedure|false|false|C0038925;C0038925|surgicalnull|ALOX5AP gene|Finding|false|false|C0038925;C0038925|flapnull|Surgical Flaps|Anatomy|false|false|C1705203;C1427618;C0013604;C0543467;C0587668;C1412362|flapnull|Edema|Finding|false|false|C0038925;C0038925|edemanull|null|Attribute|false|false|C0038925|edemanull|Focal|Modifier|false|false||focalnull|Spot (mark)|Finding|false|false|C0038925;C0038925|spot
null|THEMIS gene|Finding|false|false|C0038925;C0038925|spotnull|Leiostomus xanthurus|Entity|false|false||spotnull|View spot|Modifier|false|false||spotnull|Site of|Modifier|false|false||site ofnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778;C0038895;C1457907;C1547138;C0543467|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Level of Care - Surgery|Finding|false|false|C1515974|surgery
null|Surgical procedure finding|Finding|false|false|C1515974|surgery
null|Surgical aspects|Finding|false|false|C1515974|surgerynull|Operative Surgical Procedures|Procedure|false|false|C1515974|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Aspects of signs|Finding|true|false||signs
null|Physical findings|Finding|true|false||signsnull|Manufactured sign|Device|true|false||signsnull|Abscess|Disorder|true|false||abscessnull|null|Finding|true|false||abscessnull|fluid - substance|Drug|true|false||fluid
null|Liquid substance|Drug|true|false||fluidnull|Fluid Specimen Code|Finding|true|false||fluidnull|Fluid behavior|Modifier|false|false||fluidnull|Collection Object - UML Entity|Finding|false|false||collection
null|Item Collection|Finding|false|false||collection
null|Collections (publication)|Finding|false|false||collection
null|Collection (action)|Finding|false|false||collectionnull|Podiatry (discipline)|Title|false|false||Podiatrynull|Team|Subject|false|false||teamnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Surgical intervention (finding)|Finding|false|false||surgical interventionnull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|Intervention regimes|Procedure|false|false||intervention
null|Nursing interventions|Procedure|false|false||intervention
null|Interventional procedure|Procedure|false|false||interventionnull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false|C0230346;C4048756|line
null|Long Interspersed Elements|Drug|false|false|C0230346;C4048756|line
null|Long Interspersed Elements|Drug|false|false|C0230346;C4048756|linenull|line source specimen code|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Right upper arm structure|Anatomy|false|false|C1824218;C3715044;C1546701;C2049629;C1550648;C1517938;C1552823;C1522541;C5400986;C4761640;C3495676|right arm
null|Right arm|Anatomy|false|false|C1824218;C3715044;C1546701;C2049629;C1550648;C1517938;C1552823;C1522541;C5400986;C4761640;C3495676|right armnull|Table Cell Horizontal Align - right|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078;C0230346;C4048756|armnull|AKR1A1 wt Allele|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1824218;C3715044;C3495676;C1546701;C1522541;C5400986;C4761640;C1552823;C2049629|arm
null|null|Anatomy|false|false|C1824218;C3715044;C3495676;C1546701;C1522541;C5400986;C4761640;C1552823;C2049629|arm
null|Upper Extremity|Anatomy|false|false|C1824218;C3715044;C3495676;C1546701;C1522541;C5400986;C4761640;C1552823;C2049629|armnull|Infantile Neuroaxonal Dystrophy|Disorder|false|false||plannull|Treatment Plan|Finding|false|false||plan
null|Planned|Finding|false|false||plan
null|null|Finding|false|false||plannull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Course|Time|false|false||coursenull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Podiatry (discipline)|Title|false|false||podiatrynull|Daily|Time|false|false||dailynull|Dressing Dosage Form|Drug|false|false|C0230461|dressingnull|Ability to dress|Finding|false|false|C0230461;C4299097;C0016504|dressing
null|null|Finding|false|false|C0230461;C4299097;C0016504|dressingnull|Dressing patient (procedure)|Procedure|false|false|C0230461;C4299097;C0016504|dressing
null|Dressing of skin or wound|Procedure|false|false|C0230461;C4299097;C0016504|dressingnull|Medical dressing|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Wound Dressings (device)|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Changing|Finding|false|false|C0230461;C4299097;C0016504|changesnull|Changed status|LabModifier|false|false||changesnull|Structure of left foot|Anatomy|false|false|C1552822;C1305428;C0518459;C0392747;C0555980;C0152053;C0278286;C1705365|left footnull|Table Cell Horizontal Align - left|Finding|false|false|C0230461|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C1305428;C0518459;C0555980;C0392747;C0152053;C0278286|foot
null|Foot|Anatomy|false|false|C1305428;C0518459;C0555980;C0392747;C0152053;C0278286|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Betadine|Drug|false|false||Betadine
null|Betadine|Drug|false|false||Betadinenull|Gauzes|Device|false|false||gauzenull|Gauzes|Device|false|false||gauzenull|Cough (guaifenesin)|Drug|false|false||Cough
null|Cough (guaifenesin)|Drug|false|false||Coughnull|Coughing|Finding|false|false||Coughnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Atelectasis|Finding|false|false||atelectasisnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Remote control command - Clear|Finding|false|false||clearnull|Clear|Modifier|false|false||clear
null|Transparent (qualitative concept)|Modifier|false|false||clearnull|Coughing|Finding|false|false||coughingnull|Repeat Object|Finding|false|false||repeat
null|Repeat|Finding|false|false||repeatnull|Repeat Pattern|Time|false|false||repeatnull|Plain chest X-ray|Procedure|false|false|C1527391;C0817096|chest x-raynull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025;C0039985|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025;C0039985|chestnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||x-ray
null|roentgenographic|Finding|false|false||x-raynull|Plain x-ray|Procedure|false|false||x-ray
null|Diagnostic radiologic examination|Procedure|false|false||x-ray
null|Radiographic imaging procedure|Procedure|false|false||x-raynull|Roentgen Rays|Phenomenon|false|false||x-raynull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Cardiovascular disease+Pulmonary disease|Disorder|false|false|C0553534|cardiopulmonarynull|Cardiopulmonary|Anatomy|false|false|C4072686|cardiopulmonarynull|Comparison|Event|false|false||comparisonnull|Act Relationship Subset - previous|Time|false|false||previous
null|Previous|Time|false|false||previousnull|Chest problem|Finding|false|false|C1527391;C0817096|chestnull|Chest|Anatomy|false|false|C0741025|chest
null|Anterior thoracic region|Anatomy|false|false|C0741025|chestnull|ActClaimAttachmentCategoryCode - x-ray|Finding|false|false||x-ray
null|roentgenographic|Finding|false|false||x-raynull|Plain x-ray|Procedure|false|false||x-ray
null|Diagnostic radiologic examination|Procedure|false|false||x-ray
null|Radiographic imaging procedure|Procedure|false|false||x-raynull|Roentgen Rays|Phenomenon|false|false||x-raynull|Hospital Stay|Time|false|false||hospital staynull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Changing|Finding|true|false||changesnull|Changed status|LabModifier|false|false||changesnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|At discharge|Time|false|false||at dischargenull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Antihypertensive Agents|Drug|false|false||antihypertensivesnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|Systole|Finding|false|false||systolicnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|In Blood|Finding|false|false||blood
null|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Probable diagnosis|Finding|false|false||likely
null|Probably|Finding|false|false||likelynull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|contextual factors|Finding|false|false|C4299097;C0016504|settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|Diabetic foot ulcer|Disorder|false|false|C4299097;C0016504|diabetic foot ulcernull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false||diabeticnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C1456868;C0542559;C0085119;C0041582;C1547940;C1550672;C0555980;C0206172|foot
null|Foot|Anatomy|false|false|C1456868;C0542559;C0085119;C0041582;C1547940;C1550672;C0555980;C0206172|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C4299097;C0016504|ulcer
null|null|Finding|false|false|C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C4299097;C0016504|ulcernull|Firstly|Modifier|false|false||firstnull|First (number)|LabModifier|false|false||firstnull|Sterile maggot wound debridement|Procedure|false|false||debridement
null|Debridement|Procedure|false|false||debridementnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Systemic arterial pressure|Finding|false|false||blood pressuresnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressuresnull|null|Phenomenon|false|false||pressuresnull|Increase|Finding|false|false||increasenull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Systole|Finding|false|false||systolicnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|metoprolol|Drug|false|false||metoprolol
null|metoprolol|Drug|false|false||metoprololnull|Observation parameter|Finding|false|false||parametersnull|Systole|Finding|false|false||systolicnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Less Than|LabModifier|false|false||less thannull|Smaller|Modifier|false|false||lessnull|Less Than|LabModifier|false|false||lessnull|Hypertensive (finding)|Finding|false|false||hypertensivenull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Acute kidney injury|Disorder|false|false|C0227665;C0022646|Acute Kidney Injury
null|Kidney Failure, Acute|Disorder|false|false|C0227665;C0022646|Acute Kidney Injurynull|Admission Level of Care Code - Acute|Finding|false|false||Acute
null|Acute - Triage Code|Finding|false|false||Acutenull|acute|Time|false|false||Acutenull|Injury of kidney|Disorder|false|false|C0227665;C0022646|Kidney Injurynull|Neoplasm of uncertain or unknown behavior of kidney|Disorder|false|false|C0227665;C0022646|Kidney
null|Benign neoplasm of kidney|Disorder|false|false|C0227665;C0022646|Kidneynull|Kidney problem|Finding|false|false|C0227665;C0022646|Kidneynull|examination of kidney|Procedure|false|false|C0227665;C0022646|Kidney
null|Procedures on Kidney|Procedure|false|false|C0227665;C0022646|Kidneynull|Kidney|Anatomy|false|false|C4554465;C0869841;C0160420;C3263723;C3263722;C0812426;C0022660;C2609414;C0496927;C0496892|Kidney
null|Both kidneys|Anatomy|false|false|C4554465;C0869841;C0160420;C3263723;C3263722;C0812426;C0022660;C2609414;C0496927;C0496892|Kidneynull|Traumatic AND/OR non-traumatic injury|Disorder|false|false|C0227665;C0022646|Injury
null|Traumatic injury|Disorder|false|false|C0227665;C0022646|Injurynull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|contextual factors|Finding|false|false||settingnull|Settings (qualitative concept)|Modifier|false|false||settingnull|Sepsis|Disorder|false|false||sepsis
null|Septicemia|Disorder|false|false||sepsisnull|Sepsis <Sepsidae>|Entity|false|false||sepsisnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Hypotension|Finding|false|false||hypotensionnull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Measures (attribute)|Finding|false|false||measuresnull|Measures|LabModifier|false|false||measuresnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|BaseLine dental cement|Drug|false|false||baselinenull|baseline - TableCellVerticalAlign|Finding|false|false||baselinenull|Baseline|LabModifier|false|false||baselinenull|Chronic - Admission Level of Care Code|Finding|false|false||CHRONICnull|Provision of recurring care for chronic illness|Procedure|false|false||CHRONICnull|chronic|Time|false|false||CHRONICnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes Mellitus Type 2null|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Type 2|Finding|false|false||Type 2null|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Patient Admission|Procedure|false|false||admission, patientnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|Relationship modifier - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Dosage|LabModifier|false|false||dosesnull|Lantus|Drug|false|false||Lantus
null|Lantus|Drug|false|false||Lantusnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Humalog|Drug|false|false||Humalog
null|Humalog|Drug|false|false||Humalognull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit of Measure|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|3 times|Finding|false|false||3 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Daily|Time|false|false||dailynull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Hardness|Modifier|false|false||hardnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Diagnosis Type - Working|Finding|false|false||Workingnull|Work|Event|false|false||Workingnull|Working animal|Entity|false|false||Workingnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||diabetes
null|Diabetes|Disorder|false|false||diabetes
null|Diabetes Mellitus|Disorder|false|false||diabetesnull|Consultation|Procedure|false|false||consultnull|Team|Subject|false|false||teamnull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|Dosage|LabModifier|false|false||dosesnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Unit of Measure|LabModifier|false|false||units
null|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|Toujeo|Drug|false|false||Toujeo
null|Toujeo|Drug|false|false||Toujeonull|Unit of Measure|LabModifier|false|false||units
null|Unit - NCI Thesaurus Property|LabModifier|false|false||units
null|Unit|LabModifier|false|false||unitsnull|With meals|Time|false|false||with mealsnull|Meal (occasion for eating)|Finding|false|false||mealsnull|With meals|Time|false|false||mealsnull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Tradjenta|Drug|false|false||Trajenta
null|Tradjenta|Drug|false|false||Trajentanull|Jardiance|Drug|false|false||Jardiance
null|Jardiance|Drug|false|false||Jardiancenull|CODE STATUS|Procedure|false|false||CODE STATUSnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|What subject filter - Status|Finding|false|false||STATUSnull|null|Attribute|false|false||STATUSnull|Social status|Modifier|false|false||STATUS
null|Status|Modifier|false|false||STATUSnull|Full|Modifier|false|false||Fullnull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|Grandson|Subject|false|false||grandsonnull|Girlfriend|Subject|false|false||girlfriendnull|Marketing basis - Transitional|Finding|false|false||TRANSITIONALnull|Transitional cell morphology|Modifier|false|false||TRANSITIONALnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Every eight hours|Time|false|false||Q8Hnull|soft tissue pain in foot|Finding|false|false|C4299097;C0016504|foot pain
null|Foot pain|Finding|false|false|C4299097;C0016504|foot painnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C0016512;C2016948|foot
null|Foot|Anatomy|false|false|C0555980;C0016512;C2016948|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|BMP1 protein, human|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Phencyclidine|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|Pentachlorophenol|Drug|false|false||PCP
null|BMP1 protein, human|Drug|false|false||PCPnull|PCP - Hallucinogen-Related Disorder|Disorder|false|false||PCP
null|Pneumocystis jiroveci pneumonia|Disorder|false|false||PCP
null|Papillary craniopharyngioma|Disorder|false|false||PCPnull|obsolete serine-type Pro-X carboxypeptidase activity|Finding|false|false||PCP
null|BMP1 wt Allele|Finding|false|false||PCP
null|PGPEP1 gene|Finding|false|false||PCP
null|peptidyl carrier protein activity|Finding|false|false||PCP
null|PRCP gene|Finding|false|false||PCPnull|Primary care provider|Subject|false|false||PCPnull|Appointments|Event|false|false||appointmentnull|Pain management (procedure)|Procedure|false|false||pain managementnull|Pain Management (specialty)|Title|false|false||pain managementnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Disease Management|Procedure|false|false||managementnull|Management Occupations|Subject|false|false||managementnull|Management procedure|Event|false|false||management
null|Administration occupational activities|Event|false|false||managementnull|Osteomyelitis|Disorder|false|false||Osteomyelitisnull|Infected|Finding|false|false||infectednull|Diabetic foot ulcer|Disorder|false|false|C4299097;C0016504|diabetic foot ulcernull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false||diabeticnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C1456868;C0206172;C0555980;C0085119;C0041582;C1547940;C1550672|foot
null|Foot|Anatomy|false|false|C1456868;C0206172;C0555980;C0085119;C0041582;C1547940;C1550672|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C4299097;C0016504|ulcer
null|null|Finding|false|false|C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C4299097;C0016504|ulcernull|Surgical margins|Anatomy|false|false|C0543467;C0587668;C4761388|Surgical marginnull|Operative Surgical Procedures|Procedure|false|false|C0229985|Surgical
null|Surgical service|Procedure|false|false|C0229985|Surgicalnull|null|Finding|false|false|C0229985|marginnull|Marginal|Modifier|false|false||marginnull|Total|Modifier|false|false||totalnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C0002688;C1546539;C1552822;C0332840|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|Negative|Finding|false|false||negative fornull|Rh Negative Blood Group|Finding|false|false||negative
null|Negative|Finding|false|false||negative
null|Negative Finding|Finding|false|false||negativenull|Expression Negative|Lab|false|false||negativenull|Negative - qualifier|Modifier|false|false||negative
null|Negative Charge|Modifier|false|false||negativenull|Negative Number|LabModifier|false|false||negativenull|Osteomyelitis|Disorder|false|false||osteomyelitisnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Course|Time|false|false||coursenull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Continuous|Finding|false|false||ongoingnull|Soft Tissue Infection|Disorder|false|false|C0225317;C4532079;C0040300|soft tissue infectionnull|Neck+Chest>Soft tissue|Anatomy|false|false|C3542022;C0009450;C3714514;C0149778;C1547928|soft tissue
null|soft tissue|Anatomy|false|false|C3542022;C0009450;C3714514;C0149778;C1547928|soft tissuenull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false|C0040300;C0225317;C4532079|softnull|Soft|Modifier|false|false||softnull|Tissue Specimen Code|Finding|false|false|C0040300;C0225317;C4532079|tissuenull|Body tissue|Anatomy|false|false|C3542022;C3714514;C1547928;C0009450;C0149778|tissuenull|Communicable Diseases|Disorder|false|false|C0225317;C4532079;C0040300|infectionnull|Infection|Finding|false|false|C0225317;C4532079;C0040300|infectionnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|completion - ResponseLevel|Modifier|false|false||completion
null|Complete|Modifier|false|false||completionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|physiologic resolution|Finding|false|false||resolution
null|Resolution|Finding|false|false||resolutionnull|Resolution Property|LabModifier|false|false||resolutionnull|Hour|Time|false|false||hournull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Once - dosing instruction fragment|Finding|false|false||Oncenull|Once (schedule frequency)|Time|false|false||Oncenull|Antibiotics|Drug|false|false||antibioticnull|Right upper arm structure|Anatomy|false|false|C1824218;C3715044;C3495676;C2049629;C1522541;C5400986;C4761640;C1552823;C1546701|right arm
null|Right arm|Anatomy|false|false|C1824218;C3715044;C3495676;C2049629;C1522541;C5400986;C4761640;C1552823;C1546701|right armnull|Table Cell Horizontal Align - right|Finding|false|false|C0230346;C4048756|rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|Anorectal Malformations|Disorder|false|false|C0446516;C1140618;C1269078;C0230346;C4048756|armnull|AKR1A1 wt Allele|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|ARMC9 gene|Finding|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|armnull|Protocol Treatment Arm|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|Axillary Reverse Mapping|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|arm
null|Study Arm|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|armnull|Upper arm|Anatomy|false|false|C1546701;C3495676;C1522541;C5400986;C4761640;C1824218;C3715044;C2049629|arm
null|null|Anatomy|false|false|C1546701;C3495676;C1522541;C5400986;C4761640;C1824218;C3715044;C2049629|arm
null|Upper Extremity|Anatomy|false|false|C1546701;C3495676;C1522541;C5400986;C4761640;C1824218;C3715044;C2049629|armnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICC linenull|Peripherally Inserted Central Catheter Line Insertion|Procedure|false|false|C0230346;C4048756;C0446516;C1140618;C1269078|PICCnull|Peripherally inserted central catheter (physical object)|Device|false|false||PICCnull|Line Specimen|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||line
null|Long Interspersed Elements|Drug|false|false||linenull|line source specimen code|Finding|false|false|C0446516;C1140618;C1269078;C0230346;C4048756|linenull|Intravascular line|Device|false|false||linenull|Linear|Modifier|false|false||linenull|Line Unit of Length|LabModifier|false|false||linenull|Traumatic Wound|Disorder|false|false||wound
null|Wounds and Injuries|Disorder|false|false||wound
null|Traumatic injury|Disorder|false|false||woundnull|Route of Administration - Wound|Finding|false|false||wound
null|null|Finding|false|false||wound
null|Specimen Type - Wound|Finding|false|false||woundnull|Podiatry (discipline)|Title|false|false||podiatrynull|Daily|Time|false|false||dailynull|Dressing Dosage Form|Drug|false|false||dressingnull|null|Finding|false|false||dressing
null|Ability to dress|Finding|false|false||dressingnull|Dressing of skin or wound|Procedure|false|false||dressing
null|Dressing patient (procedure)|Procedure|false|false||dressingnull|Wound Dressings (device)|Device|false|false||dressing
null|Dress (garment)|Device|false|false||dressing
null|Medical dressing|Device|false|false||dressingnull|Dressing (unit of presentation)|LabModifier|false|false||dressingnull|Changing|Finding|false|false|C0230461;C4299097;C0016504|changesnull|Changed status|LabModifier|false|false||changesnull|Structure of left foot|Anatomy|false|false|C0392747;C0555980;C1552822|left footnull|Table Cell Horizontal Align - left|Finding|false|false|C0230461|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Foot problem|Finding|false|false|C4299097;C0016504;C0230461|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C0392747|foot
null|Foot|Anatomy|false|false|C0555980;C0392747|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Operative site|Modifier|false|false||surgical sitenull|Operative Surgical Procedures|Procedure|false|false||surgical
null|Surgical service|Procedure|false|false||surgicalnull|null|Finding|false|false|C1515974|sitenull|Anatomic Site|Anatomy|false|false|C1546778|sitenull|Study Site|Modifier|false|false||site
null|Site|Modifier|false|false||sitenull|Betadine|Drug|false|false||Betadine
null|Betadine|Drug|false|false||Betadinenull|Gauzes|Device|false|false||gauzenull|Gauzes|Device|false|false||gauzenull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes mellitus type 2null|Diabetes Mellitus|Disorder|false|false||Diabetes mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Type 2|Finding|false|false||type 2null|Type - ParameterizedDataType|Finding|false|false||type
null|SGCG gene|Finding|false|false||typenull|null|Modifier|false|false||typenull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Blood Glucose|Drug|false|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|Very|Modifier|false|false||verynull|Diabetic foot ulcer|Disorder|false|false|C4299097;C0016504|diabetic foot ulcernull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false|C4299097;C0016504|diabeticnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0041582;C1547940;C1550672;C0206172;C0085119;C0555980;C1456868;C0241863|foot
null|Foot|Anatomy|false|false|C0041582;C1547940;C1550672;C0206172;C0085119;C0555980;C1456868;C0241863|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C4299097;C0016504|ulcer
null|null|Finding|false|false|C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C4299097;C0016504|ulcernull|Blood Glucose|Drug|true|false||blood sugarsnull|Blood and lymphatic system disorders|Disorder|true|false||bloodnull|peripheral blood|Finding|true|false||blood
null|Blood|Finding|true|false||blood
null|In Blood|Finding|true|false||bloodnull|Sugars|Drug|true|false||sugars
null|Sugars|Drug|true|false||sugarsnull|sugars (lab test)|Procedure|true|false||sugarsnull|Well (answer to question)|Finding|true|false||wellnull|Well (container)|Device|true|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Diabetic|Finding|false|false||diabeticnull|Medication Regimen|Procedure|false|false||medication regimennull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Unit dose|LabModifier|false|false||dose
null|Dosage|LabModifier|false|false||dosenull|Toujeo|Drug|false|false||Toujeo
null|Toujeo|Drug|false|false||Toujeonull|Regular|Modifier|false|false||regularnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Usual|Modifier|false|false||usualnull|Tradjenta|Drug|false|false||Trajenta
null|Tradjenta|Drug|false|false||Trajentanull|Jardiance|Drug|false|false||Jardiance
null|Jardiance|Drug|false|false||Jardiancenull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Patient need for (contextual qualifier)|Finding|false|false||need fornull|Patient need for (contextual qualifier)|Finding|false|false||neednull|Needs|Modifier|false|false||neednull|Jardiance|Drug|false|false||Jardiance
null|Jardiance|Drug|false|false||Jardiancenull|Medical History|Finding|false|false||history ofnull|History of present illness (finding)|Finding|false|false||history
null|History of previous events|Finding|false|false||history
null|Historical aspects qualifier|Finding|false|false||history
null|Medical History|Finding|false|false||history
null|Concept History|Finding|false|false||historynull|History|Subject|false|false||historynull|Recurrent|Time|false|false||recurrent
null|Episodic|Time|false|false||recurrentnull|Akis|Entity|false|false||AKIsnull|Cough (guaifenesin)|Drug|false|false||Cough
null|Cough (guaifenesin)|Drug|false|false||Coughnull|Coughing|Finding|false|false||Coughnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Cough (guaifenesin)|Drug|false|false||cough
null|Cough (guaifenesin)|Drug|false|false||coughnull|Coughing|Finding|false|false||coughnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Apyrexial|Finding|false|false||afebrilenull|Leukocytosis|Disorder|true|false||leukocytosisnull|Blood leukocyte number above reference range|Finding|true|false||leukocytosisnull|Plain chest X-ray|Procedure|true|false||CXRnull|Aspects of signs|Finding|true|false|C0032225|signs
null|Physical findings|Finding|true|false|C0032225|signsnull|Manufactured sign|Device|true|false||signsnull|Pleural Diseases|Disorder|true|false|C0032225|pleuralnull|Pleura|Anatomy|false|false|C0220912;C0311392;C0032226|pleuralnull|Pleural|Modifier|false|false||pleuralnull|Effusion (substance)|Finding|false|false||effusion
null|null|Finding|false|false||effusion
null|effusion|Finding|false|false||effusionnull|Lung consolidation|Disorder|false|false||consolidationnull|Consolidation|Modifier|false|false||consolidationnull|Atelectasis|Finding|false|false||atelectasisnull|Menstruation|Finding|false|false||periodnull|Clinical Trial Period|Procedure|false|false||periodnull|per period (qualifier value)|Time|false|false||period
null|Time periods|Time|false|false||periodnull|Transaction counts and value totals - Period|LabModifier|false|false||periodnull|Operative procedure on foot|Procedure|false|false|C4299097;C0016504|foot surgerynull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0188413;C0555980;C0038895;C1457907;C1547138;C0543467|foot
null|Foot|Anatomy|false|false|C0188413;C0555980;C0038895;C1457907;C1547138;C0543467|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Level of Care - Surgery|Finding|false|false|C4299097;C0016504|surgery
null|Surgical procedure finding|Finding|false|false|C4299097;C0016504|surgery
null|Surgical aspects|Finding|false|false|C4299097;C0016504|surgerynull|Operative Surgical Procedures|Procedure|false|false|C4299097;C0016504|surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Incentives|Modifier|false|false||incentivenull|Spirometer Device|Device|false|false||spirometernull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Lasix|Drug|false|false||Lasix
null|Lasix|Drug|false|false||Lasixnull|Further|Modifier|false|false||furthernull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Regular|Modifier|false|false||regularnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Referral category - Inpatient|Finding|false|false||inpatient
null|Patient Class - Inpatient|Finding|false|false||inpatientnull|inpatient encounter|Procedure|false|false||inpatientnull|inpatient|Subject|false|false||inpatientnull|Hypotensive|Finding|false|false||hypotensivenull|Antihypertensive Agents|Drug|false|false||antihypertensivesnull|Blood pressure finding|Finding|false|false||blood pressure
null|Systemic arterial pressure|Finding|false|false||blood pressure
null|Blood Pressure|Finding|false|false||blood pressurenull|Blood pressure determination|Procedure|false|false||blood pressurenull|Blood and lymphatic system disorders|Disorder|false|false||bloodnull|peripheral blood|Finding|false|false||blood
null|Blood|Finding|false|false||blood
null|In Blood|Finding|false|false||bloodnull|Pressure (finding)|Finding|false|false||pressure
null|null|Finding|false|false||pressure
null|Baresthesia|Finding|false|false||pressurenull|null|Phenomenon|false|false||pressurenull|Pressure (property)|LabModifier|false|false||pressurenull|Table Cell Horizontal Align - right|Finding|false|false||rightnull|Right sided|Modifier|false|false||right
null|Right|Modifier|false|false||rightnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Too low|Finding|false|false||too lownull|IPSS-R Risk Category Low|Finding|false|false||low
null|IPSS Risk Category Low|Finding|false|false||low
null|low confidentiality|Finding|false|false||lownull|Low - MessageWaitingPriority|Modifier|false|false||low
null|low|Modifier|false|false||low
null|low exposure|Modifier|false|false||lownull|null|LabModifier|false|false||lownull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Intensity and Distress 1|Finding|false|false||slightnull|Slight (qualifier value)|Modifier|false|false||slight
null|Mild (qualifier value)|Modifier|false|false||slightnull|creatinine|Drug|false|false||creatinine
null|creatinine|Drug|false|false||creatininenull|Creatinine metabolic function|Finding|false|false||creatininenull|Creatinine measurement|Procedure|false|false||creatininenull|losartan|Drug|false|false||losartan
null|losartan|Drug|false|false||losartannull|Relationship modifier - Patient|Finding|false|false||Patient
null|Specimen Type - Patient|Finding|false|false||Patient
null|Mail Claim Party - Patient|Finding|false|false||Patient
null|Report source - Patient|Finding|false|false||Patient
null|null|Finding|false|false||Patient
null|Disabled Person Code - Patient|Finding|false|false||Patientnull|Patients|Subject|false|false||Patientnull|Veterinary Patient|Entity|false|false||Patientnull|Weekly|Time|false|false||weeklynull|Laboratory test finding|Lab|false|false||labsnull|Antibiotics|Drug|false|false||antibioticnull|Infusion procedures|Procedure|false|false||infusionsnull|risedronate|Drug|false|false||rise
null|risedronate|Drug|false|false||risenull|Relational and Item-Specific Encoding Task|Finding|false|false||risenull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|Antibiotics|Drug|false|false||antibioticnull|cefazolin|Drug|false|false||cefazolin
null|cefazolin|Drug|false|false||cefazolinnull|CODE STATUS|Procedure|false|false||CODE STATUSnull|MDF Attribute Type - Code|Finding|false|false||CODE
null|A Codes|Finding|false|false||CODE
null|Code|Finding|false|false||CODEnull|Coding|Event|false|false||CODEnull|What subject filter - Status|Finding|false|false||STATUSnull|null|Attribute|false|false||STATUSnull|Social status|Modifier|false|false||STATUS
null|Status|Modifier|false|false||STATUSnull|Full|Modifier|false|false||Fullnull|Contact - HL7 Attribution|Finding|false|false||CONTACT
null|Contact with|Finding|false|false||CONTACT
null|Communication Contact|Finding|false|false||CONTACTnull|contact person|Subject|false|false||CONTACTnull|Physical contact|Phenomenon|false|false||CONTACTnull|Personal Contact|Event|false|false||CONTACTnull|Grandson|Subject|false|false||grandsonnull|Girlfriend|Subject|false|false||girlfriendnull|per 30 minutes|Time|false|false||30 minutes
null|30 Minutes|Time|false|false||30 minutesnull|Minute of time|Time|false|false||minutesnull|Minute Unit of Plane Angle|LabModifier|false|false||minutes
null|Minute (diminutive)|LabModifier|false|false||minutes
null|Small|LabModifier|false|false||minutesnull|complex (molecular entity)|Drug|false|false||complexnull|Complex|Modifier|false|false||complexnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|MEDICATION LIST|Finding|false|false||Medication listnull|Pharmaceutical Preparations|Drug|false|false||Medicationnull|medication - HL7 publishing domain|Finding|false|false||Medication
null|Medications|Finding|false|false||Medicationnull|List|Finding|false|false||list
null|Sequence Data Type|Finding|false|false||listnull|Accurate (qualifier value)|Modifier|false|false||accuratenull|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||complete
null|Complete, Multiple Vitamins with Iron|Drug|false|false||completenull|Completion Status for valid values - Complete|Finding|false|false||complete
null|Data operation - complete|Finding|false|false||complete
null|Finish - dosing instruction imperative|Finding|false|false||completenull|Complete|Modifier|false|false||completenull|canagliflozin|Drug|false|false||canagliflozin
null|canagliflozin|Drug|false|false||canagliflozinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|ropinirole|Drug|false|false||rOPINIRole
null|ropinirole|Drug|false|false||rOPINIRolenull|Once a day, at bedtime|Time|false|false||QHSnull|Restless Legs Syndrome|Disorder|false|false|C1140621;C0023216|restless leg syndromenull|Restless Legs Syndrome|Disorder|false|false|C1140621;C0023216|restless legnull|Restlessness|Finding|false|false||restless
null|Agitation|Finding|false|false||restlessnull|Leg|Anatomy|false|false|C0035258;C0035258;C0039082|leg
null|Lower Extremity|Anatomy|false|false|C0035258;C0035258;C0039082|legnull|Syndrome|Disorder|false|false|C1140621;C0023216|syndromenull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Neuropathic pain|Finding|false|false||Neuropathic pain
null|Neuralgia|Finding|false|false||Neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|linagliptin|Drug|false|false||linaGLIPtin
null|linagliptin|Drug|false|false||linaGLIPtinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false||PTCH
null|PTCH1 wt Allele|Finding|false|false||PTCH
null|PTCH1 gene|Finding|false|false||PTCH
null|PTCH1 protein, human|Finding|false|false||PTCHnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Aspirin EC|Drug|false|false||Aspirin EC
null|Aspirin EC|Drug|false|false||Aspirin ECnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|null|Drug|false|false||MetronidAZOLE Topicalnull|metronidazole|Drug|false|false||MetronidAZOLE
null|metronidazole|Drug|false|false||MetronidAZOLEnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Gel - ContainerSeparator|Drug|false|false||Gel
null|Electrophoresis Gel|Drug|false|false||Gel
null|Gel|Drug|false|false||Gel
null|Gel physical state|Drug|false|false||Gelnull|Blood group antibody screen.GEL|Procedure|false|false||Gelnull|APPL1 gene|Finding|false|false||Applnull|Daily|Time|false|false||DAILYnull|Rosacea|Disorder|false|false||Rosaceanull|Rosacea <Prayinae>|Entity|false|false||Rosaceanull|nystatin|Drug|false|false||nystatin
null|nystatin|Drug|false|false||nystatinnull|Unit/gram|LabModifier|false|false||unit/gramnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|gram|LabModifier|false|false||gramnull|Topical Dosage Form|Drug|false|false||topicalnull|Topical Route of Administration|Finding|false|false||topicalnull|Topical surface|Modifier|false|false||topicalnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Every eight hours|Time|false|false||Q8Hnull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1720374;C1527415|mouth
null|Oral region|Anatomy|false|false|C1720374;C1527415|mouthnull|Every eight hours|Time|false|false||Every 8 hoursnull|Every - dosing instruction fragment|Finding|false|false|C0230028;C0226896|Everynull|Every (qualifier)|Modifier|false|false||Everynull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|soft tissue pain in foot|Finding|false|false|C4299097;C0016504|foot pain
null|Foot pain|Finding|false|false|C4299097;C0016504|foot painnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0016512;C2016948;C0555980;C1549543;C0030193|foot
null|Foot|Anatomy|false|false|C0016512;C2016948;C0555980;C1549543;C0030193|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Administration Method - Pain|Finding|false|false|C4299097;C0016504|pain
null|Pain|Finding|false|false|C4299097;C0016504|painnull|null|Attribute|false|false||painnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Precision - second|Finding|false|false||Second
null|metastatic qualifier|Finding|false|false||Second
null|Second Suffix|Finding|false|false||Secondnull|seconds|Time|false|false||Secondnull|Second Unit of Plane Angle|LabModifier|false|false||Second
null|second (number)|LabModifier|false|false||Secondnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|bisacodyl|Drug|false|false||bisacodyl
null|bisacodyl|Drug|false|false||bisacodylnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1561538;C1561539|mouth
null|Oral region|Anatomy|false|false|C1527415;C1561538;C1561539|mouthnull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|Twice a day|Time|false|false||Twice a daynull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|nafcillin|Drug|false|false||Nafcillin
null|nafcillin|Drug|false|false||Nafcillinnull|Every four hours|Time|false|false||Q4Hnull|nafcillin|Drug|false|false||nafcillin
null|nafcillin|Drug|false|false||nafcillinnull|glucose|Drug|false|false||dextrose
null|glucose|Drug|false|false||dextrose
null|glucose|Drug|false|false||dextrosenull|intravenous infusion of intravenous dextrose|Procedure|false|false||dextrosenull|OSM protein, human|Drug|false|false||osm
null|ovine sialomucin|Drug|false|false||osm
null|ovine sialomucin|Drug|false|false||osm
null|OSM protein, human|Drug|false|false||osm
null|Recombinant Oncostatin M|Drug|false|false||osm
null|Recombinant Oncostatin M|Drug|false|false||osmnull|OSM gene|Finding|false|false||osm
null|CCM2 gene|Finding|false|false||osmnull|osmole (unit of measure)|LabModifier|false|false||osmnull|gram|LabModifier|false|false||gramnull|Every - dosing instruction fragment|Finding|false|false||Everynull|Every (qualifier)|Modifier|false|false||Everynull|Hour|Time|false|false||hoursnull|Intravenous Route of Administration|Finding|false|false||Intravenousnull|Intravenous|Modifier|false|false||Intravenousnull|Bag Data Type|Finding|false|false||Bagnull|null|Device|false|false||Bagnull|Bag (unit of presentation)|LabModifier|false|false||Bag
null|Bag Dosing Unit|LabModifier|false|false||Bagnull|refill|Finding|false|false||Refillsnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Moderate - Severity of Illness Code|Finding|false|false||Moderate
null|Moderate|Finding|false|false||Moderatenull|Moderate (severity modifier)|Modifier|false|false||Moderate
null|Moderate - Allergy Severity|Modifier|false|false||Moderate
null|Moderation|Modifier|false|false||Moderatenull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|capsulenull|Capsule Shape|Modifier|false|false||capsulenull|Capsule (unit of presentation)|LabModifier|false|false||capsule
null|Capsule Dosing Unit|LabModifier|false|false||capsulenull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415|mouth
null|Oral region|Anatomy|false|false|C1527415|mouthnull|8 Hours|Time|false|false||8 hoursnull|Hour|Time|false|false||hoursnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|soft tissue pain in foot|Finding|false|false|C4299097;C0016504|foot pain
null|Foot pain|Finding|false|false|C4299097;C0016504|foot painnull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0555980;C0016512;C2016948;C1549543;C0030193|foot
null|Foot|Anatomy|false|false|C0555980;C0016512;C2016948;C1549543;C0030193|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Administration Method - Pain|Finding|false|false|C4299097;C0016504|pain
null|Pain|Finding|false|false|C4299097;C0016504|painnull|null|Attribute|false|false||painnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|sennosides, USP|Drug|false|false||Senna
null|sennosides, USP|Drug|false|false||Sennanull|Senna alexandrina|Entity|false|false||Senna
null|Senna Plant|Entity|false|false||Sennanull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|Firstly|Modifier|false|false||Firstnull|First (number)|LabModifier|false|false||Firstnull|Line Specimen|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Line
null|Long Interspersed Elements|Drug|false|false||Linenull|line source specimen code|Finding|false|false||Linenull|Intravascular line|Device|false|false||Linenull|Linear|Modifier|false|false||Linenull|Line Unit of Length|LabModifier|false|false||Linenull|sennosides, USP|Drug|false|false||sennosides
null|sennosides, USP|Drug|false|false||sennosidesnull|sennosides, USP|Drug|false|false||senna
null|sennosides, USP|Drug|false|false||sennanull|Senna alexandrina|Entity|false|false||senna
null|Senna Plant|Entity|false|false||sennanull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Twice a day|Time|false|false||Twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Constipation|Finding|false|false||constipationnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Breakfast|Finding|false|false||Breakfastnull|With breakfast|Time|false|false||Breakfastnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Lunch|Finding|false|false||Lunchnull|With lunch|Time|false|false||Lunchnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Units
null|Unit of Measure|LabModifier|false|false||Units
null|Unit|LabModifier|false|false||Unitsnull|Dinner|Finding|false|false||Dinnernull|With dinner|Time|false|false||Dinnernull|albuterol sulfate|Drug|false|false||albuterol sulfate
null|albuterol sulfate|Drug|false|false||albuterol sulfatenull|albuterol|Drug|false|false||albuterol
null|albuterol|Drug|false|false||albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|mcg/actuation|LabModifier|false|false||mcg/actuationnull|microgram|LabModifier|false|false||mcgnull|Actuation (unit of presentation)|LabModifier|false|false||actuationnull|Inhalation Route of Administration|Finding|false|false||inhalation
null|Inspiration (function)|Finding|false|false||inhalationnull|Inhalation Dosing Unit|LabModifier|false|false||inhalationnull|Every four hours|Time|false|false||Q4Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Aspirin EC|Drug|false|false||Aspirin EC
null|Aspirin EC|Drug|false|false||Aspirin ECnull|aspirin|Drug|false|false||Aspirin
null|aspirin|Drug|false|false||Aspirinnull|Daily|Time|false|false||DAILYnull|atorvastatin|Drug|false|false||Atorvastatin
null|atorvastatin|Drug|false|false||Atorvastatinnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|canagliflozin|Drug|false|false||canagliflozin
null|canagliflozin|Drug|false|false||canagliflozinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|fluticasone propionate|Drug|false|false||Fluticasone Propionate
null|fluticasone propionate|Drug|false|false||Fluticasone Propionatenull|fluticasone|Drug|false|false||Fluticasone
null|fluticasone|Drug|false|false||Fluticasonenull|propionate|Drug|false|false||Propionate
null|Propionates|Drug|false|false||Propionatenull|Puff Dosing Unit|LabModifier|false|false||PUFF
null|Picofarad|LabModifier|false|false||PUFFnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|furosemide|Drug|false|false||Furosemide
null|furosemide|Drug|false|false||Furosemidenull|Daily|Time|false|false||DAILYnull|gabapentin|Drug|false|false||Gabapentin
null|gabapentin|Drug|false|false||Gabapentinnull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Neuropathic pain|Finding|false|false||Neuropathic pain
null|Neuralgia|Finding|false|false||Neuropathic painnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|PTCH1 protein, human|Drug|false|false||PTCHnull|PTCH gene|Finding|false|false||PTCH
null|PTCH1 wt Allele|Finding|false|false||PTCH
null|PTCH1 gene|Finding|false|false||PTCH
null|PTCH1 protein, human|Finding|false|false||PTCHnull|QPM|Time|false|false||QPM
null|Once a day, in the evening|Time|false|false||QPMnull|linagliptin|Drug|false|false||linaGLIPtin
null|linagliptin|Drug|false|false||linaGLIPtinnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Daily|Time|false|false||DAILYnull|losartan potassium|Drug|false|false||Losartan Potassium
null|losartan potassium|Drug|false|false||Losartan Potassiumnull|losartan|Drug|false|false||Losartan
null|losartan|Drug|false|false||Losartannull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|Daily|Time|false|false||DAILYnull|metoprolol succinate|Drug|false|false||Metoprolol Succinate
null|metoprolol succinate|Drug|false|false||Metoprolol Succinatenull|metoprolol|Drug|false|false||Metoprolol
null|metoprolol|Drug|false|false||Metoprololnull|succinate|Drug|false|false||Succinate
null|Succinates|Drug|false|false||Succinatenull|Daily|Time|false|false||DAILYnull|null|Drug|false|false||MetronidAZOLE Topicalnull|metronidazole|Drug|false|false||MetronidAZOLE
null|metronidazole|Drug|false|false||MetronidAZOLEnull|Topical Dosage Form|Drug|false|false||Topicalnull|Topical Route of Administration|Finding|false|false||Topicalnull|Topical surface|Modifier|false|false||Topicalnull|Gel - ContainerSeparator|Drug|false|false||Gel
null|Electrophoresis Gel|Drug|false|false||Gel
null|Gel|Drug|false|false||Gel
null|Gel physical state|Drug|false|false||Gelnull|Blood group antibody screen.GEL|Procedure|false|false||Gelnull|APPL1 gene|Finding|false|false||Applnull|Daily|Time|false|false||DAILYnull|Rosacea|Disorder|false|false||Rosaceanull|Rosacea <Prayinae>|Entity|false|false||Rosaceanull|nitroglycerin|Drug|false|false||Nitroglycerin
null|nitroglycerin|Drug|false|false||Nitroglycerinnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Angina Pectoris|Finding|false|false||angina
null|null|Finding|false|false||anginanull|null|Attribute|false|false||anginanull|nystatin|Drug|false|false||nystatin
null|nystatin|Drug|false|false||nystatinnull|Unit/gram|LabModifier|false|false||unit/gramnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|gram|LabModifier|false|false||gramnull|Topical Dosage Form|Drug|false|false||topicalnull|Topical Route of Administration|Finding|false|false||topicalnull|Topical surface|Modifier|false|false||topicalnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|oxycodone|Drug|false|false||OxyCODONE
null|oxycodone|Drug|false|false||OxyCODONEnull|Oxycodone measurement|Procedure|false|false||OxyCODONEnull|Acetaminophen [EPC]|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophen
null|acetaminophen|Drug|false|false||Acetaminophennull|Acetaminophen measurement|Procedure|false|false||Acetaminophennull|Tablet Dosage Form|Drug|false|false||TABnull|Tablet Dosing Unit|LabModifier|false|false||TABnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||Pain
null|Pain|Finding|false|false||Painnull|null|Attribute|false|false||Painnull|Severe - Severity of Illness Code|Finding|false|false||Severe
null|Intensity and Distress 5|Finding|false|false||Severe
null|Severe - Triage Code|Finding|false|false||Severe
null|Severe (severity modifier)|Finding|false|false||Severe
null|Allergy Severity - Severe|Finding|false|false||Severenull|pantoprazole|Drug|false|false||Pantoprazole
null|pantoprazole|Drug|false|false||Pantoprazolenull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ropinirole|Drug|false|false||rOPINIRole
null|ropinirole|Drug|false|false||rOPINIRolenull|Once a day, at bedtime|Time|false|false||QHSnull|Restless Legs Syndrome|Disorder|false|false|C1140621;C0023216|restless leg syndromenull|Restless Legs Syndrome|Disorder|false|false|C1140621;C0023216|restless legnull|Restlessness|Finding|false|false||restless
null|Agitation|Finding|false|false||restlessnull|Leg|Anatomy|false|false|C0039082;C0035258;C0035258|leg
null|Lower Extremity|Anatomy|false|false|C0039082;C0035258;C0035258|legnull|Syndrome|Disorder|false|false|C1140621;C0023216|syndromenull|insulin, regular, human|Drug|false|false||Insulin
null|Insulin [EPC]|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|INS protein, human|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Therapeutic Insulin|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|Insulin Drug Class|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulin
null|insulin, regular, human|Drug|false|false||Insulinnull|INS gene|Finding|false|false||Insulinnull|Insulin measurement|Procedure|false|false||Insulinnull|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glargine
null|insulin glargine|Drug|false|false||insulin glarginenull|insulin, regular, human|Drug|false|false||insulin
null|Insulin [EPC]|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|INS protein, human|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Therapeutic Insulin|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|Insulin Drug Class|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulin
null|insulin, regular, human|Drug|false|false||insulinnull|INS gene|Finding|false|false||insulinnull|Insulin measurement|Procedure|false|false||insulinnull|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glargine
null|insulin glargine|Drug|false|false||glarginenull|Unit per Milliliter|LabModifier|false|false||unit/mLnull|Storage Unit|Device|false|false||unit
null|Unit device|Device|false|false||unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||unit
null|Unit of Measure|LabModifier|false|false||unit
null|Unit|LabModifier|false|false||unit
null|Enzyme Unit|LabModifier|false|false||unitnull|per milliliter|LabModifier|false|false||/mLnull|Subcutaneous Route of Administration|Finding|false|false||subcutaneousnull|subcutaneous|Modifier|false|false||subcutaneousnull|Once a day, at bedtime|Time|false|false||QHSnull|Once a day, at bedtime|Time|false|false||QHSnull|trazodone|Drug|false|false||TraZODone
null|trazodone|Drug|false|false||TraZODonenull|Once a day, at bedtime|Time|false|false||QHSnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Insomnia homeopathic medication|Drug|false|false||insomnianull|Sleeplessness|Finding|false|false||insomnianull|Referral category - Outpatient|Finding|false|false||Outpatient
null|Patient Class - Outpatient|Finding|false|false||Outpatientnull|Outpatients|Subject|false|false||Outpatientnull|AML Lab Table|Finding|false|false||Lab
null|LAT2 gene|Finding|false|false||Lab
null|EWS Lab Table|Finding|false|false||Labnull|Laboratory|Device|false|false||Labnull|Labrador retriever|Entity|false|false||Lab
null|Laboratory|Entity|false|false||Labnull|Work|Event|false|false||Worknull|International Statistical Classification of Diseases and Related Health Problems, Tenth Revision (ICD-10)|Finding|false|false||ICD-10null|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|Weekly|Time|false|false||weeklynull|Laboratory Procedures|Procedure|false|false|C4318744|LAB TESTnull|AML Lab Table|Finding|false|false|C4318744|LAB
null|LAT2 gene|Finding|false|false|C4318744|LAB
null|EWS Lab Table|Finding|false|false|C4318744|LABnull|Laboratory|Device|false|false||LABnull|Labrador retriever|Entity|false|false||LAB
null|Laboratory|Entity|false|false||LABnull|Tests (qualifier value)|Finding|false|false|C4318744|TEST
null|Testing|Finding|false|false|C4318744|TESTnull|Laboratory Procedures|Procedure|false|false|C4318744|TESTnull|Test - temporal region|Anatomy|false|false|C0022885;C0456984;C0022885;C5420098;C5420670;C1825793;C0039593;C0392366|TESTnull|Test Result|Lab|false|false|C4318744|TESTnull|Test Dosing Unit|LabModifier|false|false||TESTnull|complete blood count with differential|Procedure|false|false|C2263086|CBC with differentialnull|Complete Blood Count|Procedure|false|false|C2263086|CBCnull|Nuclear cap binding complex location|Anatomy|false|false|C0545131;C0009555;C0005845;C1549478|CBCnull|Amount type - Differential|Finding|false|false|C2263086|differentialnull|Differential (qualifier value)|Modifier|false|false||differential
null|Different|Modifier|false|false||differential
null|Differential - view|Modifier|false|false||differentialnull|Blood Urea Nitrogen|Drug|false|false||BUN
null|Blood Urea Nitrogen|Drug|false|false||BUNnull|Blood urea nitrogen measurement|Procedure|false|false|C2263086|BUNnull|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|Aspartate Transaminase|Drug|false|false|C1185650|AST
null|SGOT - Glutamate oxaloacetate transaminase|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|AST
null|SLC17A5 protein, human|Drug|false|false|C1185650|ASTnull|Atypical Spitz Nevus|Disorder|false|false|C1185650|ASTnull|SLC17A5 wt Allele|Finding|false|false|C1185650|AST
null|SLC17A5 gene|Finding|false|false|C1185650|AST
null|GOT1 gene|Finding|false|false|C1185650|ASTnull|Asterion|Anatomy|false|false|C2257651;C1415274;C1140170;C4522245;C0004002;C0242192;C1121182;C1415181;C1420113;C5960784;C1266129;C1370889;C4553172|ASTnull|Asturian Language|Entity|false|false||ASTnull|Atlantic Standard Time|Time|false|false||ASTnull|Alanine Transaminase|Drug|false|false||ALT
null|Alanine Transaminase|Drug|false|false||ALTnull|Liposarcoma, well differentiated|Disorder|false|false|C1185650|ALT
null|Atypical Lipoma|Disorder|false|false|C1185650|ALTnull|null|Finding|false|false|C1185650|ALT
null|Alternative Billing Concepts|Finding|false|false|C1185650|ALT
null|GPT gene|Finding|false|false|C1185650|ALTnull|Antibiotic Lock Therapy|Procedure|false|false|C1185650|ALTnull|Southern Altai Language|Entity|false|false||ALTnull|Total|Modifier|false|false||Totalnull|Alkaline Phosphatase|Drug|false|false||ALK PHOS
null|Alkaline Phosphatase|Drug|false|false||ALK PHOSnull|Alkaline phosphatase measurement|Procedure|false|false||ALK PHOSnull|ALK protein, human|Drug|false|false||ALK
null|ALK protein, human|Drug|false|false||ALKnull|ALK protein, human|Finding|false|false||ALK
null|ALK gene|Finding|false|false||ALK
null|ALK wt Allele|Finding|false|false||ALKnull|Phos <Photinae>|Entity|false|false||PHOSnull|Extended Rotated Sidebent|Finding|false|false||ESR
null|ESR1 wt Allele|Finding|false|false||ESR
null|ESR1 gene|Finding|false|false||ESRnull|Erythrocyte sedimentation rate measurement|Procedure|false|false||ESR
null|Electron Spin Resonance Spectroscopy|Procedure|false|false||ESRnull|null|LabModifier|false|false||ESRnull|C-Reactive Protein, human|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-reactive protein|Drug|false|false||CRP
null|C-Reactive Protein, human|Drug|false|false||CRPnull|CRP wt Allele|Finding|false|false||CRP
null|CRP gene|Finding|false|false||CRP
null|CSRP1 gene|Finding|false|false||CRP
null|PPIAP10 gene|Finding|false|false||CRPnull|Pidgin and Creole language|Entity|false|false||CRPnull|Authorization Mode - Fax|Finding|false|false||FAX
null|Fax Number|Finding|false|false||FAXnull|Facsimile Machine|Device|false|false||FAX
null|Telefacsimile|Device|false|false||FAXnull|Clinic|Device|false|false||CLINIC
null|Ambulatory Care Facilities|Device|false|false||CLINICnull|Clinic|Entity|false|false||CLINIC
null|Ambulatory Care Facilities|Entity|false|false||CLINICnull|Patient location type - Clinic|Modifier|false|false||CLINIC
null|Person location type - Clinic|Modifier|false|false||CLINICnull|Authorization Mode - Fax|Finding|false|false||FAX
null|Fax Number|Finding|false|false||FAXnull|Facsimile Machine|Device|false|false||FAX
null|Telefacsimile|Device|false|false||FAXnull|Walkers|Device|false|false||Walkernull|Diagnostic, Therapeutic, and Research Equipment|Device|false|false||EQUIPMENT
null|Equipment|Device|false|false||EQUIPMENT
null|Equipment used|Device|false|false||EQUIPMENT
null|Scientific Equipment|Device|false|false||EQUIPMENTnull|Walkers|Device|false|false||Walkernull|Diagnosis Classification - Diagnosis|Finding|false|false||DIAGNOSIS
null|diagnosis aspects|Finding|false|false||DIAGNOSISnull|Diagnosis|Procedure|false|false||DIAGNOSISnull|null|Attribute|false|false||DIAGNOSISnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|Leftnull|Left sided|Modifier|false|false||Left
null|Left|Modifier|false|false||Leftnull|Hallux structure|Anatomy|false|false|C0332840;C1552822;C0002688;C1546539|halluxnull|Amputated structure (morphologic abnormality)|Disorder|false|false|C0018534|amputationnull|Amputation Specimen Code|Finding|false|false|C0018534|amputationnull|Amputation|Procedure|false|false|C0018534|amputationnull|International Statistical Classification of Diseases and Related Health Problems, Tenth Revision (ICD-10)|Finding|false|false||ICD-10null|Disruptive, Impulse Control, and Conduct Disorders|Disorder|false|false||ICD
null|Type II Mucolipidosis|Disorder|false|false||ICDnull|International Classification of Diseases|Finding|false|false||ICD
null|GNPTAB wt Allele|Finding|false|false||ICDnull|Icd Regimen|Procedure|false|false||ICDnull|between lunch and dinner|Time|false|false||ICDnull|Language Ability Proficiency - Good|Finding|false|false||Good
null|Language Proficiency - Good|Finding|false|false||Goodnull|Specimen Quality - Good|Modifier|false|false||Good
null|Good|Modifier|false|false||Goodnull|month|Time|false|false||monthsnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|ADMIN.FACILITY|Finding|false|false||Facilitynull|Facility (object)|Device|false|false||Facilitynull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Osteomyelitis|Disorder|false|false|C0018534|Osteomyelitisnull|Table Cell Horizontal Align - left|Finding|false|false|C0018534|leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Hallux structure|Anatomy|false|false|C1552822;C0029443|halluxnull|Neoplasm Metastasis|Disorder|false|false||SECONDARYnull|metastatic qualifier|Finding|false|false||SECONDARYnull|Secondary to|Modifier|false|false||SECONDARYnull|second (number)|LabModifier|false|false||SECONDARYnull|Diagnosis|Procedure|false|false||DIAGNOSESnull|Hypertensive disease|Disorder|false|false||Hypertensionnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type 2 Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Type 2 Diabetesnull|Type 2|Finding|false|false||Type 2null|Type - ParameterizedDataType|Finding|false|false||Type
null|SGCG gene|Finding|false|false||Typenull|null|Modifier|false|false||Typenull|Diabetes Mellitus|Disorder|false|false||Diabetes Mellitusnull|Diabetes Mellitus, Non-Insulin-Dependent|Disorder|false|false||Diabetes
null|Diabetes|Disorder|false|false||Diabetes
null|Diabetes Mellitus|Disorder|false|false||Diabetesnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Production Class Code - Pleasure|Finding|false|false||pleasure
null|pleasurable emotion|Finding|false|false||pleasurenull|Pleasure - Animals raised for recreation|Entity|false|false||pleasurenull|care of - AddressPartType|Finding|false|false||care ofnull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Organization unit type - Hospital|Finding|false|false||HOSPITALnull|Hospitals|Device|false|false||HOSPITALnull|Hospitals|Entity|false|false||HOSPITALnull|Hospital environment|Modifier|false|false||HOSPITALnull|Diabetic foot ulcer|Disorder|false|false|C4299097;C0016504|diabetic foot ulcernull|Diabetic Foot|Disorder|false|false|C4299097;C0016504|diabetic footnull|Diabetic|Finding|false|false|C4299097;C0016504|diabeticnull|Foot Ulcer|Disorder|false|false|C4299097;C0016504|foot ulcernull|Foot problem|Finding|false|false|C4299097;C0016504|footnull|Lower extremity>Foot|Anatomy|false|false|C0241863;C1456868;C0085119;C0206172;C0555980;C0041582;C1547940;C1550672|foot
null|Foot|Anatomy|false|false|C0241863;C1456868;C0085119;C0206172;C0555980;C0041582;C1547940;C1550672|footnull|Foot Unit of Length|LabModifier|false|false||footnull|Specimen Type - Ulcer|Finding|false|false|C4299097;C0016504|ulcer
null|null|Finding|false|false|C4299097;C0016504|ulcer
null|Ulcer|Finding|false|false|C4299097;C0016504|ulcernull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower extremity>Toes|Anatomy|false|false||toe
null|Toes|Anatomy|false|false||toenull|Very|Modifier|false|false||verynull|Infected|Finding|false|false||infectednull|Communicable Diseases|Disorder|false|false|C1442209;C0262950|infectionnull|Infection|Finding|false|false||infectionnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|bone
null|null|Finding|false|false|C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C0009450;C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C0009450;C1546560;C1550616|bonenull|Done (qualifier value)|Modifier|false|false||DONEnull|Large|LabModifier|false|false||bignull|Table Cell Horizontal Align - left|Finding|false|false||leftnull|Left sided|Modifier|false|false||left
null|Left|Modifier|false|false||leftnull|Lower extremity>Toes|Anatomy|false|false||toe
null|Toes|Anatomy|false|false||toenull|BAD protein, human|Drug|false|false||bad
null|BAD protein, human|Drug|false|false||badnull|Brachial Amyotrophic Diplegia|Disorder|false|false||badnull|BAD gene|Finding|false|false||badnull|Banda language|Entity|false|false||badnull|Bad|Modifier|false|false||badnull|Specimen Type - Bone|Finding|false|false|C1442209;C0262950|bone
null|null|Finding|false|false|C1442209;C0262950|bonenull|Skeletal bone|Anatomy|false|false|C1546560;C1550616|bone
null|XXX bone|Anatomy|false|false|C1546560;C1550616|bonenull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Communicable Diseases|Disorder|false|false||infectionnull|Infection|Finding|false|false||infectionnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|On IV|Finding|false|false||on IVnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|Leave from Employment|Finding|false|false||LEAVEnull|null|Event|false|false||LEAVEnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Injection of antibiotic|Procedure|false|false||antibiotic infusionnull|Antibiotics|Drug|false|false||antibioticnull|Infusion Pump|Device|false|false||infusion pumpnull|Location Equipment - Infusion pump|Modifier|false|false||infusion pumpnull|Infusion route|Finding|false|false||infusionnull|Infusion procedures|Procedure|false|false||infusionnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Nurses|Subject|false|false||nursenull|House (environment)|Device|false|false||housenull|Home environment|Modifier|false|false||housenull|Education (procedure)|Procedure|false|false||teachnull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||antibiotics
null|Antibiotics|Drug|false|false||antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||antibiotics
null|Antibiotics, Gynecological|Drug|false|false||antibiotics
null|antibiotics, intestinal|Drug|false|false||antibiotics
null|Antibiotic throat preparations|Drug|false|false||antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||antibiotics
null|Antibiotics for systemic use|Drug|false|false||antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||antibioticsnull|matrix metalloproteinase 7 activity|Finding|false|false||pumpnull|null|Device|false|false||pumpnull|Pump Dosing Unit|LabModifier|false|false||pumpnull|Hour|Time|false|false||hoursnull|Diabetic|Finding|false|false||diabeticnull|Medication Regimen|Procedure|false|false||medication regimennull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Close|Finding|false|false||close
null|Closed|Finding|false|false||closenull|Track (course)|Device|false|false||tracknull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Sugars|Drug|false|false||sugars
null|Sugars|Drug|false|false||sugarsnull|sugars (lab test)|Procedure|false|false||sugarsnull|4 times|Finding|false|false||4 timesnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Event Log|Finding|false|false|C0228228|lognull|lateral occipital gyrus (human only)|Anatomy|false|false|C1708728|lognull|Logarithm|LabModifier|false|false||lognull|Appointments|Event|false|false||appointmentnull|Medication Regimen|Procedure|false|false||medication regimennull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Team|Subject|false|false||teamnull|Antibiotics|Drug|false|false||antibioticnull|GDC Regimen Terminology|Finding|false|false||regimennull|Treatment Protocols|Procedure|false|false||regimennull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Care team|Finding|false|false||Care Teamnull|null|Attribute|false|false||Care Teamnull|In care (finding)|Finding|false|false||Care
null|Continuity Assessment Record and Evaluation|Finding|false|false||Carenull|care activity|Event|false|false||Carenull|Team|Subject|false|false||Teamnull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions