CUI | Concept | Semantic Group | Negated | Family History | Location | Document Text
null|MDF Attribute Type - Name|Finding|false|false||Name
null|Person Name|Finding|false|false||Name
null|Name|Finding|false|false||Namenull|Name (property) (qualifier value)|Modifier|false|false||Namenull|Storage Unit|Device|false|false||Unit
null|Unit device|Device|false|false||Unitnull|Unit - NCI Thesaurus Property|LabModifier|false|false||Unit
null|Unit of Measure|LabModifier|false|false||Unit
null|Unit|LabModifier|false|false||Unit
null|Enzyme Unit|LabModifier|false|false||Unitnull|null|Attribute|false|false||Admission Datenull|Date of admission|Time|false|false||Admission Datenull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|null|Attribute|false|false||Discharge Datenull|Discharge date|Time|false|false||Discharge Datenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient date of birth|Time|false|false||Date of Birthnull|Entity Name Part Qualifier - birth|Finding|false|false||Birth
null|Childbirth|Finding|false|false||Birth
null|birth (history)|Finding|false|false||Birth
null|Name Given at Birth|Finding|false|false||Birth
null|Birth|Finding|false|false||Birthnull|Sex Behavior|Finding|false|false||Sex
null|PLXNA3 gene|Finding|false|false||Sex
null|Coitus|Finding|false|false||Sex
null|null|Finding|false|false||Sexnull|null|Attribute|false|false||Sexnull|sex|Subject|false|false||Sex
null|Gender|Subject|false|false||Sexnull|ActInformationPrivacyReason - service|Finding|false|false||Servicenull|Software Service|Device|false|false||Servicenull|Services|Event|false|false||Servicenull|Obstetrics and gynecology (specialty)|Title|false|false||OBSTETRICS/GYNECOLOGYnull|Obstetrics service|Procedure|false|false||OBSTETRICSnull|Obstetric Patient|Subject|false|false||OBSTETRICSnull|Discipline of obstetrics|Title|false|false||OBSTETRICSnull|Gynecology|Title|false|false||GYNECOLOGYnull|Hypersensitivity|Finding|false|false||Allergiesnull|null|Attribute|false|false||Allergiesnull|codeine|Drug|false|false||Codeine
null|codeine|Drug|false|false||Codeinenull|gabapentin|Drug|false|false||gabapentin
null|gabapentin|Drug|false|false||gabapentinnull|morphine|Drug|false|false||morphine
null|morphine|Drug|false|false||morphinenull|amoxicillin|Drug|false|false||Amoxicillin
null|amoxicillin|Drug|false|false||Amoxicillinnull|metronidazole|Drug|false|false||metronidazole
null|metronidazole|Drug|false|false||metronidazolenull|propoxyphene|Drug|false|false||propoxyphene
null|propoxyphene|Drug|false|false||propoxyphenenull|Propoxyphene measurement|Procedure|false|false||propoxyphenenull|rofecoxib|Drug|false|false||rofecoxib
null|rofecoxib|Drug|false|false||rofecoxibnull|Macrobid|Drug|false|false||Macrobid
null|Macrobid|Drug|false|false||Macrobidnull|furosemide|Drug|false|false||furosemide
null|furosemide|Drug|false|false||furosemidenull|Amitiza|Drug|false|false||Amitiza
null|Amitiza|Drug|false|false||Amitizanull|sulfa|Drug|false|false||Sulfanull|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamide Anti-Infective Agents|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamides|Drug|false|false||Sulfonamide
null|Sulfonamide [EPC]|Drug|false|false||Sulfonamidenull|Antibiotics FOR TREATMENT OF HEMORRHOIDS AND ANAL FISSURES FOR TOPICAL USE|Drug|false|false||Antibiotics
null|Antibiotics|Drug|false|false||Antibiotics
null|Antibiotics, ophthalmologic|Drug|false|false||Antibiotics
null|Antibiotics, Gynecological|Drug|false|false||Antibiotics
null|antibiotics, intestinal|Drug|false|false||Antibiotics
null|Antibiotic throat preparations|Drug|false|false||Antibiotics
null|Antibiotics, Antitubercular|Drug|false|false||Antibiotics
null|Antibiotics for systemic use|Drug|false|false||Antibiotics
null|Antifungal Antibiotics, Topical|Drug|false|false||Antibioticsnull|Tylenol|Drug|false|false||Tylenol
null|Tylenol|Drug|false|false||Tylenolnull|hydromorphone|Drug|false|false||Hydromorphone
null|hydromorphone|Drug|false|false||Hydromorphonenull|Toradol|Drug|false|false||Toradol
null|Toradol|Drug|false|false||Toradolnull|Attending (action)|Finding|false|false||Attendingnull|Attending (provider role)|Subject|false|false||Attendingnull|Chief complaint (finding)|Finding|false|false||Chief Complaintnull|Complaint (finding)|Finding|false|false||Complaintnull|null|Attribute|false|false||Complaintnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Visit Priority Code - Elective|Finding|false|false||elective
null|Act Priority - elective|Finding|false|false||elective
null|Admission Type - Elective|Finding|false|false||electivenull|elective|Time|false|false||electivenull|Gynecologic Surgical Procedures|Procedure|false|false||gynecologic surgerynull|Gynecologic|Modifier|false|false||gynecologicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Urinary tract|Anatomy|false|false||urinarynull|urinary|Modifier|false|false||urinarynull|cellular entity retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Urinary Retention|Finding|false|false||retention
null|Retention of content|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Transfer - product ownership|Finding|false|false||transfer
null|Transfer Technique|Finding|false|false||transfer
null|ActClass - transfer|Finding|false|false||transfer
null|null|Finding|false|false||transfernull|Transfer (immobility management)|Procedure|false|false||transfernull|Anaphylaxis;non medication|Disorder|false|false||Anaphylaxisnull|anaphylaxis|Finding|false|false||Anaphylaxis
null|Anaphylactic shock|Finding|false|false||Anaphylaxisnull|United States Military Commissioned Officer O4 (qualifier value)|Finding|false|false||Majornull|Major <Sympycninae>|Entity|false|false||Majornull|Major|Modifier|false|false||Majornull|Operative Surgical Procedures|Procedure|false|false||Surgical
null|Surgical service|Procedure|false|false||Surgicalnull|Invasive procedure|Procedure|false|false||Invasive Procedurenull|Open approach|Modifier|false|false||Invasive Procedurenull|Invasive|Modifier|false|false||Invasivenull|Procedure (set of actions)|Finding|false|false||Procedurenull|Interventional procedure|Procedure|false|false||Procedurenull|null|Attribute|false|false||Procedurenull|Act Class - procedure|Event|false|false||Procedurenull|Stage level 2|Finding|false|false||Stage 2null|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|Posterior repair of vagina|Procedure|false|false||posterior colporrhaphy
null|Repair of rectocele|Procedure|false|false||posterior colporrhaphynull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Suture of vagina|Procedure|false|false||colporrhaphynull|Rectocele|Disorder|false|false||rectocelenull|Enterocele|Disorder|false|false||enterocelenull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|History of present illness (finding)|Finding|false|false||History of Present Illnessnull|null|Attribute|false|false||History of Present Illnessnull|Medical History|Finding|false|false||History ofnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Present illness|Finding|false|false||Present Illnessnull|Present|Finding|false|false||Present
null|Presentation|Finding|false|false||Presentnull|Illness (finding)|Finding|false|false||Illnessnull|cervical cancer|Disorder|false|false|C0027530|cervical CAnull|Neck|Anatomy|false|false|C4048328|cervicalnull|Cervical|Modifier|false|false||cervicalnull|Radical hysterectomy|Procedure|false|false||radical hysterectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Lymphedema|Disorder|false|false||lymphedemanull|Urinary Retention|Finding|false|false|C0042027|urinary retentionnull|Bladder retention of urine|Attribute|false|false||urinary retentionnull|Urinary tract|Anatomy|false|false|C0080274|urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Retention of content|Finding|false|false||retention
null|cellular entity retention|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Frequently|Time|false|false||frequentlynull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Asthma|Disorder|false|false||Asthmanull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Ichthyosis Bullosa of Siemens|Disorder|false|false||IBS
null|Irritable Bowel Syndrome|Disorder|false|false||IBSnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Fibromyalgia|Disorder|false|false||fibromyalgianull|Visit Priority Code - Elective|Finding|false|false||elective
null|Act Priority - elective|Finding|false|false||elective
null|Admission Type - Elective|Finding|false|false||electivenull|elective|Time|false|false||electivenull|Gynecologic|Modifier|false|false||gynecologicnull|Level of Care - Surgery|Finding|false|false||surgery
null|Surgical procedure finding|Finding|false|false||surgery
null|Surgical aspects|Finding|false|false||surgerynull|Operative Surgical Procedures|Procedure|false|false||surgerynull|General surgery specialty|Title|false|false||surgery
null|Surgery specialty|Title|false|false||surgerynull|Stage level 2|Finding|false|false||stage 2null|Tumor stage|Attribute|false|false||stagenull|Stage|Time|false|false||stage
null|Phase|Time|false|false||stagenull|Posterior repair of vagina|Procedure|false|false||posterior colporrhaphy
null|Repair of rectocele|Procedure|false|false||posterior colporrhaphynull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Suture of vagina|Procedure|false|false||colporrhaphynull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C0332835|graft
null|Grafting procedure|Procedure|false|false|C0332835|graftnull|Transplanted tissue|Anatomy|false|false|C1546653;C1961139;C3683798;C0181074;C1705210|graftnull|Urinary Retention|Finding|false|false|C0042027|urinary retentionnull|Bladder retention of urine|Attribute|false|false|C0042027|urinary retentionnull|Urinary tract|Anatomy|false|false|C0080274;C0149771;C0333117;C0080274;C1753315;C0035280;C0205792;C5700171|urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false|C0042027|retention
null|Retention (Psychology)|Finding|false|false|C0042027|retention
null|Retention of content|Finding|false|false|C0042027|retention
null|cellular entity retention|Finding|false|false|C0042027|retentionnull|Retention - dental|Attribute|false|false||retentionnull|Rectocele|Disorder|false|false|C0042027|rectocelenull|Enterocele|Disorder|false|false|C0042027|enterocelenull|PMH - past medical history|Finding|false|false||Past Medical History
null|Medical History|Finding|false|false||Past Medical Historynull|Medical History|Finding|false|false||Medical Historynull|Medical referral type|Finding|false|false||Medical
null|Medical|Finding|false|false||Medical
null|Medical school type|Finding|false|false||Medicalnull|Medical service|Procedure|false|false||Medicalnull|Medical History|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|History of present illness (finding)|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|cervical cancer|Disorder|false|false|C0027530|Cervical CAnull|Neck|Anatomy|false|false|C4048328|Cervicalnull|Cervical|Modifier|false|false||Cervicalnull|Radical hysterectomy|Procedure|false|false||radical hysterectomynull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Lymphedema|Disorder|false|false||lymphedemanull|Attention deficit hyperactivity disorder|Disorder|false|false||ADHDnull|Anxiety Disorders|Disorder|false|false||Anxiety
null|Anxiety|Disorder|false|false||Anxietynull|Anxiety symptoms|Finding|false|false||Anxietynull|Cancer patients and suicide and depression|Disorder|false|false||Depression
null|Mental Depression|Disorder|false|false||Depression
null|Depressive disorder|Disorder|false|false||Depression
null|Depressed mood|Disorder|false|false||Depressionnull|Depression - motion|Finding|false|false||Depression
null|null|Finding|false|false||Depressionnull|Depression - recess|Modifier|false|false||Depressionnull|Asthma|Disorder|false|false||Asthmanull|Insomnia homeopathic medication|Drug|false|false||Insomnianull|Sleeplessness|Finding|false|false||Insomnianull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Raynaud Disease|Disorder|false|false||Raynaudnull|Ichthyosis Bullosa of Siemens|Disorder|false|false||IBS
null|Irritable Bowel Syndrome|Disorder|false|false||IBSnull|Fibromyalgia|Disorder|false|false||Fibromyalgianull|Social and personal history|Finding|false|false||Social History
null|Social History|Finding|false|false||Social Historynull|Social|Finding|false|false||Socialnull|History of present illness (finding)|Finding|false|false||History
null|History of previous events|Finding|false|false||History
null|Historical aspects qualifier|Finding|false|false||History
null|Medical History|Finding|false|false||History
null|Concept History|Finding|false|false||Historynull|History|Subject|false|false||Historynull|Family Medical History|Finding|false|false||Family Historynull|Entity Name Part Type - family|Finding|false|false||Family
null|Last Name|Finding|false|false||Family
null|Living Arrangement - Family|Finding|false|false||Family
null|Family (taxonomic)|Finding|false|false||Family
null|Family Collection|Finding|false|false||Familynull|Family|Subject|false|false||Familynull|History of present illness (finding)|Finding|false|true||History
null|History of previous events|Finding|false|true||History
null|Historical aspects qualifier|Finding|false|true||History
null|Medical History|Finding|false|true||History
null|Concept History|Finding|false|true||Historynull|History|Subject|false|false||Historynull|Atopy|Finding|false|false||atopy
null|MS4A2 wt Allele|Finding|false|false||atopynull|SON gene|Finding|false|false||sonnull|Son (person)|Subject|false|false||sonnull|Songhay Languages|Entity|false|false||sonnull|Daughter|Subject|false|false||daughternull|Frequently|Time|false|false||frequentnull|Allergy - Charge Type Reason|Finding|false|false||allergy
null|Allergic disposition|Finding|false|false||allergy
null|Hypersensitivity|Finding|false|false||allergy
null|Response to antigens|Finding|false|false||allergy
null|History of allergies|Finding|false|false||allergy
null|Allergic Reaction|Finding|false|false||allergynull|Allergy Specialty|Title|false|false||allergynull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epinull|Exocrine pancreatic insufficiency|Disorder|false|false||epinull|Eysenck personality inventory|Finding|false|false||epi
null|TFPI wt Allele|Finding|false|false||epi
null|TFPI gene|Finding|false|false||epinull|Electronic Portal Imaging|Procedure|false|false||epi
null|Echo-Planar Imaging|Procedure|false|false||epinull|Peripheral Electronic Nerve Stimulation|Procedure|false|false||pensnull|physical examination (physical finding)|Finding|false|false||Physical Examnull|Physical Examination|Procedure|false|false||Physical Examnull|physical examination (physical finding)|Finding|false|false||Physical
null|Physical|Finding|false|false||Physicalnull|Physical Examination|Procedure|false|false||Physicalnull|Exam|Finding|false|false||Examnull|Medical Examination|Procedure|false|false||Examnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|false|false||acute
null|Acute - Triage Code|Finding|false|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Slightly (qualifier value)|Modifier|false|false||slightly
null|Slight (qualifier value)|Modifier|false|false||slightlynull|Muffled voice|Finding|false|false||muffled voicenull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Somewhat|Finding|false|false|C1123023;C4520765|somewhatnull|Flushing|Finding|false|false|C1123023;C4520765|flushed skinnull|Flushing|Finding|false|false|C1123023;C4520765|flushednull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099;C2984079;C0016382;C0016382|skin
null|Skin|Anatomy|false|false|C0178298;C0496955;C1546781;C0444099;C2984079;C0016382;C0016382|skinnull|HEENT|Anatomy|false|false||HEENTnull|Moist mucous membranes|Finding|false|false|C0025255;C0026724|Moist mucous membranesnull|Moist|Modifier|false|false||Moistnull|moisture of mucous membranes (physical finding)|Finding|false|false|C0025255;C0026724|mucous membranesnull|Mucous Membrane|Anatomy|false|false|C0153932;C0264511;C0240211;C1547225;C2230150;C1846919;C3889123;C2753459;C0026727;C0517391|mucous membranesnull|Mucus (substance)|Finding|false|false|C0025255;C0026724|mucous
null|mucus layer|Finding|false|false|C0025255;C0026724|mucousnull|Mucous appearance|Modifier|false|false||mucousnull|Membrane Tissue|Anatomy|false|false|C1846919;C3889123;C2753459;C0026727;C0517391;C2230150;C0240211;C0153932;C0264511;C1547225|membranesnull|Mild Severity of Illness Code|Finding|false|false|C0026724;C0025255|mildnull|Mild (qualifier value)|Modifier|false|false||mild
null|Mild Allergy Severity|Modifier|false|false||mildnull|Lip swelling|Finding|false|false|C0023759;C0026724;C0025255|lip swellingnull|Benign neoplasm of the lip|Disorder|false|false|C0026724;C0025255;C0023759|lip
null|Lymphoid interstitial pneumonia|Disorder|false|false|C0026724;C0025255;C0023759|lipnull|SMG1 wt Allele|Finding|false|false|C0023759;C0025255;C0026724|lip
null|SMG1 gene|Finding|false|false|C0023759;C0025255;C0026724|lipnull|Lip structure|Anatomy|false|false|C1846919;C3889123;C0240211;C0153932;C0264511|lipnull|Swelling|Finding|false|false||swelling
null|Edema|Finding|false|false||swellingnull|Benign neoplasm of tongue|Disorder|false|false|C0040408|tonguenull|Procedure on tongue|Procedure|false|false|C0040408|tonguenull|Tongue|Anatomy|false|false|C0872394;C0153933|tonguenull|Edema|Finding|false|false||edematousnull|Angioedema|Finding|true|false||angioedemanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Jugular venous pressure|Finding|false|false||JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|false|false||wheezesnull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Rhonchi|Finding|false|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Protective muscle spasm|Finding|true|false||guardingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|Peripheral edema|Finding|false|false||edema, peripheralnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Peripheral pulse|Finding|false|false||peripheral pulsesnull|Peripheral|Modifier|false|false||peripheralnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to person|Finding|false|false||oriented to personnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Exam|Finding|false|false||EXAMnull|Medical Examination|Procedure|false|false||EXAMnull|Well (answer to question)|Finding|false|false||Wellnull|Well (container)|Device|false|false||Wellnull|Microplate Well|Modifier|false|false||Well
null|Good|Modifier|false|false||Well
null|Healthy|Modifier|false|false||Wellnull|Females|Subject|false|false||female
null|Woman|Subject|false|false||femalenull|Female, Self-Report|Modifier|false|false||female
null|Female Phenotype|Modifier|false|false||femalenull|patient appears in no acute distress (physical finding)|Finding|false|false||in no acute distressnull|Admission Level of Care Code - Acute|Finding|true|false||acute
null|Acute - Triage Code|Finding|true|false||acutenull|acute|Time|false|false||acutenull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Somewhat|Finding|false|false||somewhatnull|Flushing|Finding|false|false|C1123023;C4520765|flushed skinnull|Flushing|Finding|false|false|C1123023;C4520765|flushednull|Neoplasm of uncertain or unknown behavior of skin|Disorder|false|false|C1123023;C4520765|skin
null|Skin and subcutaneous tissue disorders|Disorder|false|false|C1123023;C4520765|skinnull|Skin Specimen Source Code|Finding|false|false|C1123023;C4520765|skin
null|Skin Specimen|Finding|false|false|C1123023;C4520765|skinnull|Skin, Human|Anatomy|false|false|C1546781;C0444099;C0016382;C0016382;C0178298;C0496955|skin
null|Skin|Anatomy|false|false|C1546781;C0444099;C0016382;C0016382;C0178298;C0496955|skinnull|Prominent|Modifier|false|false||prominentnull|Zygomatic bone|Anatomy|false|false||malarnull|Distribution [PK]|Finding|false|false|C0015450;C4266571|distribution
null|Distribution|Finding|false|false|C0015450;C4266571|distributionnull|Spatial Distribution|Modifier|false|false||distributionnull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C5779816;C1704711;C3160739;C1423759;C2828055;C1414531|face
null|Face|Anatomy|false|false|C5779816;C1704711;C3160739;C1423759;C2828055;C1414531|facenull|Face (spatial concept)|Modifier|false|false||facenull|HEENT|Anatomy|false|false||HEENTnull|Moist mucous membranes|Finding|false|false|C0026724;C0025255|Moist mucous membranesnull|Moist|Modifier|false|false||Moistnull|moisture of mucous membranes (physical finding)|Finding|false|false|C0026724;C0025255|mucous membranesnull|Mucous Membrane|Anatomy|false|false|C0517391;C2230150;C1423759;C2828055;C1414531;C2753459;C0026727;C3160739;C2051406|mucous membranesnull|Mucus (substance)|Finding|false|false|C0025255;C0026724|mucous
null|mucus layer|Finding|false|false|C0025255;C0026724|mucousnull|Mucous appearance|Modifier|false|false||mucousnull|Membrane Tissue|Anatomy|false|false|C3160739;C2753459;C0026727;C2051406;C1423759;C2828055;C1414531;C2230150;C0517391|membranesnull|patient appearance regarding mental status exam|Procedure|false|false|C0025255;C0026724;C0015450;C4266571|appearancenull|null|Attribute|false|false||appearancenull|Personal appearance|Subject|false|false||appearancenull|Appearance|Modifier|false|false||appearancenull|Kind of quantity - Appearance|LabModifier|false|false||appearancenull|FANCONI ANEMIA, COMPLEMENTATION GROUP E|Disorder|false|false|C0025255;C0026724;C0015450;C4266571|facenull|FANCE wt Allele|Finding|false|false|C0026724;C0025255;C0015450;C4266571|face
null|FANCE gene|Finding|false|false|C0026724;C0025255;C0015450;C4266571|face
null|ELOVL6 gene|Finding|false|false|C0026724;C0025255;C0015450;C4266571|facenull|Head>Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C2051406|face
null|Face|Anatomy|false|false|C3160739;C1423759;C2828055;C1414531;C2051406|facenull|Face (spatial concept)|Modifier|false|false||facenull|null|Finding|false|false||unchangednull|About The Same|Modifier|false|false||unchangednull|Benign neoplasm of tongue|Disorder|false|false|C0040408|tonguenull|Procedure on tongue|Procedure|false|false|C0040408|tonguenull|Tongue|Anatomy|false|false|C0153933;C0013604;C0872394|tonguenull|Edema|Finding|true|false|C0040408|edematousnull|Angioedema|Finding|true|false||angioedemanull|Passive joint movement of neck (finding)|Finding|false|false|C0027530;C3159206|Neck
null|Neck problem|Finding|false|false|C0027530;C3159206|Necknull|dendritic spine neck|Anatomy|false|false|C0812434;C0684335|Neck
null|Neck|Anatomy|false|false|C0812434;C0684335|Necknull|Jugular venous pressure|Finding|false|false||JVPnull|Elevated|Modifier|false|false||elevated
null|High|Modifier|false|false||elevatednull|Regular|Modifier|false|false||Regularnull|Amount type - Rate|Finding|false|false||ratenull|Rating (action)|Event|false|false||ratenull|Rate|LabModifier|false|false||ratenull|Rhythm|Finding|false|false||rhythm
null|rhythmic process (biological)|Finding|false|false||rhythmnull|Heart murmur|Finding|true|false||murmursnull|Lung|Anatomy|false|false||Lungsnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Auscultation|Procedure|false|false||auscultationnull|Wheezing|Finding|false|false||wheezesnull|Basilar Rales|Finding|false|false||rales
null|Rales|Finding|false|false||ralesnull|Rhonchi|Finding|false|false||rhonchinull|Malignant neoplasm of abdomen|Disorder|false|false|C0230168;C0000726|Abdomennull|Abdomen problem|Finding|false|false|C0230168;C0000726|Abdomennull|Abdomen|Anatomy|false|false|C0153662;C0941288|Abdomen
null|Abdominal Cavity|Anatomy|false|false|C0153662;C0941288|Abdomennull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||Softnull|Soft|Modifier|false|false||Softnull|Bowel sounds|Finding|false|false|C0021853|bowel soundsnull|Intestines|Anatomy|false|false|C0232693|bowelnull|null|Device|false|false||soundsnull|null|Phenomenon|false|false||soundsnull|Protective muscle spasm|Finding|true|false||guardingnull|Place - dosing instruction imperative|Finding|false|false||placenull|null|Procedure|false|false||placenull|put - instruction imperative|Event|false|false||placenull|Place|Modifier|false|false||placenull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|Feels warm|Finding|false|false||Warmnull|warming process|Phenomenon|false|false||Warmnull|Sequence Chromatogram|Finding|false|false||tracenull|Trace Dosing Unit|LabModifier|false|false||trace
null|trace amount|LabModifier|false|false||trace
null|unknown - trace|LabModifier|false|false||tracenull|Peripheral edema|Finding|false|false||edema, peripheralnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Peripheral pulse|Finding|false|false||peripheral pulsesnull|Peripheral|Modifier|false|false||peripheralnull|null|Drug|false|false||pulsesnull|Physiologic pulse|Finding|false|false||pulsesnull|Pulse taking|Procedure|false|false||pulsesnull|Neurology speciality|Title|false|false||Neuronull|Neurologic (qualifier value)|Modifier|false|false||Neuronull|Alert brand of caffeine|Drug|false|false||alert
null|Alert brand of caffeine|Drug|false|false||alertnull|Mentally alert|Finding|false|false||alert
null|Consciousness clear|Finding|false|false||alert
null|Alert note|Finding|false|false||alert
null|Alert|Finding|false|false||alertnull|null|Attribute|false|false||alertnull|Oriented to person|Finding|false|false||oriented to personnull|Oriented to place|Finding|false|false||orientednull|Orientation, Spatial|Modifier|false|false||orientednull|Person Info|Finding|false|false||personnull|null|Attribute|false|false||personnull|Persons|Subject|false|false||personnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Gynecology|Title|false|false||GYNnull|Gynecologic|Modifier|false|false||GYNnull|Floor (anatomic)|Anatomy|false|false|C0030685;C0582103;C4284036;C0600083;C1546601;C0012621;C2926602|Floornull|floor (object)|Device|false|false||Floornull|Floor - story of building|Entity|false|false||Floornull|Body Substance Discharge|Finding|false|false|C3714591|discharge
null|Discharge Body Fluid|Finding|false|false|C3714591|discharge
null|Body Fluid Discharge|Finding|false|false|C3714591|discharge
null|null|Finding|false|false|C3714591|dischargenull|Patient Discharge|Procedure|false|false|C3714591|dischargenull|Exam|Finding|false|false|C3714591|examnull|Medical Examination|Procedure|false|false|C3714591|examnull|United States Military Commissioned Officer O10 (qualifier value)|Finding|false|false||Gen
null|GEN1 wt Allele|Finding|false|false||Gen
null|GEN1 gene|Finding|false|false||Gennull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Respiratory, thoracic and mediastinal disorders|Disorder|false|false||Respnull|Respiratory rate|Attribute|false|false||Respnull|Visible|Modifier|false|false||visiblenull|Respiratory distress|Finding|true|false||respiratory distressnull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|Emotional distress|Finding|true|false||distress
null|Distress|Finding|true|false||distressnull|Full|Modifier|false|false||fullnull|Sentence|Finding|false|false||sentencesnull|Absence of Biallelic TCRgamma Deletion|Disorder|false|false|C0449202;C0000726|Abdnull|ABD (body structure)|Anatomy|false|false|C3811055|Abd
null|Abdomen|Anatomy|false|false|C3811055|Abdnull|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Disorder|false|false||softnull|Soft|Modifier|false|false||softnull|Hereditary Multiple Exostoses|Disorder|false|false||Extnull|EXT1 wt Allele|Finding|false|false||Ext
null|EXT1 gene|Finding|false|false||Extnull|All extremities|Anatomy|false|false||extremities
null|Limb structure|Anatomy|false|false||extremitiesnull|Admission activity|Procedure|false|false||ADMISSION
null|Hospital admission|Procedure|false|false||ADMISSIONnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood tryptase|Procedure|false|false||BLOOD TRYPTASEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|TRYPTASE|Drug|false|false||TRYPTASE
null|TRYPTASE|Drug|false|false||TRYPTASEnull|Tryptase measurement|Procedure|false|false||TRYPTASEnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Body Substance Discharge|Finding|false|false||DISCHARGE
null|Discharge Body Fluid|Finding|false|false||DISCHARGE
null|Body Fluid Discharge|Finding|false|false||DISCHARGE
null|null|Finding|false|false||DISCHARGEnull|Patient Discharge|Procedure|false|false||DISCHARGEnull|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C0014792;C1114281|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|MCOLN1 protein, human|Drug|false|false||Mg-2
null|MCOLN1 protein, human|Drug|false|false||Mg-2null|MCOLN1 wt Allele|Finding|false|false||Mg-2null|Laboratory test finding|Lab|false|false||LABSnull|Blood and lymphatic system disorders|Disorder|false|false|C0023516|BLOODnull|peripheral blood|Finding|false|false|C0023516|BLOOD
null|Blood|Finding|false|false|C0023516|BLOOD
null|In Blood|Finding|false|false|C0023516|BLOODnull|Leukocytes|Anatomy|false|false|C0851353;C0005768;C0229664;C0005767|WBCnull|Erythrocytes|Drug|false|false|C0014792|RBCnull|Erythrocytes|Anatomy|false|false|C1114281;C0014792|RBCnull|null|Attribute|false|false|C0014792|RBCnull|Hemoglobin|Drug|false|false||Hgb
null|Hemoglobin|Drug|false|false||Hgbnull|CYGB gene|Finding|false|false||Hgbnull|Hemoglobin concentration|Lab|false|false||Hgbnull|Hemopoietic stem cell transplant|Procedure|false|false||Hct
null|Hematocrit Measurement|Procedure|false|false||Hctnull|Merkel cell polyomavirus|Disorder|false|false||MCVnull|Erythrocyte Mean Corpuscular Volume Measurement|Procedure|false|false||MCV
null|Cisplatin-Methotrexate-Vinblastine Regimen|Procedure|false|false||MCVnull|Mean Corpuscular Volume|Lab|false|false||MCVnull|Microvolt|LabModifier|false|false||MCVnull|methacholine|Drug|false|false||MCH
null|methacholine|Drug|false|false||MCHnull|mesaconyl-CoA hydratase activity|Finding|false|false||MCH
null|PMCH gene|Finding|false|false||MCHnull|Mean corpuscular hemoglobin determination|Procedure|false|false||MCHnull|Mean corpuscular hemoglobin concentration determination|Procedure|false|false||MCHCnull|Primed lymphocyte test|Procedure|false|false||Pltnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Lymph|Finding|false|false||Lymphsnull|Monos|Drug|false|false||Monos
null|Mono-S|Drug|false|false||Monos
null|Monos|Drug|false|false||Monosnull|SARCOIDOSIS, EARLY-ONSET|Disorder|false|false||Eos
null|Familial eosinophilia|Disorder|false|false||Eosnull|PRSS33 gene|Finding|false|false||Eos
null|IKZF4 gene|Finding|false|false||Eosnull|Eos <Loriini>|Entity|false|false||Eosnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|Proliferating trichilemmal tumor|Disorder|false|false||PTTnull|Partial thromboplastin time, activated (procedure)|Procedure|false|false||PTT
null|Partial Thromboplastin Time|Procedure|false|false||PTTnull|Blood Glucose|Drug|false|false||BLOOD Glucosenull|Blood glucose measurement|Procedure|false|false||BLOOD Glucosenull|Finding of blood glucose level|Lab|false|false||BLOOD Glucosenull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucose
null|glucose|Drug|false|false||Glucosenull|Glucose measurement|Procedure|false|false||Glucosenull|Glucose^1.5H post dose glucagon|Lab|false|false||Glucosenull|Bicarbonates|Drug|false|false||HCO3
null|Bicarbonates|Drug|false|false||HCO3null|Bicarbonate measurement|Procedure|false|false||HCO3null|Blood calcium measurement|Procedure|false|false||BLOOD Calciumnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|calcium|Drug|false|false||Calcium
null|CALCIUM SUPPLEMENTS|Drug|false|false||Calcium
null|Calcium, Dietary|Drug|false|false||Calcium
null|Calcium [EPC]|Drug|false|false||Calcium
null|Calcium Drug Class|Drug|false|false||Calciumnull|Calcium metabolic function|Finding|false|false||Calciumnull|Calcium measurement|Procedure|false|false||Calciumnull|Phos <Photinae>|Entity|false|false||Phosnull|Blood tryptase|Procedure|false|false||BLOOD TRYPTASEnull|Blood and lymphatic system disorders|Disorder|false|false||BLOODnull|peripheral blood|Finding|false|false||BLOOD
null|Blood|Finding|false|false||BLOOD
null|In Blood|Finding|false|false||BLOODnull|TRYPTASE|Drug|false|false||TRYPTASE
null|TRYPTASE|Drug|false|false||TRYPTASEnull|Tryptase measurement|Procedure|false|false||TRYPTASEnull|Paroxysmal nocturnal dyspnea|Disorder|false|false||PNDnull|NPPA wt Allele|Finding|false|false||PND
null|NPPA gene|Finding|false|false||PNDnull|Imaging problem|Finding|false|false||IMAGINGnull|Diagnostic Imaging|Procedure|false|false||IMAGING
null|Imaging Techniques|Procedure|false|false||IMAGINGnull|Imaging Technology|Title|false|false||IMAGINGnull|Micro (prefix)|Finding|false|false||MICRO
null|Microbiology - Laboratory Class|Finding|false|false||MICROnull|Microbiology procedure|Procedure|false|false||MICROnull|Unit Of Measure Prefix - micro|LabModifier|false|false||MICROnull|BRIEF Health Literacy Screening Tool|Finding|false|false||Brief
null|Behavior Rating Inventory of Executive Function|Finding|false|false||Briefnull|Brief|Time|false|false||Briefnull|Shortened|Modifier|false|false||Briefnull|Hospital course|Finding|false|false||Hospital Coursenull|null|Attribute|false|false||Hospital Coursenull|Organization unit type - Hospital|Finding|false|false||Hospitalnull|Hospitals|Device|false|false||Hospitalnull|Hospitals|Entity|false|false||Hospitalnull|Hospital environment|Modifier|false|false||Hospitalnull|Course|Time|false|false||Coursenull|cervical cancer|Disorder|false|false|C0027530|cervical CAnull|Neck|Anatomy|false|false|C4048328|cervicalnull|Cervical|Modifier|false|false||cervicalnull|Radicals (chemistry)|Drug|false|false||radicalnull|Radical (qualifier value)|Modifier|false|false||radicalnull|Consent Type - Hysterectomy|Finding|false|false||hysterectomynull|Hysterectomy|Procedure|false|false||hysterectomynull|Chronic - Admission Level of Care Code|Finding|false|false||chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||chronicnull|chronic|Time|false|false||chronicnull|Lymphedema|Disorder|false|false||lymphedemanull|Urinary Retention|Finding|false|false|C0042027|urinary retentionnull|Bladder retention of urine|Attribute|false|false||urinary retentionnull|Urinary tract|Anatomy|false|false|C0080274|urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Retention of content|Finding|false|false||retention
null|cellular entity retention|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Asthma|Disorder|false|false||Asthmanull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Fibromyalgia|Disorder|false|false||fibromyalgianull|Operative report|Finding|false|false||operative reportnull|Operative|Time|false|false||operativenull|Report (document)|Finding|false|false||reportnull|Reporting|Procedure|false|false||reportnull|null|Attribute|false|false||reportnull|Full|Modifier|false|false||fullnull|Details|Modifier|false|false||detailsnull|Postoperative Period|Time|false|false||post-operativenull|Course|Time|false|false||coursenull|Uncomplicated|Modifier|false|false||uncomplicatednull|Stat (do immediately)|Time|false|false||Immediatelynull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Toradol|Drug|false|false||toradol
null|Toradol|Drug|false|false||toradolnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Pruritus|Finding|false|false||itchynull|Once - dosing instruction fragment|Finding|false|false||Oncenull|Once (schedule frequency)|Time|false|false||Oncenull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Observation of Sensation|Finding|false|false|C0040408|sensation
null|Sensory perception|Finding|false|false|C0040408|sensationnull|sensory exam|Procedure|false|false|C0040408|sensationnull|Sensation quality|Modifier|false|false||sensationnull|Benign neoplasm of tongue|Disorder|false|false|C0040408|tonguenull|Procedure on tongue|Procedure|false|false|C0040408|tonguenull|Tongue|Anatomy|false|false|C0153933;C2229507;C0036658;C0542538;C0872394|tonguenull|Lip swelling|Finding|false|false|C0023759|lip swellingnull|Benign neoplasm of the lip|Disorder|false|false|C0023759|lip
null|Lymphoid interstitial pneumonia|Disorder|false|false|C0023759|lipnull|SMG1 wt Allele|Finding|false|false|C0023759|lip
null|SMG1 gene|Finding|false|false|C0023759|lipnull|Lip structure|Anatomy|false|false|C0240211;C0392747;C1846919;C3889123;C0036537;C0153932;C0264511;C0013604;C0038999;C4319952;C1299586|lipnull|Swelling|Finding|false|false|C0023759|swelling
null|Edema|Finding|false|false|C0023759|swellingnull|Has difficulty doing (qualifier value)|Finding|false|false|C0023759|difficultynull|Bodily secretions|Finding|false|false|C0023759|secretionsnull|Changing|Finding|false|false||change innull|Changed status|LabModifier|false|false||change innull|Changing|Finding|false|false|C0023759|changenull|Change - procedure|Procedure|false|false|C0023759|changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Dyspnea|Finding|true|false||SOBnull|Flushing|Finding|true|false||flushingnull|Stridor|Finding|true|false||stridornull|Wheezing|Finding|true|false||wheezenull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|penclomedine|Drug|false|false||pen
null|penclomedine|Drug|false|false||pennull|TSPAN33 gene|Finding|false|false||pen
null|PUM3 gene|Finding|false|false||pen
null|PCSK1N gene|Finding|false|false||pennull|Pre-filled Pen Syringe|Device|false|false||pennull|Pen (unit of presentation)|LabModifier|false|false||pennull|Solu-Medrol|Drug|false|false||Solumedrol
null|Solu-Medrol|Drug|false|false||Solumedrolnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|hydroxyzine|Drug|false|false||Hydroxyzine
null|hydroxyzine|Drug|false|false||Hydroxyzinenull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Has patient|Finding|false|false||patient hasnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Numerous|LabModifier|false|false||numerousnull|Drug Allergy|Finding|false|false||drug allergiesnull|Pharmaceutical Preparations|Drug|false|false||drug
null|Pharmacologic Substance|Drug|false|false||drugnull|Drug problem|Finding|false|false||drugnull|Hypersensitivity|Finding|false|false||allergiesnull|null|Attribute|false|false||allergiesnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|midazolam|Drug|false|false||Midazolam
null|midazolam|Drug|false|false||Midazolamnull|rocuronium|Drug|false|false||Rocuronium
null|rocuronium|Drug|false|false||Rocuroniumnull|fentanyl|Drug|false|false||Fentanyl
null|fentanyl|Drug|false|false||Fentanylnull|Fentanyl measurement|Procedure|false|false||Fentanylnull|dexamethasone|Drug|false|false||Dexamethasone
null|dexamethasone|Drug|false|false||Dexamethasonenull|hydromorphone|Drug|false|false||Hydromorphone
null|hydromorphone|Drug|false|false||Hydromorphonenull|ondansetron|Drug|false|false||Ondansetron
null|ondansetron|Drug|false|false||Ondansetronnull|lidocaine|Drug|false|false||Lidocaine
null|lidocaine|Drug|false|false||Lidocainenull|Lidocaine measurement|Procedure|false|false||Lidocainenull|propofol|Drug|false|false||Propofol
null|propofol|Drug|false|false||Propofolnull|cefazolin|Drug|false|false||Cefazolin
null|cefazolin|Drug|false|false||Cefazolinnull|glycopyrrolate|Drug|false|false||Glycopyrrolate
null|glycopyrrolate|Drug|false|false||Glycopyrrolatenull|phenylephrine|Drug|false|false||Phenylephrine
null|phenylephrine|Drug|false|false||Phenylephrinenull|ketorolac|Drug|false|false||Ketorolac
null|ketorolac|Drug|false|false||Ketorolacnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|BP 100|Drug|false|false||BP 100
null|BP 100|Drug|false|false||BP 100null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Wheezing|Finding|true|false||wheezenull|Patient Condition Code - Poor|Finding|true|false||poor
null|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|true|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Air (substance)|Drug|true|false||air
null|air|Drug|true|false||air
null|air|Drug|true|false||airnull|ACUTE INSULIN RESPONSE|Finding|true|false||air
null|AIRN gene|Finding|true|false||air
null|AI/RHEUM|Finding|true|false||airnull|Movement|Finding|false|false||movementnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Persistent|Time|false|false||persistentnull|Dysphonia|Disorder|false|false||voice changenull|Change in voice (finding)|Finding|false|false||voice changenull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|More|LabModifier|false|false||morenull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epinull|Exocrine pancreatic insufficiency|Disorder|false|false||epinull|Eysenck personality inventory|Finding|false|false||epi
null|TFPI wt Allele|Finding|false|false||epi
null|TFPI gene|Finding|false|false||epinull|Electronic Portal Imaging|Procedure|false|false||epi
null|Echo-Planar Imaging|Procedure|false|false||epinull|Peripheral Electronic Nerve Stimulation|Procedure|false|false||pensnull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|compromise|Finding|false|false||compromisenull|post operative (finding)|Finding|false|false||Post operativenull|SLC35G1 gene|Finding|false|false||Post
null|DESI1 gene|Finding|false|false||Postnull|Post Device|Device|false|false||Postnull|Post|Time|false|false||Postnull|Operative|Time|false|false||operativenull|In care (finding)|Finding|false|false||care
null|Continuity Assessment Record and Evaluation|Finding|false|false||carenull|care activity|Event|false|false||carenull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Stat (do immediately)|Time|false|false||immediatelynull|Dilaudid|Drug|false|false||dilaudid
null|Dilaudid|Drug|false|false||dilaudidnull|Toradol|Drug|false|false||toradol
null|Toradol|Drug|false|false||toradolnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Difficult (qualifier value)|Finding|false|false||difficultnull|Allergic Reaction|Finding|false|false||allergic reaction
null|Hypersensitivity|Finding|false|false||allergic reactionnull|Allergic|Finding|false|false||allergicnull|Reaction|Finding|false|false||reactionnull|Insertion of pack into vagina|Procedure|false|false|C0042232|vaginal packingnull|Vaginal Dosage Form|Drug|false|false|C0042232|vaginalnull|Vaginal Route of Administration|Finding|false|false|C0042232|vaginal
null|Vaginal (intended site)|Finding|false|false|C0042232|vaginalnull|Vagina|Anatomy|false|false|C1272941;C4521343;C1522570;C0184967;C1270937|vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Packing Dosage Form|Drug|false|false||packingnull|Insertion of pack (procedure)|Procedure|false|false|C0042232|packingnull|Packing material|Device|false|false||packingnull|Packing (action)|Event|false|false||packingnull|Postoperative Period|Time|false|false||post-operativenull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|monitoring of urine output for fluid balance|Procedure|false|false||urine outputnull|null|Attribute|false|false||urine output
null|null|Attribute|false|false||urine outputnull|Urine volume finding|LabModifier|false|false||urine outputnull|Portion of urine|Finding|false|false||urine
null|null|Finding|false|false||urine
null|Urine|Finding|false|false||urine
null|In Urine|Finding|false|false||urine
null|Urine specimen|Finding|false|false||urinenull|system output|Finding|false|false||outputnull|Measurement of fluid output|Procedure|false|false||outputnull|Adequate|Modifier|false|false||adequate
null|Sufficient|Modifier|false|false||adequatenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Able (qualifier value)|Finding|false|false||ablenull|Ability|Subject|false|false||ablenull|subscriber - self|Finding|false|false||self
null|Self|Finding|false|false||selfnull|Catheterization|Procedure|false|false||catheterizationnull|TELANGIECTASIA, IMPAIRED INTELLECTUAL DEVELOPMENT, MICROCEPHALY, METAPHYSEAL DYSPLASIA, EYE ABNORMALITIES, AND SHORT STATURE|Disorder|false|false||timesnull|Time|Time|false|false||timesnull|Times|LabModifier|false|false||timesnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Observation of Sensation|Finding|false|false||sensation
null|Sensory perception|Finding|false|false||sensationnull|sensory exam|Procedure|false|false||sensationnull|Sensation quality|Modifier|false|false||sensationnull|Neoplasm of uncertain or unknown behavior of bladder|Disorder|false|false|C0005682|bladder
null|Benign neoplasm of bladder|Disorder|false|false|C0005682|bladder
null|Carcinoma in situ of bladder|Disorder|false|false|C0005682|bladdernull|Procedures on bladder|Procedure|false|false|C0005682|bladdernull|Urinary Bladder|Anatomy|false|false|C0496930;C0154017;C0154091;C0872388|bladdernull|Fullness|Modifier|false|false||fullnessnull|Anaphylaxis;non medication|Disorder|false|false||Anaphylaxisnull|anaphylaxis|Finding|false|false||Anaphylaxis
null|Anaphylactic shock|Finding|false|false||Anaphylaxisnull|Recovery Room|Device|false|false||PACUnull|Recovery Room|Entity|false|false||PACUnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Pruritus|Finding|false|false||pruritisnull|Once - dosing instruction fragment|Finding|false|false||Oncenull|Once (schedule frequency)|Time|false|false||Oncenull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Lip swelling|Finding|false|false|C0023759|swollen lipsnull|Swelling|Finding|false|false||swollennull|Lip structure|Anatomy|false|false|C0240211;C0872394;C0205382;C0153933|lipsnull|Benign neoplasm of tongue|Disorder|false|false|C0040408;C0023759|tonguenull|Procedure on tongue|Procedure|false|false|C0040408;C0023759|tonguenull|Tongue|Anatomy|false|false|C0872394;C0153933|tonguenull|vocal|Finding|false|false|C0023759|vocalnull|Changing|Finding|false|false||changesnull|Changed status|LabModifier|false|false||changesnull|Dyspnea|Finding|true|false||SOBnull|Flushing|Finding|false|false||flushingnull|Stridor|Finding|true|false||stridornull|Wheezing|Finding|true|false||wheezenull|Precipitating Factors|Attribute|false|false||triggernull|Triggered by|Modifier|false|false||triggernull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|penclomedine|Drug|false|false||pen
null|penclomedine|Drug|false|false||pennull|TSPAN33 gene|Finding|false|false||pen
null|PUM3 gene|Finding|false|false||pen
null|PCSK1N gene|Finding|false|false||pennull|Pre-filled Pen Syringe|Device|false|false||pennull|Pen (unit of presentation)|LabModifier|false|false||pennull|Solu-Medrol|Drug|false|false||Solumedrol
null|Solu-Medrol|Drug|false|false||Solumedrolnull|famotidine|Drug|false|false||Famotidine
null|famotidine|Drug|false|false||Famotidinenull|hydroxyzine|Drug|false|false||Hydroxyzine
null|hydroxyzine|Drug|false|false||Hydroxyzinenull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Initial (abbreviation)|Finding|false|false||initialnull|Initially|Time|false|false||initialnull|Firstly|Modifier|false|false||initialnull|BP 100|Drug|false|false||BP 100
null|BP 100|Drug|false|false||BP 100null|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|nicotinamide adenine dinucleotide (NAD)|Drug|false|false||NAD
null|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide|Drug|false|false||NADnull|NEUTROPHIL ACTIN DYSFUNCTION|Disorder|false|false||NAD
null|Dysplastic Nevus|Disorder|false|false||NAD
null|Neuroaxonal Dystrophies|Disorder|false|false||NADnull|patient appears in no acute distress (physical finding)|Finding|false|false||NADnull|Wheezing|Finding|true|false||wheezenull|Patient Condition Code - Poor|Finding|true|false||poor
null|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group|Finding|true|false||poornull|Poverty|Subject|false|false||poornull|Language Proficiency - Poor|Modifier|false|false||poor
null|Specimen Quality - Poor|Modifier|false|false||poor
null|Poor - grade|Modifier|false|false||poor
null|Poor - qualifier|Modifier|false|false||poornull|Air (substance)|Drug|true|false||air
null|air|Drug|true|false||air
null|air|Drug|true|false||airnull|ACUTE INSULIN RESPONSE|Finding|true|false||air
null|AIRN gene|Finding|true|false||air
null|AI/RHEUM|Finding|true|false||airnull|Movement|Finding|false|false||movementnull|Exam|Finding|false|false||examnull|Medical Examination|Procedure|false|false||examnull|Persistent|Time|false|false||persistentnull|Dysphonia|Disorder|false|false||voice changenull|Change in voice (finding)|Finding|false|false||voice changenull|Authorization Mode - Voice|Finding|false|false||voice
null|Voice G-code|Finding|false|false||voice
null|Voice|Finding|false|false||voicenull|TelecommunicationCapabilities - voice|Modifier|false|false||voicenull|Changing|Finding|false|false||changenull|Change - procedure|Procedure|false|false||changenull|Delta (difference)|LabModifier|false|false||change
null|Changed status|LabModifier|false|false||changenull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|More|LabModifier|false|false||morenull|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|epinephrine|Drug|false|false||epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||epinull|Exocrine pancreatic insufficiency|Disorder|false|false||epinull|Eysenck personality inventory|Finding|false|false||epi
null|TFPI wt Allele|Finding|false|false||epi
null|TFPI gene|Finding|false|false||epinull|Electronic Portal Imaging|Procedure|false|false||epi
null|Echo-Planar Imaging|Procedure|false|false||epinull|Peripheral Electronic Nerve Stimulation|Procedure|false|false||pensnull|Hemodynamically stable|Finding|false|false||hemodynamically stablenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|compromise|Finding|false|false||compromisenull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Feeling comfortable|Finding|false|false||comfortablenull|BORNHOLM EYE DISEASE|Disorder|false|false||bednull|Bachelor of Education|Finding|false|false||bednull|Beds|Device|false|false||bednull|Patient Location - Bed|Modifier|false|false||bednull|More|LabModifier|false|false||morenull|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|epinephrine|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epi
null|Tissue Factor Pathway Inhibitor, human|Drug|false|false||Epinull|Exocrine pancreatic insufficiency|Disorder|false|false||Epinull|Eysenck personality inventory|Finding|false|false||Epi
null|TFPI wt Allele|Finding|false|false||Epi
null|TFPI gene|Finding|false|false||Epinull|Electronic Portal Imaging|Procedure|false|false||Epi
null|Echo-Planar Imaging|Procedure|false|false||Epinull|Peripheral Electronic Nerve Stimulation|Procedure|false|false||pensnull|epinephrine|Drug|false|false||epinephrine
null|epinephrine|Drug|false|false||epinephrine
null|epinephrine|Drug|false|false||epinephrinenull|Epinephrine measurement|Procedure|false|false||epinephrinenull|Drops - Drug Form|Drug|false|false||gttnull|Gestational Trophoblastic Neoplasms|Disorder|false|false||gttnull|Glucose tolerance test|Procedure|false|false||gttnull|Drop Dosing Unit|LabModifier|false|false||gtt
null|Medical Drop|LabModifier|false|false||gttnull|Feeling comfortable|Finding|false|false||comfortablenull|Cell Respiration|Finding|false|false||respiration
null|Respiration|Finding|false|false||respirationnull|respiratory system process|Phenomenon|false|false||respirationnull|Vocalization (finding)|Finding|false|false||vocalizationnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|oralnull|Oral|Modifier|false|false||oralnull|Structure|Modifier|false|false||structuresnull|Ativan|Drug|false|false||Ativan
null|Ativan|Drug|false|false||Ativannull|Ambien|Drug|false|false||Ambien
null|Ambien|Drug|false|false||Ambiennull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|propranolol|Drug|false|false||propranolol
null|propranolol|Drug|false|false||propranololnull|Essential Tremor|Disorder|false|false||essential tremornull|Essential|Modifier|false|false||essentialnull|Tremor|Finding|false|false||tremornull|Explanation|Finding|false|false||explanationnull|Adrenergic beta-Antagonists|Drug|false|false||beta blockersnull|Greek letter beta|Finding|false|false||betanull|Beta <eudicots>|Entity|false|false||betanull|Beta Distribution|LabModifier|false|false||betanull|Bronchoconstriction [PE]|Finding|false|false||bronchoconstriction
null|Bronchoconstriction|Finding|false|false||bronchoconstrictionnull|Respiratory compromise|Finding|false|false||respiratory compromisenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|compromise|Finding|false|false||compromisenull|Anaphylaxis;non medication|Disorder|false|false||anaphylaxisnull|anaphylaxis|Finding|false|false||anaphylaxis
null|Anaphylactic shock|Finding|false|false||anaphylaxisnull|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|Floor (anatomic)|Anatomy|false|false||floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Persistent|Time|false|false||persistentnull|Flushing|Finding|false|false|C0015450|facial flushing
null|Face goes red|Finding|false|false|C0015450|facial flushingnull|Face|Anatomy|false|false|C5848177;C0016382;C0016382|facialnull|Facial|Modifier|false|false||facialnull|Flushing|Finding|false|false|C0015450|flushingnull|Apyrexial|Finding|false|false||afebrilenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Respiratory compromise|Finding|true|false||respiratory compromisenull|Respiratory attachment|Finding|false|false||respiratory
null|respiratory|Finding|false|false||respiratory
null|null|Finding|false|false||respiratory
null|Respiratory specimen|Finding|false|false||respiratorynull|Respiratory rate|Attribute|false|false||respiratorynull|compromise|Finding|true|false||compromisenull|systemic symptoms|Finding|true|false||systemic symptomsnull|Systemic Route of Administration|Finding|false|false||systemic
null|Systemic|Finding|false|false||systemicnull|Symptoms aspect|Finding|false|false||symptoms
null|Symptoms|Finding|false|false||symptomsnull|Symptomatic|Finding|false|false||Symptomaticnull|Continuity Assessment Record and Evaluation|Finding|false|false||care
null|In care (finding)|Finding|false|false||carenull|care activity|Event|false|false||carenull|hydroxyzine|Drug|false|false||hydroxyzine
null|hydroxyzine|Drug|false|false||hydroxyzinenull|eucerin|Drug|false|false||eucerin
null|eucerin|Drug|false|false||eucerinnull|Lotion|Drug|false|false||lotionnull|Step (specific stage)|Finding|false|false|C3714591|step
null|Treatment Step|Finding|false|false|C3714591|step
null|PTPN5 gene|Finding|false|false|C3714591|stepnull|Stair (equipment)|Device|false|false||stepnull|Increment|LabModifier|false|false||stepnull|Floor (anatomic)|Anatomy|false|false|C1261552;C1419107;C1704379|floornull|floor (object)|Device|false|false||floornull|Floor - story of building|Entity|false|false||floornull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Breast Feeding|Finding|false|false||nursingnull|RNAx nursing therapy actions|Procedure|false|false||nursingnull|Discipline of Nursing|Title|false|false||nursingnull|Constriction in throat|Finding|false|false|C0230069;C3665375;C0031354;C1760025|throat constrictionnull|Throat Homeopathic Medication|Drug|false|false|C0230069;C3665375;C0031354|throatnull|Specimen Type - Throat|Finding|false|false|C0230069;C3665375;C0031354;C1760025|throat
null|null|Finding|false|false|C0230069;C3665375;C0031354;C1760025|throatnull|Throat|Anatomy|false|false|C0236071;C0009813;C1550663;C1547926;C1950455;C1261287|throat
null|Anterior portion of neck|Anatomy|false|false|C0236071;C0009813;C1550663;C1547926;C1950455;C1261287|throat
null|Pharyngeal structure|Anatomy|false|false|C0236071;C0009813;C1550663;C1547926;C1950455;C1261287|throatnull|Stenosis|Finding|false|false|C0230069;C3665375;C0031354;C1760025|constrictionnull|Constriction procedure|Procedure|false|false|C0230069;C3665375;C0031354;C1760025|constrictionnull|constriction location|Anatomy|false|false|C0236071;C0009813;C1550663;C1547926;C1261287|constrictionnull|LOOP,CONSTRICTION ADJUSTABLE DEVICE ACTIS|Device|false|false||constrictionnull|epinephrine|Drug|false|false||Epinephrine
null|epinephrine|Drug|false|false||Epinephrine
null|epinephrine|Drug|false|false||Epinephrinenull|Epinephrine measurement|Procedure|false|false||Epinephrinenull|Solu-Medrol|Drug|false|false||solumedrol
null|Solu-Medrol|Drug|false|false||solumedrolnull|Relationship modifier - Patient|Finding|false|false||patient
null|Specimen Type - Patient|Finding|false|false||patient
null|Mail Claim Party - Patient|Finding|false|false||patient
null|Report source - Patient|Finding|false|false||patient
null|null|Finding|false|false||patient
null|Disabled Person Code - Patient|Finding|false|false||patientnull|Patients|Subject|false|false||patientnull|Veterinary Patient|Entity|false|false||patientnull|Relief brand of phenylephrine|Drug|false|false||relief
null|Relief brand of phenylephrine|Drug|false|false||reliefnull|Feeling relief|Finding|false|false||reliefnull|Allergy - Charge Type Reason|Finding|false|false||Allergy
null|Allergic disposition|Finding|false|false||Allergy
null|Hypersensitivity|Finding|false|false||Allergy
null|Response to antigens|Finding|false|false||Allergy
null|History of allergies|Finding|false|false||Allergy
null|Allergic Reaction|Finding|false|false||Allergynull|Allergy Specialty|Title|false|false||Allergynull|New medications|Drug|false|false||new medicationsnull|Query Status Code - new|Finding|false|false||new
null|Act Status - new|Finding|false|false||newnull|Newar Language|Entity|false|false||newnull|New|Modifier|false|false||newnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Organization unit type - Hospital|Finding|false|false||hospitalnull|Hospitals|Device|false|false||hospitalnull|Hospitals|Entity|false|false||hospitalnull|Hospital environment|Modifier|false|false||hospitalnull|Hypersensitivity|Finding|false|false||allergiesnull|null|Attribute|false|false||allergiesnull|In addition to|Finding|false|false||addition
null|Add - instruction imperative|Finding|false|false||additionnull|TRYPTASE|Drug|false|false||tryptase
null|TRYPTASE|Drug|false|false||tryptasenull|Tryptase measurement|Procedure|false|false||tryptasenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Chronic - Admission Level of Care Code|Finding|false|false||Chronicnull|Provision of recurring care for chronic illness|Procedure|false|false||Chronicnull|chronic|Time|false|false||Chronicnull|Edema|Finding|false|false||edemanull|null|Attribute|false|false||edemanull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|metolazone|Drug|false|false||Metolazone
null|metolazone|Drug|false|false||Metolazonenull|spironolactone|Drug|false|false||spironolactone
null|spironolactone|Drug|false|false||spironolactonenull|Potassium Drug Class|Drug|false|false||potassium
null|Dietary Potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|potassium|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassium
null|Potassium supplement|Drug|false|false||potassiumnull|Potassium metabolic function|Finding|false|false||potassiumnull|Potassium measurement|Procedure|false|false||potassiumnull|Hypotensive|Finding|false|false||hypotensivenull|Asthma|Disorder|false|false||Asthmanull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Use - dosing instruction imperative|Finding|false|false||use
null|utilization qualifier|Finding|false|false||use
null|Usage|Finding|false|false||usenull|Weekly|Time|false|false||per weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Gastroesophageal reflux disease|Disorder|false|false||GERDnull|Nexium|Drug|false|false||Nexium
null|Nexium|Drug|false|false||Nexiumnull|Initially|Time|false|false||initiallynull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Request - ActReason|Finding|false|false||request
null|request - ActMood|Finding|false|false||request
null|Question (inquiry)|Finding|false|false||requestnull|null|Event|false|false||requestnull|null|Time|false|false||prior tonull|null|Time|false|false||priornull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Attention deficit hyperactivity disorder|Disorder|false|false||ADHDnull|Adderall|Drug|false|false||Adderall
null|Adderall|Drug|false|false||Adderallnull|On admission|Time|false|false||on admissionnull|Admission activity|Procedure|false|false||admission
null|Hospital admission|Procedure|false|false||admissionnull|Anxiety Disorders|Disorder|false|false||Anxiety
null|Anxiety|Disorder|false|false||Anxietynull|Anxiety symptoms|Finding|false|false||Anxietynull|Cancer patients and suicide and depression|Disorder|false|false||depression
null|Mental Depression|Disorder|false|false||depression
null|Depressive disorder|Disorder|false|false||depression
null|Depressed mood|Disorder|false|false||depressionnull|Depression - motion|Finding|false|false||depression
null|null|Finding|false|false||depressionnull|Depression - recess|Modifier|false|false||depressionnull|Fibromyalgia|Disorder|false|false||fibromyalgianull|lorazepam|Drug|false|false||lorazepam
null|lorazepam|Drug|false|false||lorazepamnull|Insomnia homeopathic medication|Drug|false|false||Insomnianull|Sleeplessness|Finding|false|false||Insomnianull|zolpidem|Drug|false|false||zolpidem
null|zolpidem|Drug|false|false||zolpidemnull|Postoperative Period|Time|false|false||post-operativenull|Day 1|Time|false|false||day 1null|Transaction counts and value totals - day|Finding|false|false||day
null|Precision - day|Finding|false|false||daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Oral Dosage Form|Drug|false|false|C0226896|oralnull|Oral Route of Administration|Finding|false|false|C0226896|oral
null|Oral (intended site)|Finding|false|false|C0226896|oralnull|Oral cavity|Anatomy|false|false|C1527415;C4521986;C1272919|oralnull|Oral|Modifier|false|false||oralnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Referral category - Outpatient|Finding|false|false||outpatient
null|Patient Class - Outpatient|Finding|false|false||outpatientnull|Outpatients|Subject|false|false||outpatientnull|Follow-up status|Finding|false|false||follow-upnull|follow-up|Procedure|false|false||follow-upnull|Follow - dosing instruction imperative|Finding|false|false||follow
null|Follow|Finding|false|false||follownull|Followed by|Time|false|false||follownull|Appointments|Event|false|false||appointmentnull|Allergy and Immunology|Title|false|false||Allergy and Immunologynull|Allergy - Charge Type Reason|Finding|false|false||Allergy
null|Allergic disposition|Finding|false|false||Allergy
null|Hypersensitivity|Finding|false|false||Allergy
null|Response to antigens|Finding|false|false||Allergy
null|History of allergies|Finding|false|false||Allergy
null|Allergic Reaction|Finding|false|false||Allergynull|Allergy Specialty|Title|false|false||Allergynull|Diagnostic Service Section ID - Immunology|Finding|false|false||Immunologynull|Immunology|Title|false|false||Immunologynull|immunology aspects|Modifier|false|false||Immunologynull|Medications on admission|Finding|false|false||Medications on Admissionnull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|On admission|Time|false|false||on Admissionnull|Admission activity|Procedure|false|false||Admission
null|Hospital admission|Procedure|false|false||Admissionnull|albuterol sulfate|Drug|false|false||Albuterol sulfate
null|albuterol sulfate|Drug|false|false||Albuterol sulfatenull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfate
null|Sulfates, Inorganic|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|sulfate ion|Drug|false|false||sulfate
null|Sulfates, Unspecified or Sulfate Ion|Drug|false|false||sulfatenull|NEB protein, human|Drug|false|false||Neb
null|NEB protein, human|Drug|false|false||Neb
null|Nebulizer solution|Drug|false|false||Nebnull|NEB gene|Finding|false|false||Neb
null|mitotic nuclear membrane disassembly|Finding|false|false||Nebnull|three times a day at institution-specified times|Time|false|false||TID
null|Three times daily|Time|false|false||TIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|albuterol|Drug|false|false||Albuterol
null|albuterol|Drug|false|false||Albuterolnull|ProAir|Drug|false|false||ProAir HFA
null|ProAir|Drug|false|false||ProAir HFAnull|ProAir|Drug|false|false||ProAir
null|ProAir|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAir
null|Pro-Air Procaterol|Drug|false|false||ProAirnull|Facial Hemiatrophy|Disorder|false|false||HFAnull|High frequency audiometry|Procedure|false|false||HFAnull|microgram|LabModifier|false|false||mcgnull|Inhalant dose form|Drug|false|false||INH
null|isoniazid|Drug|false|false||INH
null|isoniazid|Drug|false|false||INHnull|Inhalation Route of Administration|Finding|false|false||INHnull|Ingush language|Entity|false|false||INHnull|Inhalation Dosing Unit|LabModifier|false|false||INHnull|Puff Dosing Unit|LabModifier|false|false||puff
null|Picofarad|LabModifier|false|false||puffnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|cephalexin|Drug|false|false||Cephalexin
null|cephalexin|Drug|false|false||Cephalexinnull|Adderall-XR|Drug|false|false||Adderall XR
null|Adderall-XR|Drug|false|false||Adderall XRnull|Adderall|Drug|false|false||Adderall
null|Adderall|Drug|false|false||Adderallnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|ergocalciferol|Drug|false|false||Ergocalciferol (vitamin D2)
null|ergocalciferol|Drug|false|false||Ergocalciferol (vitamin D2)
null|ergocalciferol|Drug|false|false||Ergocalciferol (vitamin D2)null|Ergocalciferol Drug Product|Drug|false|false||Ergocalciferol
null|Ergocalciferol Drug Product|Drug|false|false||Ergocalciferol
null|ergocalciferol|Drug|false|false||Ergocalciferol
null|ergocalciferol|Drug|false|false||Ergocalciferol
null|ergocalciferol|Drug|false|false||Ergocalciferolnull|ergocalciferol|Drug|false|false||vitamin D2
null|ergocalciferol|Drug|false|false||vitamin D2
null|ergocalciferol|Drug|false|false||vitamin D2null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitamin
null|Vitamins|Drug|false|false||vitaminnull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Nexium|Drug|false|false||Nexium
null|Nexium|Drug|false|false||Nexiumnull|Every morning|Time|false|false||QAMnull|Vivelle|Drug|false|false||Vivelle
null|Vivelle|Drug|false|false||Vivelle
null|Vivelle|Drug|false|false||Vivellenull|Patch - Extended Release Film|Drug|false|false||Patch
null|Human patch material|Drug|false|false||Patch
null|Body tissue patch material|Drug|false|false||Patchnull|Plaque (lesion)|Finding|false|false||Patchnull|Patch Dosage Form|Device|false|false||Patch
null|Surgical patch|Device|false|false||Patchnull|Patch (unit of presentation)|LabModifier|false|false||Patch
null|Patch Dosing Unit|LabModifier|false|false||Patchnull|Weekly|Time|false|false||/ weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|Diflucan|Drug|false|false||Diflucan
null|Diflucan|Drug|false|false||Diflucannull|hydroxyzine hydrochloride|Drug|false|false||Hydroxyzine HCl
null|hydroxyzine hydrochloride|Drug|false|false||Hydroxyzine HClnull|hydroxyzine|Drug|false|false||Hydroxyzine
null|hydroxyzine|Drug|false|false||Hydroxyzinenull|Flinders medical centre-7 marker|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HCl
null|hydrochloride|Drug|false|false||HClnull|Hairy Cell Leukemia|Disorder|false|false||HClnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|ibuprofen|Drug|false|false||Ibuprofen
null|ibuprofen|Drug|false|false||Ibuprofennull|Every eight hours|Time|false|false||Q8Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Linzess|Drug|false|false||Linzess
null|Linzess|Drug|false|false||Linzessnull|microgram|LabModifier|false|false||mcgnull|Ativan|Drug|false|false||Ativan
null|Ativan|Drug|false|false||Ativannull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|metolazone|Drug|false|false||Metolazone
null|metolazone|Drug|false|false||Metolazonenull|Zofran|Drug|false|false||Zofran
null|Zofran|Drug|false|false||Zofrannull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|oxycodone|Drug|false|false||Oxycodone
null|oxycodone|Drug|false|false||Oxycodonenull|Oxycodone measurement|Procedure|false|false||Oxycodonenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|potassium chloride|Drug|false|false||Potassium chloride
null|potassium chloride|Drug|false|false||Potassium chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||chloride
null|Chlorides|Drug|false|false||chloridenull|Chloride metabolic function|Finding|false|false||chloridenull|Chloride measurement|Procedure|false|false||chloridenull|Oral Liquid Product|Drug|false|false|C0226896|Oral Liquidnull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1304698;C1272919;C1273619;C1527415;C4521986;C0301571|Oralnull|Oral|Modifier|false|false||Oralnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false|C0226896|Liquidnull|Liquid diet|Procedure|false|false|C0226896|Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|30mL|LabModifier|false|false||30mlnull|Four times daily|Time|false|false||QIDnull|propranolol|Drug|false|false||Propranolol
null|propranolol|Drug|false|false||Propranololnull|Once a day, at bedtime|Time|false|false||QHSnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Ambien|Drug|false|false||Ambien
null|Ambien|Drug|false|false||Ambiennull|Once a day, at bedtime|Time|false|false||QHSnull|null|Finding|false|false||catheternull|catheter device|Device|false|false||catheter
null|XXX>Catheter|Device|false|false||catheternull|docusate sodium|Drug|false|false||Docusate sodium
null|docusate sodium|Drug|false|false||Docusate sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|Lactobacillus|Entity|false|false||LACTOBACILLUSnull|combination - answer to question|Finding|false|false||COMBINATIONnull|combination of objects|Entity|false|false||COMBINATIONnull|Combined|Modifier|false|false||COMBINATIONnull|Medication.discharge|Finding|false|false||Discharge Medicationsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Pharmaceutical Preparations|Drug|false|false||Medicationsnull|Medications|Finding|false|false||Medicationsnull|null|Attribute|false|false||Medications
null|null|Attribute|false|false||Medicationsnull|docusate sodium|Drug|false|false||Docusate Sodium
null|docusate sodium|Drug|false|false||Docusate Sodiumnull|docusate|Drug|false|false||Docusate
null|docusate|Drug|false|false||Docusatenull|Sodium supplements|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|sodium|Drug|false|false||Sodium
null|Sodium Drug Class|Drug|false|false||Sodiumnull|Sodium metabolic function|Finding|false|false||Sodiumnull|Sodium measurement|Procedure|false|false||Sodiumnull|Liquid Dosage Form|Drug|false|false||Liquid
null|Liquid substance|Drug|false|false||Liquidnull|Liquid (finding)|Finding|false|false||Liquidnull|Liquid diet|Procedure|false|false||Liquidnull|Liquid (state of matter)|Modifier|false|false||Liquidnull|BID protein, human|Drug|false|false||BID
null|BID protein, human|Drug|false|false||BIDnull|Body integrity dysphoria|Disorder|false|false||BIDnull|BID gene|Finding|false|false||BIDnull|Twice a day|Time|false|false||BIDnull|docusate sodium|Drug|false|false||docusate sodium
null|docusate sodium|Drug|false|false||docusate sodiumnull|docusate|Drug|false|false||docusate
null|docusate|Drug|false|false||docusatenull|Sodium supplements|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|sodium|Drug|false|false||sodium
null|Sodium Drug Class|Drug|false|false||sodiumnull|Sodium metabolic function|Finding|false|false||sodiumnull|Sodium measurement|Procedure|false|false||sodiumnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1561538;C1561539;C1527415|mouth
null|Oral region|Anatomy|false|false|C1561538;C1561539;C1527415|mouthnull|Twice a day|Time|false|false||twice a daynull|Transaction counts and value totals - day|Finding|false|false|C0230028;C0226896|day
null|Precision - day|Finding|false|false|C0230028;C0226896|daynull|Land Dayak Languages|Entity|false|false||daynull|day|Time|false|false||day
null|Daily|Time|false|false||daynull|PRSS30P gene|Finding|false|false||Dispnull|Dispense (activity)|Event|false|false||Dispnull|capsule (pharmacologic)|Drug|false|false|C0524463;C1325531|Capsulenull|Microbial anatomical capsule structure|Anatomy|false|false|C0006935|Capsule
null|Structure of organ capsule|Anatomy|false|false|C0006935|Capsulenull|Capsule Shape|Modifier|false|false||Capsulenull|Capsule (unit of presentation)|LabModifier|false|false||Capsule
null|Capsule Dosing Unit|LabModifier|false|false||Capsulenull|refill|Finding|false|false||Refillsnull|bisacodyl|Drug|false|false||Bisacodyl
null|bisacodyl|Drug|false|false||Bisacodylnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Constipation|Finding|false|false||Constipationnull|bisacodyl|Drug|false|false||bisacodyl
null|bisacodyl|Drug|false|false||bisacodylnull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Release - action (qualifier value)|Finding|false|false||release
null|Released (action)|Finding|false|false||releasenull|Discharge (release)|Procedure|false|false||release
null|Release (procedure)|Procedure|false|false||release
null|Patient Discharge|Procedure|false|false||releasenull|Oral cavity|Anatomy|false|false|C0009806|mouth
null|Oral region|Anatomy|false|false|C0009806|mouthnull|Constipation|Finding|false|false|C0230028;C0226896|constipationnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|metolazone|Drug|false|false||Metolazone
null|metolazone|Drug|false|false||Metolazonenull|Daily|Time|false|false||DAILYnull|Nexium|Drug|false|false||NexIUM
null|Nexium|Drug|false|false||NexIUMnull|esomeprazole magnesium|Drug|false|false||esomeprazole magnesium
null|esomeprazole magnesium|Drug|false|false||esomeprazole magnesiumnull|esomeprazole|Drug|false|false||esomeprazole
null|esomeprazole|Drug|false|false||esomeprazolenull|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||magnesium
null|magnesium|Drug|false|false||magnesium
null|magnesium|Drug|false|false||magnesium
null|Magnesium Drug Class|Drug|false|false||magnesium
null|Magnesium supplements, alimentary tract and metabolism|Drug|false|false||magnesiumnull|Magnesium measurement|Procedure|false|false||magnesiumnull|Oral Dosage Form|Drug|false|false|C0226896|Oralnull|Oral Route of Administration|Finding|false|false|C0226896|Oral
null|Oral (intended site)|Finding|false|false|C0226896|Oralnull|Oral cavity|Anatomy|false|false|C1272919;C1527415;C4521986|Oralnull|Oral|Modifier|false|false||Oralnull|Once - dosing instruction fragment|Finding|false|false||oncenull|Once (schedule frequency)|Time|false|false||oncenull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|Unit dose|LabModifier|false|false||Dose
null|Dosage|LabModifier|false|false||Dosenull|oxycodone|Drug|false|false||OxycoDONE
null|oxycodone|Drug|false|false||OxycoDONEnull|Oxycodone measurement|Procedure|false|false||OxycoDONEnull|Immediate Release Dosage Form|Drug|false|false||Immediate Releasenull|Query Priority - Immediate|Finding|false|false||Immediate
null|immediate - ResponseCode|Finding|false|false||Immediatenull|Immediate|Time|false|false||Immediate
null|Stat (do immediately)|Time|false|false||Immediatenull|Release - action (qualifier value)|Finding|false|false||Release
null|Released (action)|Finding|false|false||Releasenull|Discharge (release)|Procedure|false|false||Release
null|Release (procedure)|Procedure|false|false||Release
null|Patient Discharge|Procedure|false|false||Releasenull|Every six hours|Time|false|false||Q6Hnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Administration Method - Pain|Finding|false|false||pain
null|Pain|Finding|false|false||painnull|null|Attribute|false|false||painnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|oxycodone|Drug|false|false||oxycodone
null|oxycodone|Drug|false|false||oxycodonenull|Oxycodone measurement|Procedure|false|false||oxycodonenull|Tablet Dosage Form|Drug|false|false||tabletnull|Tablet (unit of presentation)|LabModifier|false|false||tablet
null|Tablet Dosing Unit|LabModifier|false|false||tabletnull|Oral Route of Administration|Finding|false|false|C0230028;C0226896|by mouthnull|Oral cavity|Anatomy|false|false|C1527415;C1415473;C1419996;C1708271;C5780798;C5575450;C1366514;C0751781|mouth
null|Oral region|Anatomy|false|false|C1527415;C1415473;C1419996;C1708271;C5780798;C5575450;C1366514;C0751781|mouthnull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false|C0230028;C0226896|hrsnull|HARS1 wt Allele|Finding|false|false|C0230028;C0226896|hrs
null|HARS1 gene|Finding|false|false|C0230028;C0226896|hrs
null|HGS wt Allele|Finding|false|false|C0230028;C0226896|hrs
null|HGS gene|Finding|false|false|C0230028;C0226896|hrs
null|ATN1 wt Allele|Finding|false|false|C0230028;C0226896|hrs
null|SRSF5 gene|Finding|false|false|C0230028;C0226896|hrsnull|Hour|Time|false|false||hrsnull|Tablet Dosage Form|Drug|false|false||Tabletnull|Tablet (unit of presentation)|LabModifier|false|false||Tablet
null|Tablet Dosing Unit|LabModifier|false|false||Tabletnull|refill|Finding|false|false||Refillsnull|propranolol|Drug|false|false||Propranolol
null|propranolol|Drug|false|false||Propranololnull|Daily|Time|false|false||DAILYnull|spironolactone|Drug|false|false||Spironolactone
null|spironolactone|Drug|false|false||Spironolactonenull|Daily|Time|false|false||DAILYnull|zolpidem tartrate|Drug|false|false||Zolpidem Tartrate
null|zolpidem tartrate|Drug|false|false||Zolpidem Tartratenull|zolpidem|Drug|false|false||Zolpidem
null|zolpidem|Drug|false|false||Zolpidemnull|tartrate|Drug|false|false||Tartrate
null|Tartrates|Drug|false|false||Tartrate
null|tartrate|Drug|false|false||Tartratenull|trimethoprim|Drug|false|false||Trimethoprim
null|trimethoprim|Drug|false|false||Trimethoprimnull|Daily|Time|false|false||DAILYnull|Vivelle|Drug|false|false||Vivelle
null|Vivelle|Drug|false|false||Vivelle
null|Vivelle|Drug|false|false||Vivellenull|estradiol|Drug|false|false||estradiol
null|estradiol|Drug|false|false||estradiol
null|estradiol|Drug|false|false||estradiolnull|Estradiol measurement|Procedure|false|false||estradiolnull|Transdermal Route of Administration|Finding|false|false||Transdermal
null|transdermal|Finding|false|false||Transdermal
null|Transdermal (intended site)|Finding|false|false||Transdermalnull|Weekly|Time|false|false||/weeknull|Transaction counts and value totals - week|Finding|false|false||weeknull|week|Time|false|false||weeknull|lorazepam|Drug|false|false||Lorazepam
null|lorazepam|Drug|false|false||Lorazepamnull|Daily|Time|false|false||DAILYnull|CIAO3 gene|Finding|false|false||PRNnull|As required|Time|false|false||PRN
null|Pro Re Nata|Time|false|false||PRNnull|Anxiety Disorders|Disorder|false|false||anxiety
null|Anxiety|Disorder|false|false||anxietynull|Anxiety symptoms|Finding|false|false||anxietynull|potassium chloride|Drug|false|false||Potassium Chloride
null|potassium chloride|Drug|false|false||Potassium Chloridenull|Potassium Drug Class|Drug|false|false||Potassium
null|Dietary Potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|potassium|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassium
null|Potassium supplement|Drug|false|false||Potassiumnull|Potassium metabolic function|Finding|false|false||Potassiumnull|Potassium measurement|Procedure|false|false||Potassiumnull|chloride ion|Drug|false|false||Chloride
null|Chlorides|Drug|false|false||Chloridenull|Chloride metabolic function|Finding|false|false||Chloridenull|Chloride measurement|Procedure|false|false||Chloridenull|mEq|LabModifier|false|false||mEqnull|Daily|Time|false|false||DAILYnull|Duration brand of oxymetazoline|Drug|false|false||Durationnull|Duration (temporal concept)|Time|false|false||Durationnull|24 Hours|Time|false|false||24 Hoursnull|Hour|Time|false|false||Hoursnull|Hold - dosing instruction fragment|Finding|false|false||Hold
null|hold - Data Operation|Finding|false|false||Holdnull|Hold (action)|Event|false|false||Holdnull|Discharge disposition|Finding|false|false||Discharge Dispositionnull|null|Attribute|false|false||Discharge Dispositionnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Patient disposition|Procedure|false|false||Dispositionnull|null|Attribute|false|false||Dispositionnull|Disposition|Modifier|false|false||Dispositionnull|Visit User Code - Home|Finding|false|false||Home
null|Address type - Home|Finding|false|false||Homenull|home health encounter|Procedure|false|false||Homenull|Organization unit type - Home|Entity|false|false||Homenull|Person location type - Home|Modifier|false|false||Home
null|Home environment|Modifier|false|false||Homenull|discharge diagnosis|Finding|false|false||Discharge Diagnosisnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Diagnosis Classification - Diagnosis|Finding|false|false||Diagnosis
null|diagnosis aspects|Finding|false|false||Diagnosisnull|Diagnosis|Procedure|false|false||Diagnosisnull|null|Attribute|false|false||Diagnosisnull|Urinary Retention|Finding|false|false|C0042027|urinary retentionnull|Bladder retention of urine|Attribute|false|false|C0042027|urinary retentionnull|Urinary tract|Anatomy|false|false|C0080274;C0333117;C0080274;C1753315;C0035280;C5700171|urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false|C0042027|retention
null|Retention (Psychology)|Finding|false|false|C0042027|retention
null|Retention of content|Finding|false|false|C0042027|retention
null|cellular entity retention|Finding|false|false|C0042027|retentionnull|Retention - dental|Attribute|false|false||retentionnull|Rectocele|Disorder|false|false||rectocelenull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Disease|Disorder|false|false||Conditionnull|Logical Condition|Finding|false|false||Conditionnull|null|Attribute|false|false||Conditionnull|Condition|Modifier|false|false||Conditionnull|Mental state|Finding|false|false||Mental Statusnull|null|Attribute|false|false||Mental Status
null|null|Attribute|false|false||Mental Statusnull|Psyche structure|Finding|false|false||Mentalnull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Remote control command - Clear|Finding|false|false||Clearnull|Clear|Modifier|false|false||Clear
null|Transparent (qualitative concept)|Modifier|false|false||Clearnull|Coherent|Finding|false|false||coherentnull|Level of consciousness|Finding|false|false||Level of Consciousnessnull|null|Attribute|false|false||Level of Consciousnessnull|Consciousness related finding|Finding|false|false||Consciousness
null|Conscious|Finding|false|false||Consciousness
null|null|Finding|false|false||Consciousnessnull|Alert brand of caffeine|Drug|false|false||Alert
null|Alert brand of caffeine|Drug|false|false||Alertnull|Mentally alert|Finding|false|false||Alert
null|Consciousness clear|Finding|false|false||Alert
null|Alert note|Finding|false|false||Alert
null|Alert|Finding|false|false||Alertnull|null|Attribute|false|false||Alertnull|Interaction|Finding|false|false||interactivenull|Activity Status|Modifier|false|false||Activity Statusnull|Activity (animal life circumstance)|Finding|false|false||Activity
null|Physical activity|Finding|false|false||Activitynull|Activities|Event|false|false||Activitynull|null|Modifier|false|false||Activitynull|What subject filter - Status|Finding|false|false||Statusnull|null|Attribute|false|false||Statusnull|Social status|Modifier|false|false||Status
null|Status|Modifier|false|false||Statusnull|Referral category - Ambulatory|Finding|false|false||Ambulatory
null|Ambulatory (qualifier value)|Finding|false|false||Ambulatory
null|Ambulatory|Finding|false|false||Ambulatory
null|Level of Care - Ambulatory|Finding|false|false||Ambulatorynull|ambulatory encounter|Procedure|false|false||Ambulatorynull|Specialty Type - Ambulatory|Title|false|false||Ambulatorynull|Coordination of Benefits - Independent|Finding|false|false||Independent
null|Religious Affiliation - Independent|Finding|false|false||Independent
null|Independence|Finding|false|false||Independent
null|Independently able|Finding|false|false||Independentnull|Discharge instructions|Finding|false|false||Discharge Instructionsnull|hospital discharge instructions (treatment)|Procedure|false|false||Discharge Instructionsnull|null|Attribute|false|false||Discharge Instructionsnull|Body Substance Discharge|Finding|false|false||Discharge
null|Discharge Body Fluid|Finding|false|false||Discharge
null|Body Fluid Discharge|Finding|false|false||Discharge
null|null|Finding|false|false||Dischargenull|Patient Discharge|Procedure|false|false||Dischargenull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructionsnull|FBXW7-AS1 gene|Finding|false|false||Dearnull|Gynecology service|Entity|false|false||Gynecology servicenull|Gynecology|Title|false|false||Gynecologynull|ActInformationPrivacyReason - service|Finding|false|false||servicenull|Software Service|Device|false|false||servicenull|Services|Event|false|false||servicenull|Stage level 2|Finding|false|false||Stage 2null|Tumor stage|Attribute|false|false||Stagenull|Stage|Time|false|false||Stage
null|Phase|Time|false|false||Stagenull|null|Procedure|false|false||placement
null|Implantation procedure|Procedure|false|false||placement
null|Clinical act of insertion|Procedure|false|false||placementnull|Placement|Modifier|false|false||placementnull|Posterior repair of vagina|Procedure|false|false||posterior colporrhaphy
null|Repair of rectocele|Procedure|false|false||posterior colporrhaphynull|Posterior pituitary disease|Disorder|false|false||posteriornull|Dorsal|Modifier|false|false||posteriornull|Suture of vagina|Procedure|false|false||colporrhaphynull|Graft Dosage Form|Drug|false|false|C0332835|graft
null|Graft material|Drug|false|false|C0332835|graftnull|Graft - Specimen Source Codes|Finding|false|false|C0332835|graftnull|Graft Procedures on the Head|Procedure|false|false|C0332835|graft
null|Grafting procedure|Procedure|false|false|C0332835|graftnull|Transplanted tissue|Anatomy|false|false|C0205792;C0080274;C0149771;C0181074;C1705210;C1546653;C1961139;C3683798|graftnull|Urinary Retention|Finding|false|false|C0042027;C0332835|urinary retentionnull|Bladder retention of urine|Attribute|false|false|C0042027|urinary retentionnull|Urinary tract|Anatomy|false|false|C0080274;C5700171|urinarynull|urinary|Modifier|false|false||urinarynull|Urinary Retention|Finding|false|false||retention
null|Retention (Psychology)|Finding|false|false||retention
null|Retention of content|Finding|false|false||retention
null|cellular entity retention|Finding|false|false||retentionnull|Retention - dental|Attribute|false|false||retentionnull|Rectocele|Disorder|false|false|C0332835|rectocelenull|Enterocele|Disorder|false|false|C0332835|enterocelenull|Procedure (set of actions)|Finding|false|false||procedurenull|Interventional procedure|Procedure|false|false||procedurenull|null|Attribute|false|false||procedurenull|Act Class - procedure|Event|false|false||procedurenull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Computer Operation|Procedure|false|false||operation
null|Operative Surgical Procedures|Procedure|false|false||operationnull|Operation Activity|Event|false|false||operationnull|severe allergic reaction|Finding|false|false||severe allergic reactionnull|Severe - Severity of Illness Code|Finding|false|false||severe
null|Intensity and Distress 5|Finding|false|false||severe
null|Severe - Triage Code|Finding|false|false||severe
null|Severe (severity modifier)|Finding|false|false||severe
null|Allergy Severity - Severe|Finding|false|false||severenull|Allergic Reaction|Finding|false|false||allergic reaction
null|Hypersensitivity|Finding|false|false||allergic reactionnull|Allergic|Finding|false|false||allergicnull|Reaction|Finding|false|false||reactionnull|Inventory of Callous-Unemotional Traits|Finding|false|false|C0228479|ICUnull|Structure of intraculminate fissure|Anatomy|false|false|C4554035|ICUnull|intensive care unit|Device|false|false||ICUnull|intensive care unit|Entity|false|false||ICUnull|Preventive monitoring|Procedure|false|false||monitoringnull|null|Event|false|false||monitoringnull|Then - dosing instruction fragment|Finding|false|false||thennull|Then|Time|false|false||thennull|Well (answer to question)|Finding|false|false||wellnull|Well (container)|Device|false|false||wellnull|Microplate Well|Modifier|false|false||well
null|Good|Modifier|false|false||well
null|Healthy|Modifier|false|false||wellnull|Patient Condition Code - Stable|Finding|false|false||stablenull|Stable status|Modifier|false|false||stablenull|Disease|Disorder|false|false||conditionnull|Logical Condition|Finding|false|false||conditionnull|null|Attribute|false|false||conditionnull|Condition|Modifier|false|false||conditionnull|Body Substance Discharge|Finding|false|false||discharge
null|Discharge Body Fluid|Finding|false|false||discharge
null|Body Fluid Discharge|Finding|false|false||discharge
null|null|Finding|false|false||dischargenull|Patient Discharge|Procedure|false|false||dischargenull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|Appointments|Event|false|false||appointmentsnull|Instructions|Finding|false|false||instructions
null|Instruction [Publication Type]|Finding|false|false||instructionsnull|null|Attribute|false|false||instructionsnull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener brand of docusate sodium|Drug|false|false||stool softener
null|Stool Softener|Drug|false|false||stool softenernull|Feces|Finding|false|false||stoolnull|Stool seat|Device|false|false||stoolnull|Colace|Drug|false|false||colace
null|Colace|Drug|false|false||colacenull|Narcotics|Drug|false|false||narcotics
null|Narcotics|Drug|false|false||narcoticsnull|Constipation|Finding|false|false||constipationnull|Narcotics|Drug|false|false||narcotic
null|Narcotics|Drug|false|false||narcoticnull|Sedatives|Drug|false|false||sedativenull|Pharmaceutical Preparations|Drug|false|false||medicationsnull|Medications|Finding|false|false||medicationsnull|null|Attribute|false|false||medications
null|null|Attribute|false|false||medicationsnull|Alcohols|Drug|false|false||alcohol
null|Alcohols|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcohol
null|ethanol|Drug|false|false||alcoholnull|Alcohol - Recreational Drug Use Code|Finding|false|false||alcoholnull|Greater Than|LabModifier|false|false||more thannull|More|LabModifier|false|false||morenull|Acetaminophen [EPC]|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophen
null|acetaminophen|Drug|false|false||acetaminophennull|Acetaminophen measurement|Procedure|false|false||acetaminophennull|acetaminophen|Drug|false|false||APAP
null|acetaminophen|Drug|false|false||APAPnull|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED|Disorder|false|false||APAPnull|HGS protein, human|Drug|false|false||hrs
null|HGS protein, human|Drug|false|false||hrsnull|Dentatorubral-Pallidoluysian Atrophy|Disorder|false|false||hrsnull|HARS1 wt Allele|Finding|false|false||hrs
null|HARS1 gene|Finding|false|false||hrs
null|HGS wt Allele|Finding|false|false||hrs
null|HGS gene|Finding|false|false||hrs
null|ATN1 wt Allele|Finding|false|false||hrs
null|SRSF5 gene|Finding|false|false||hrsnull|Hour|Time|false|false||hrsnull|Strenuous Exercise|Finding|false|false||strenuous activitynull|Strenuous|Modifier|false|false||strenuousnull|Activity (animal life circumstance)|Finding|false|false||activity
null|Physical activity|Finding|false|false||activitynull|Activities|Event|false|false||activitynull|null|Modifier|false|false||activitynull|Appointments|Event|false|false||appointmentnull|Carcinoma in situ of vagina|Disorder|false|false|C0042232;C1519910;C4482396|vagina
null|Benign neoplasm vagina|Disorder|false|false|C0042232;C1519910;C4482396|vagina
null|Vaginal Diseases|Disorder|false|false|C0042232;C1519910;C4482396|vaginanull|Procedure on vagina|Procedure|false|false|C0042232;C1519910;C4482396|vaginanull|Pelvis>Vagina|Anatomy|false|false|C0869896;C0154002;C0686277;C0042251|vagina
null|Mouse Vagina|Anatomy|false|false|C0869896;C0154002;C0686277;C0042251|vagina
null|Vagina|Anatomy|false|false|C0869896;C0154002;C0686277;C0042251|vaginanull|Tampons|Device|true|false||tamponsnull|Douching procedure|Procedure|true|false||douchingnull|Sex Behavior|Finding|true|false||sex
null|PLXNA3 gene|Finding|true|false||sex
null|Coitus|Finding|true|false||sex
null|null|Finding|true|false||sexnull|null|Attribute|true|false||sexnull|sex|Subject|false|false||sex
null|Gender|Subject|false|false||sexnull|week|Time|false|false||weeksnull|Heavy (weight) (qualifier value)|Modifier|false|false||heavy
null|Heavy (amount)|Modifier|false|false||heavynull|Lifting|Event|true|false||liftingnull|Physical object|Entity|false|false||objectsnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|null|Finding|false|false||regular dietnull|Regular|Modifier|false|false||regularnull|Diet (animal life circumstance)|Drug|false|false||diet
null|Diet|Drug|false|false||dietnull|diet - supply|Finding|false|false||dietnull|Diet therapy|Procedure|false|false||dietnull|Incision care|Procedure|false|false|C2338258|Incision carenull|Surgical wound|Disorder|false|false|C2338258|Incisionnull|Surgical incisions|Procedure|false|false|C2338258|Incisionnull|Cranial incision point|Anatomy|false|false|C0150258;C0332803;C0580931;C2362566;C1947933;C0184898|Incisionnull|In care (finding)|Finding|false|false|C2338258|care
null|Continuity Assessment Record and Evaluation|Finding|false|false|C2338258|carenull|care activity|Event|false|false|C2338258|carenull|Water Specimen|Drug|false|false||water
null|water|Drug|false|false||water
null|water|Drug|false|false||waternull|Water - Specimen Source Codes|Finding|false|false||waternull|Hydrotherapy|Procedure|false|false|C2338258|waternull|Does run (finding)|Finding|false|false||run
null|Running (physical activity)|Finding|false|false||run
null|Go Jogging or Running Question|Finding|false|false||run
null|Run action|Finding|false|false||runnull|Rundi language|Entity|false|false||runnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0020311;C0184898|incisionnull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Bathing|Procedure|false|false||bathnull|6 weeks|Time|false|false||6 weeksnull|week|Time|false|false||weeksnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|Fever symptoms (finding)|Finding|false|false||fever
null|Fever|Finding|false|false||fevernull|Severe - Severity of Illness Code|Finding|false|false|C0000726|severe
null|Intensity and Distress 5|Finding|false|false|C0000726|severe
null|Severe - Triage Code|Finding|false|false|C0000726|severe
null|Severe (severity modifier)|Finding|false|false|C0000726|severe
null|Allergy Severity - Severe|Finding|false|false|C0000726|severenull|Abdominal Pain|Finding|false|false|C0000726|abdominal painnull|Abdomen|Anatomy|false|false|C0000737;C1549543;C0030193;C5203119;C1547231;C0205082;C1547227;C1561581|abdominalnull|Abdominal (qualifier value)|Modifier|false|false||abdominalnull|Administration Method - Pain|Finding|false|false|C0000726|pain
null|Pain|Finding|false|false|C0000726|painnull|null|Attribute|false|false||painnull|Has difficulty doing (qualifier value)|Finding|false|false||difficultynull|Abnormal vaginal bleeding|Finding|false|false|C0042232|vaginal bleeding
null|Vaginal Hemorrhage|Finding|false|false|C0042232|vaginal bleedingnull|Vaginal Dosage Form|Drug|false|false|C0042232|vaginalnull|Vaginal Route of Administration|Finding|false|false|C0042232|vaginal
null|Vaginal (intended site)|Finding|false|false|C0042232|vaginalnull|Vagina|Anatomy|false|false|C3814046;C0332568;C1704436;C3540603;C1425478;C1425244;C0019080;C0578503;C2979982;C4521343;C1522570;C1272941|vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Hemorrhage|Finding|false|false|C0042232|bleedingnull|Pad Dosage Form|Drug|false|false|C3669270|padnull|Pad Mass|Disorder|false|false|C0042232;C3669270|pad
null|Peripheral Arterial Diseases|Disorder|false|false|C0042232;C3669270|padnull|PADI4 wt Allele|Finding|false|false|C3669270;C0042232|pad
null|PADI4 gene|Finding|false|false|C3669270;C0042232|pad
null|DHX40 gene|Finding|false|false|C3669270;C0042232|padnull|PAD Regimen|Procedure|false|false|C0042232;C3669270|padnull|Strucure of thick cushion of skin|Anatomy|false|false|C3540603;C1425478;C1425244;C0332568;C1704436;C3814046;C2347441|padnull|Pad Device|Device|false|false||pad
null|Pads|Device|false|false||padnull|Pad (unit of presentation)|LabModifier|false|false||pad
null|Pad Dosing Unit|LabModifier|false|false||padnull|Abnormal Vaginal Discharge|Finding|false|false|C0042232|abnormal vaginal dischargenull|Observation Interpretation - Abnormal|Finding|false|false||abnormal
null|Abnormal|Finding|false|false||abnormalnull|Vaginal discharge symptom|Finding|false|false|C0042232|vaginal discharge
null|Vaginal Discharge|Finding|false|false|C0042232|vaginal dischargenull|Vaginal Dosage Form|Drug|false|false|C0042232|vaginalnull|Vaginal Route of Administration|Finding|false|false|C0042232|vaginal
null|Vaginal (intended site)|Finding|false|false|C0042232|vaginalnull|Vagina|Anatomy|false|false|C1272941;C0030685;C0566986;C0600083;C1546601;C0012621;C2926602;C4521343;C1522570;C0227791;C0438692|vaginalnull|Vaginal|Modifier|false|false||vaginalnull|Body Substance Discharge|Finding|false|false|C0042232|discharge
null|Discharge Body Fluid|Finding|false|false|C0042232|discharge
null|Body Fluid Discharge|Finding|false|false|C0042232|discharge
null|null|Finding|false|false|C0042232|dischargenull|Patient Discharge|Procedure|false|false|C0042232|dischargenull|Erythema|Disorder|false|false||rednessnull|Redness|Finding|false|false||rednessnull|Red color|Modifier|false|false||rednessnull|Body Substance Discharge|Finding|false|false||drainage
null|Body Fluid Discharge|Finding|false|false||drainagenull|Drainage procedure|Procedure|false|false||drainagenull|Surgical wound|Disorder|false|false|C2338258|incisionnull|Surgical incisions|Procedure|false|false|C2338258|incisionnull|Cranial incision point|Anatomy|false|false|C0332803;C0184898|incisionnull|Nausea and vomiting|Finding|false|false||nausea/vomitingnull|Nausea|Finding|false|false||nauseanull|null|Attribute|false|false||nauseanull|Vomiting|Finding|false|false||vomitingnull|Unable|Finding|false|false||unablenull|Liquid substance|Drug|false|false||fluidsnull|Mouse Body Fluid or Substance|Finding|false|false||fluidsnull|Fluid Therapy|Procedure|false|false||fluidsnull|Food allergenic extracts|Drug|false|false||food
null|Food|Drug|false|false||food
null|Food allergenic extracts|Drug|false|false||foodnull|Pharmaceutical Preparations|Drug|false|false||medicationnull|medication - HL7 publishing domain|Finding|false|false||medication
null|Medications|Finding|false|false||medicationnull|HL7 Committee ID In RIM - Medical records|Finding|false|false||medical records
null|Medical Records|Finding|false|false||medical recordsnull|null|Attribute|false|false||medical recordsnull|Medical referral type|Finding|false|false||medical
null|Medical|Finding|false|false||medical
null|Medical school type|Finding|false|false||medicalnull|Medical service|Procedure|false|false||medicalnull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Quantity limited request - Records|Finding|false|false||records
null|Records|Finding|false|false||recordsnull|Query Quantity Unit - Records|Modifier|false|false||recordsnull|Hospitalization|Procedure|false|false||hospitalizationnull|Doctor - Title|Finding|false|false||doctornull|Physicians|Subject|false|false||doctornull|At home|Finding|false|false||at homenull|Visit User Code - Home|Finding|false|false||home
null|Address type - Home|Finding|false|false||homenull|home health encounter|Procedure|false|false||homenull|Organization unit type - Home|Entity|false|false||homenull|Person location type - Home|Modifier|false|false||home
null|Home environment|Modifier|false|false||homenull|follow-up|Procedure|false|false||Followupnull|Instructions|Finding|false|false||Instructions
null|Instruction [Publication Type]|Finding|false|false||Instructionsnull|null|Attribute|false|false||Instructions