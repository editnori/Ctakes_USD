 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|35,39
No|40,42
:|42,43
_|46,47
_|47,48
_|48,49
<EOL>|49,50
<EOL>|51,52
Admission|52,61
Date|62,66
:|66,67
_|69,70
_|70,71
_|71,72
Discharge|86,95
Date|96,100
:|100,101
_|104,105
_|105,106
_|106,107
<EOL>|107,108
<EOL>|109,110
Date|110,114
of|115,117
Birth|118,123
:|123,124
_|126,127
_|127,128
_|128,129
Sex|142,145
:|145,146
M|149,150
<EOL>|150,151
<EOL>|152,153
Service|153,160
:|160,161
MEDICINE|162,170
<EOL>|170,171
<EOL>|172,173
No|185,187
Allergies|188,197
/|197,198
ADRs|198,202
on|203,205
File|206,210
<EOL>|210,211
<EOL>|212,213
Attending|213,222
:|222,223
_|224,225
_|225,226
_|226,227
.|227,228
<EOL>|228,229
<EOL>|230,231
chest|248,253
pain|254,258
<EOL>|258,259
<EOL>|260,261
Major|261,266
Surgical|267,275
or|276,278
Invasive|279,287
Procedure|288,297
:|297,298
<EOL>|298,299
_|299,300
_|300,301
_|301,302
-|303,304
bedside|305,312
pericardiocentesis|313,331
at|332,334
_|335,336
_|336,337
_|337,338
<EOL>|338,339
<EOL>|339,340
<EOL>|341,342
HISTORY|371,378
OF|379,381
PRESENTING|382,392
ILLNESS|393,400
:|400,401
Mr.|402,405
_|406,407
_|407,408
_|408,409
is|410,412
a|413,414
_|415,416
_|416,417
_|417,418
<EOL>|418,419
male|419,423
with|424,428
rheumatoid|429,439
arthritis|440,449
,|449,450
DMARD|451,456
holiday|457,464
,|464,465
and|466,469
recent|470,476
,|476,477
brief|478,483
<EOL>|483,484
hospitalization|484,499
for|500,503
presumptive|504,515
pericarditis|516,528
,|528,529
returned|530,538
to|539,541
<EOL>|542,543
outside|543,550
<EOL>|550,551
hospital|551,559
with|560,564
probable|565,573
cardiac|574,581
tamponade|582,591
now|592,595
post-bedside|596,608
<EOL>|608,609
pericardiocentesis|609,627
with|628,632
drain|633,638
placement|639,648
prior|649,654
to|655,657
transfer|658,666
.|666,667
<EOL>|667,668
Importantly|668,679
,|679,680
patient|681,688
was|689,692
hospitalized|693,705
at|706,708
_|709,710
_|710,711
_|711,712
on|713,715
_|716,717
_|717,718
_|718,719
with|720,724
acute|725,730
pleuritic|731,740
chest|741,746
pain|747,751
of|752,754
two|755,758
-|758,759
day|759,762
duration|763,771
in|772,774
the|775,778
<EOL>|778,779
context|779,786
of|787,789
constellation|790,803
of|804,806
fatigue|807,814
,|814,815
malaise|816,823
,|823,824
upper|825,830
respiratory|831,842
<EOL>|842,843
symptoms|843,851
,|851,852
and|853,856
non-productive|857,871
cough|872,877
.|877,878
While|879,884
CTA|885,888
exonerated|889,899
<EOL>|899,900
pulmonary|900,909
embolism|910,918
,|918,919
thickened|920,929
pericardium|930,941
and|942,945
small|946,951
effusion|952,960
<EOL>|961,962
were|962,966
<EOL>|966,967
noted|967,972
,|972,973
suggesting|974,984
pericarditis|985,997
.|997,998
ECG|999,1002
revealed|1003,1011
subtle|1012,1018
diffuse|1019,1026
ST|1027,1029
<EOL>|1029,1030
elevations|1030,1040
in|1041,1043
keeping|1044,1051
with|1052,1056
pericarditis|1057,1069
.|1069,1070
Echocardiogram|1071,1085
<EOL>|1086,1087
confirmed|1087,1096
<EOL>|1096,1097
said|1097,1101
effusion|1102,1110
,|1110,1111
though|1112,1118
no|1119,1121
features|1122,1130
of|1131,1133
tamponade|1134,1143
were|1144,1148
appreciated|1149,1160
.|1160,1161
<EOL>|1161,1162
He|1162,1164
was|1165,1168
discharged|1169,1179
the|1180,1183
same|1184,1188
day|1189,1192
with|1193,1197
ibuprofen|1198,1207
600|1208,1211
mg|1212,1214
TID|1215,1218
and|1219,1222
<EOL>|1222,1223
colchicine|1223,1233
0.6|1234,1237
mg|1238,1240
BID|1241,1244
.|1244,1245
He|1246,1248
had|1249,1252
persistence|1253,1264
of|1265,1267
minor|1268,1273
residual|1274,1282
<EOL>|1283,1284
chest|1284,1289
<EOL>|1289,1290
pain|1290,1294
,|1294,1295
which|1296,1301
began|1302,1307
to|1308,1310
worsen|1311,1317
two|1318,1321
days|1322,1326
later|1327,1332
,|1332,1333
but|1334,1337
was|1338,1341
tolerable|1342,1351
<EOL>|1351,1352
until|1352,1357
yesterday|1358,1367
evening|1368,1375
when|1376,1380
it|1381,1383
evolved|1384,1391
to|1392,1394
severe|1395,1401
,|1401,1402
unrelenting|1403,1414
<EOL>|1414,1415
pain|1415,1419
across|1420,1426
his|1427,1430
precordium|1431,1441
likened|1442,1449
to|1450,1452
"|1453,1454
wearing|1454,1461
shoulder|1462,1470
pads|1471,1475
<EOL>|1475,1476
bearing|1476,1483
down|1484,1488
on|1489,1491
him|1492,1495
.|1495,1496
"|1496,1497
He|1498,1500
notes|1501,1506
a|1507,1508
new|1509,1512
concurrent|1513,1523
substernal|1524,1534
chest|1535,1540
<EOL>|1540,1541
pain|1541,1545
that|1546,1550
"|1551,1552
goes|1552,1556
straight|1557,1565
to|1566,1568
his|1569,1572
back|1573,1577
.|1577,1578
"|1578,1579
He|1580,1582
then|1583,1587
became|1588,1594
dyspneic|1595,1603
,|1603,1604
<EOL>|1604,1605
prompting|1605,1614
him|1615,1618
to|1619,1621
seek|1622,1626
care|1627,1631
.|1631,1632
He|1633,1635
arrived|1636,1643
at|1644,1646
_|1647,1648
_|1648,1649
_|1649,1650
hypotensive|1651,1662
<EOL>|1662,1663
with|1663,1667
SBP|1668,1671
in|1672,1674
the|1675,1678
80|1679,1681
-|1681,1682
range|1682,1687
.|1687,1688
He|1689,1691
was|1692,1695
borderline|1696,1706
tachycardic|1707,1718
and|1719,1722
in|1723,1725
<EOL>|1725,1726
mild|1726,1730
respiratory|1731,1742
distress|1743,1751
,|1751,1752
but|1753,1756
oxygenation|1757,1768
was|1769,1772
acceptable|1773,1783
.|1783,1784
He|1785,1787
<EOL>|1787,1788
rapidly|1788,1795
received|1796,1804
three|1805,1810
liters|1811,1817
of|1818,1820
fluid|1821,1826
for|1827,1830
presumptive|1831,1842
tamponade|1843,1852
<EOL>|1852,1853
within|1853,1859
the|1860,1863
confines|1864,1872
of|1873,1875
poor|1876,1880
windows|1881,1888
on|1889,1891
bedside|1892,1899
echocardiogram|1900,1914
.|1914,1915
<EOL>|1915,1916
Pericardiocentesis|1916,1934
yielded|1935,1942
400|1943,1946
cc|1947,1949
or|1950,1952
more|1953,1957
of|1958,1960
serous|1961,1967
fluid|1968,1973
and|1974,1977
a|1978,1979
<EOL>|1979,1980
pericardial|1980,1991
drain|1992,1997
was|1998,2001
placed|2002,2008
.|2008,2009
Hemodynamics|2010,2022
rapidly|2023,2030
improved|2031,2039
.|2039,2040
On|2041,2043
<EOL>|2043,2044
arrival|2044,2051
to|2052,2054
_|2055,2056
_|2056,2057
_|2057,2058
ED|2059,2061
,|2061,2062
patient|2063,2070
was|2071,2074
indeed|2075,2081
hemodynamically|2082,2097
stable|2098,2104
<EOL>|2104,2105
but|2105,2108
was|2109,2112
then|2113,2117
in|2118,2120
moderate|2121,2129
respiratory|2130,2141
distress|2142,2150
,|2150,2151
requiring|2152,2161
<EOL>|2161,2162
non-rebreather|2162,2176
.|2176,2177
He|2178,2180
was|2181,2184
given|2185,2190
Lasix|2191,2196
20|2197,2199
mg|2200,2202
IV.|2203,2206
Bedside|2207,2214
<EOL>|2214,2215
echocardiogram|2215,2229
was|2230,2233
limited|2234,2241
,|2241,2242
but|2243,2246
preliminarily|2247,2260
suggestive|2261,2271
of|2272,2274
<EOL>|2275,2276
small|2276,2281
<EOL>|2281,2282
residual|2282,2290
effusion|2291,2299
.|2299,2300
In|2301,2303
the|2304,2307
CCU|2308,2311
,|2311,2312
patient|2313,2320
notes|2321,2326
resurgence|2327,2337
of|2338,2340
said|2341,2345
<EOL>|2345,2346
chest|2346,2351
pain|2352,2356
.|2356,2357
His|2358,2361
dyspnea|2362,2369
is|2370,2372
improving|2373,2382
.|2382,2383
An|2384,2386
additional|2387,2397
250|2398,2401
cc|2402,2404
was|2405,2408
<EOL>|2408,2409
drained|2409,2416
.|2416,2417
<EOL>|2418,2419
<EOL>|2420,2421
<EOL>|2442,2443
Cardiac|2468,2475
-|2487,2488
Pericarditis|2488,2500
,|2500,2501
as|2502,2504
above|2505,2510
.|2510,2511
<EOL>|2511,2512
-|2512,2513
Hypertension|2513,2525
.|2525,2526
<EOL>|2526,2527
-|2527,2528
Dyslipidemia|2528,2540
.|2540,2541
<EOL>|2542,2543
<EOL>|2544,2545
Other|2546,2551
PMH|2552,2555
:|2555,2556
<EOL>|2558,2559
-|2559,2560
Rheumatoid|2560,2570
arthritis|2571,2580
.|2580,2581
<EOL>|2582,2583
-|2583,2584
Remote|2584,2590
traumatic|2591,2600
DVT|2601,2604
.|2604,2605
<EOL>|2605,2606
-|2606,2607
Cholecystectomy|2607,2622
.|2622,2623
<EOL>|2623,2624
-|2624,2625
Appendectomy|2625,2637
.|2637,2638
<EOL>|2638,2639
-|2639,2640
Tonsillectomy|2640,2653
.|2653,2654
<EOL>|2654,2655
-|2655,2656
Left|2656,2660
wrist|2661,2666
reconstruction|2667,2681
.|2681,2682
<EOL>|2682,2683
-|2683,2684
Right|2684,2689
rotator|2690,2697
cuff|2698,2702
reconstruction|2703,2717
.|2717,2718
<EOL>|2718,2719
<EOL>|2719,2720
<EOL>|2721,2722
:|2736,2737
<EOL>|2737,2738
_|2738,2739
_|2739,2740
_|2740,2741
<EOL>|2741,2742
:|2756,2757
<EOL>|2757,2758
paternal|2758,2766
history|2767,2774
of|2775,2777
ureothelial|2778,2789
carcinoma|2790,2799
.|2799,2800
<EOL>|2800,2801
Maternal|2801,2809
history|2810,2817
of|2818,2820
diabetes|2821,2829
.|2829,2830
<EOL>|2831,2832
<EOL>|2832,2833
<EOL>|2834,2835
ADMISSION|2850,2859
PHYSICAL|2860,2868
EXAMINATION|2869,2880
:|2880,2881
<EOL>|2883,2884
=|2884,2885
=|2885,2886
=|2886,2887
=|2887,2888
=|2888,2889
=|2889,2890
=|2890,2891
=|2891,2892
=|2892,2893
=|2893,2894
=|2894,2895
=|2895,2896
=|2896,2897
=|2897,2898
=|2898,2899
=|2899,2900
=|2900,2901
=|2901,2902
=|2902,2903
=|2903,2904
=|2904,2905
=|2905,2906
=|2906,2907
=|2907,2908
=|2908,2909
=|2909,2910
=|2910,2911
=|2911,2912
=|2912,2913
=|2913,2914
=|2914,2915
=|2915,2916
=|2916,2917
<EOL>|2917,2918
VS|2919,2921
:|2921,2922
T|2923,2924
96.7|2925,2929
,|2929,2930
HR|2931,2933
81|2934,2936
,|2936,2937
BP|2938,2940
136|2941,2944
/|2944,2945
81|2945,2947
,|2947,2948
O2|2949,2951
94|2952,2954
%|2954,2955
6L|2956,2958
<EOL>|2959,2960
GENERAL|2961,2968
:|2968,2969
obese|2970,2975
male|2976,2980
in|2981,2983
mild|2984,2988
to|2989,2991
moderate|2992,3000
respiratory|3001,3012
distress|3013,3021
.|3021,3022
<EOL>|3024,3025
HEENT|3026,3031
:|3031,3032
anicteric|3033,3042
sclerae|3043,3050
.|3050,3051
Oropharynx|3052,3062
clear|3063,3068
.|3068,3069
<EOL>|3071,3072
NECK|3073,3077
:|3077,3078
JVP|3079,3082
at|3083,3085
mandibular|3086,3096
angle|3097,3102
.|3102,3103
<EOL>|3104,3105
CARDIAC|3106,3113
:|3113,3114
tachycardic|3115,3126
,|3126,3127
regular|3128,3135
with|3136,3140
rare|3141,3145
ectopy|3146,3152
,|3152,3153
S1|3154,3156
/|3156,3157
S2|3157,3159
within|3160,3166
<EOL>|3167,3168
the|3168,3171
<EOL>|3171,3172
confines|3172,3180
of|3181,3183
body|3184,3188
habitus|3189,3196
.|3196,3197
Subtle|3198,3204
pericardial|3205,3216
rub|3217,3220
.|3220,3221
Pericardial|3222,3233
<EOL>|3233,3234
drain|3234,3239
with|3240,3244
serosanguinous|3245,3259
fluid|3260,3265
.|3265,3266
Sternal|3267,3274
tenderness|3275,3285
.|3285,3286
<EOL>|3287,3288
LUNGS|3289,3294
:|3294,3295
Conversational|3296,3310
dyspnea|3311,3318
but|3319,3322
tachypnea|3323,3332
is|3333,3335
slowing|3336,3343
.|3343,3344
Diffuse|3345,3352
<EOL>|3352,3353
wheezing|3353,3361
and|3362,3365
crackles|3366,3374
in|3375,3377
bilateral|3378,3387
lung|3388,3392
fields|3393,3399
.|3399,3400
<EOL>|3402,3403
ABDOMEN|3404,3411
:|3411,3412
obese|3413,3418
,|3418,3419
soft|3420,3424
,|3424,3425
non-tender|3426,3436
.|3436,3437
<EOL>|3437,3438
EXTREMITIES|3439,3450
:|3450,3451
Warm|3452,3456
,|3456,3457
well|3458,3462
perfused|3463,3471
,|3471,3472
2|3473,3474
+|3474,3475
pitting|3476,3483
edema|3484,3489
to|3490,3492
knees|3493,3498
.|3498,3499
<EOL>|3501,3502
SKIN|3503,3507
:|3507,3508
Chronic|3509,3516
bilateral|3517,3526
venous|3527,3533
stasis|3534,3540
dermatitis|3541,3551
.|3551,3552
<EOL>|3554,3555
PULSES|3556,3562
:|3562,3563
Distal|3564,3570
pulses|3571,3577
palpable|3578,3586
and|3587,3590
symmetric|3591,3600
.|3600,3601
<EOL>|3603,3604
NEURO|3605,3610
:|3610,3611
non-focal|3612,3621
.|3621,3622
<EOL>|3622,3623
<EOL>|3623,3624
DISCHARGE|3624,3633
PHYSICAL|3634,3642
EXAMINATION|3643,3654
:|3654,3655
<EOL>|3657,3658
=|3658,3659
=|3659,3660
=|3660,3661
=|3661,3662
=|3662,3663
=|3663,3664
=|3664,3665
=|3665,3666
=|3666,3667
=|3667,3668
=|3668,3669
=|3669,3670
=|3670,3671
=|3671,3672
=|3672,3673
=|3673,3674
=|3674,3675
=|3675,3676
=|3676,3677
=|3677,3678
=|3678,3679
=|3679,3680
=|3680,3681
=|3681,3682
=|3682,3683
=|3683,3684
=|3684,3685
=|3685,3686
=|3686,3687
=|3687,3688
=|3688,3689
=|3689,3690
=|3690,3691
<EOL>|3691,3692
GENERAL|3692,3699
:|3699,3700
obese|3701,3706
male|3707,3711
in|3712,3714
mild|3715,3719
to|3720,3722
moderate|3723,3731
respiratory|3732,3743
distress|3744,3752
.|3752,3753
<EOL>|3755,3756
HEENT|3757,3762
:|3762,3763
anicteric|3764,3773
sclerae|3774,3781
.|3781,3782
Oropharynx|3783,3793
clear|3794,3799
.|3799,3800
<EOL>|3802,3803
NECK|3804,3808
:|3808,3809
JVP|3810,3813
not|3814,3817
appreciated|3818,3829
.|3829,3830
<EOL>|3831,3832
CARDIAC|3833,3840
:|3840,3841
normal|3842,3848
rate|3849,3853
and|3854,3857
rhythm|3858,3864
,|3864,3865
S1|3866,3868
/|3868,3869
S2|3869,3871
within|3872,3878
the|3879,3882
confines|3883,3891
of|3892,3894
<EOL>|3894,3895
body|3895,3899
habitus|3900,3907
.|3907,3908
No|3909,3911
pericardial|3912,3923
rub|3924,3927
appreciated|3928,3939
.|3939,3940
<EOL>|3941,3942
LUNGS|3943,3948
:|3948,3949
Decreased|3950,3959
respiratory|3960,3971
effort|3972,3978
compared|3979,3987
to|3988,3990
yesterday|3991,4000
.|4000,4001
<EOL>|4001,4002
Expiratory|4002,4012
wheezing|4013,4021
and|4022,4025
bibasilar|4026,4035
crackles|4036,4044
.|4044,4045
<EOL>|4045,4046
ABDOMEN|4047,4054
:|4054,4055
obese|4056,4061
,|4061,4062
soft|4063,4067
,|4067,4068
non-tender|4069,4079
,|4079,4080
non-distended|4081,4094
.|4094,4095
<EOL>|4095,4096
EXTREMITIES|4097,4108
:|4108,4109
Warm|4110,4114
,|4114,4115
well|4116,4120
perfused|4121,4129
,|4129,4130
1|4131,4132
to|4133,4135
2|4136,4137
+|4137,4138
pitting|4139,4146
edema|4147,4152
to|4153,4155
<EOL>|4155,4156
knees|4156,4161
.|4161,4162
<EOL>|4164,4165
SKIN|4166,4170
:|4170,4171
Chronic|4172,4179
venous|4180,4186
stasis|4187,4193
dermatitis|4194,4204
.|4204,4205
<EOL>|4207,4208
PULSES|4209,4215
:|4215,4216
Distal|4217,4223
pulses|4224,4230
palpable|4231,4239
and|4240,4243
symmetric|4244,4253
.|4253,4254
<EOL>|4256,4257
NEURO|4258,4263
:|4263,4264
non-focal|4265,4274
.|4274,4275
<EOL>|4275,4276
<EOL>|4277,4278
Pertinent|4278,4287
Results|4288,4295
:|4295,4296
<EOL>|4296,4297
ADMISSION|4297,4306
LABS|4307,4311
:|4311,4312
<EOL>|4312,4313
=|4313,4314
=|4314,4315
=|4315,4316
=|4316,4317
=|4317,4318
=|4318,4319
=|4319,4320
=|4320,4321
=|4321,4322
=|4322,4323
=|4323,4324
=|4324,4325
=|4325,4326
=|4326,4327
=|4327,4328
<EOL>|4328,4329
_|4329,4330
_|4330,4331
_|4331,4332
10|4333,4335
:|4335,4336
57PM|4336,4340
WBC|4343,4346
-|4346,4347
16|4347,4349
.|4349,4350
9|4350,4351
*|4351,4352
RBC|4353,4356
-|4356,4357
4|4357,4358
.|4358,4359
63|4359,4361
HGB|4362,4365
-|4365,4366
14.2|4366,4370
HCT|4371,4374
-|4374,4375
43.1|4375,4379
MCV|4380,4383
-|4383,4384
93|4384,4386
<EOL>|4387,4388
MCH|4388,4391
-|4391,4392
30.7|4392,4396
MCHC|4397,4401
-|4401,4402
32.9|4402,4406
RDW|4407,4410
-|4410,4411
13.1|4411,4415
RDWSD|4416,4421
-|4421,4422
44.1|4422,4426
<EOL>|4426,4427
_|4427,4428
_|4428,4429
_|4429,4430
10|4431,4433
:|4433,4434
57PM|4434,4438
NEUTS|4441,4446
-|4446,4447
85|4447,4449
.|4449,4450
5|4450,4451
*|4451,4452
LYMPHS|4453,4459
-|4459,4460
4|4460,4461
.|4461,4462
3|4462,4463
*|4463,4464
MONOS|4465,4470
-|4470,4471
9.4|4471,4474
EOS|4475,4478
-|4478,4479
0|4479,4480
.|4480,4481
1|4481,4482
*|4482,4483
<EOL>|4484,4485
BASOS|4485,4490
-|4490,4491
0.2|4491,4494
IM|4495,4497
_|4498,4499
_|4499,4500
_|4500,4501
AbsNeut|4502,4509
-|4509,4510
14|4510,4512
.|4512,4513
43|4513,4515
*|4515,4516
AbsLymp|4517,4524
-|4524,4525
0|4525,4526
.|4526,4527
72|4527,4529
*|4529,4530
AbsMono|4531,4538
-|4538,4539
1|4539,4540
.|4540,4541
58|4541,4543
*|4543,4544
<EOL>|4545,4546
AbsEos|4546,4552
-|4552,4553
0|4553,4554
.|4554,4555
01|4555,4557
*|4557,4558
AbsBaso|4559,4566
-|4566,4567
0.04|4567,4571
<EOL>|4571,4572
_|4572,4573
_|4573,4574
_|4574,4575
10|4576,4578
:|4578,4579
57PM|4579,4583
_|4586,4587
_|4587,4588
_|4588,4589
PTT|4590,4593
-|4593,4594
27.2|4594,4598
_|4599,4600
_|4600,4601
_|4601,4602
<EOL>|4602,4603
_|4603,4604
_|4604,4605
_|4605,4606
10|4607,4609
:|4609,4610
57PM|4610,4614
GLUCOSE|4617,4624
-|4624,4625
269|4625,4628
*|4628,4629
UREA|4630,4634
N|4635,4636
-|4636,4637
20|4637,4639
CREAT|4640,4645
-|4645,4646
0.9|4646,4649
SODIUM|4650,4656
-|4656,4657
135|4657,4660
<EOL>|4661,4662
POTASSIUM|4662,4671
-|4671,4672
5.3|4672,4675
CHLORIDE|4676,4684
-|4684,4685
106|4685,4688
TOTAL|4689,4694
CO2|4695,4698
-|4698,4699
18|4699,4701
*|4701,4702
ANION|4703,4708
GAP|4709,4712
-|4712,4713
11|4713,4715
<EOL>|4715,4716
_|4716,4717
_|4717,4718
_|4718,4719
10|4720,4722
:|4722,4723
57PM|4723,4727
CALCIUM|4730,4737
-|4737,4738
7|4738,4739
.|4739,4740
4|4740,4741
*|4741,4742
PHOSPHATE|4743,4752
-|4752,4753
3.1|4753,4756
MAGNESIUM|4757,4766
-|4766,4767
1.6|4767,4770
<EOL>|4770,4771
_|4771,4772
_|4772,4773
_|4773,4774
10|4775,4777
:|4777,4778
57PM|4778,4782
cTropnT|4785,4792
-|4792,4793
<|4793,4794
0|4794,4795
.|4795,4796
01|4796,4798
<EOL>|4798,4799
_|4799,4800
_|4800,4801
_|4801,4802
11|4803,4805
:|4805,4806
03PM|4806,4810
LACTATE|4813,4820
-|4820,4821
2.0|4821,4824
<EOL>|4824,4825
_|4825,4826
_|4826,4827
_|4827,4828
01|4829,4831
:|4831,4832
05AM|4832,4836
PLEURAL|4837,4844
FLUID|4845,4850
STUDIES|4851,4858
_|4859,4860
_|4860,4861
_|4861,4862
<EOL>|4863,4864
Polys|4864,4869
-|4869,4870
94|4870,4872
*|4872,4873
Lymphs|4874,4880
-|4880,4881
2|4881,4882
*|4882,4883
Monos|4884,4889
-|4889,4890
4|4890,4891
*|4891,4892
<EOL>|4892,4893
<EOL>|4893,4894
IMAGING|4894,4901
:|4901,4902
<EOL>|4902,4903
=|4903,4904
=|4904,4905
=|4905,4906
=|4906,4907
=|4907,4908
=|4908,4909
=|4909,4910
=|4910,4911
<EOL>|4911,4912
_|4912,4913
_|4913,4914
_|4914,4915
TTE|4916,4919
<EOL>|4919,4920
The|4920,4923
left|4924,4928
atrium|4929,4935
is|4936,4938
normal|4939,4945
in|4946,4948
size|4949,4953
.|4953,4954
The|4955,4958
inferior|4959,4967
vena|4968,4972
cava|4973,4977
is|4978,4980
<EOL>|4981,4982
dilated|4982,4989
(|4990,4991
>|4991,4992
2.5|4992,4995
cm|4996,4998
)|4998,4999
.|4999,5000
There|5001,5006
is|5007,5009
normal|5010,5016
left|5017,5021
ventricular|5022,5033
<EOL>|5033,5034
wall|5034,5038
thickness|5039,5048
with|5049,5053
a|5054,5055
normal|5056,5062
cavity|5063,5069
size|5070,5074
.|5074,5075
There|5076,5081
is|5082,5084
suboptimal|5085,5095
<EOL>|5096,5097
image|5097,5102
quality|5103,5110
to|5111,5113
assess|5114,5120
regional|5121,5129
left|5130,5134
ventricular|5135,5146
<EOL>|5146,5147
function|5147,5155
.|5155,5156
Overall|5157,5164
left|5165,5169
ventricular|5170,5181
systolic|5182,5190
function|5191,5199
is|5200,5202
normal|5203,5209
.|5209,5210
<EOL>|5211,5212
Quantitative|5212,5224
biplane|5225,5232
left|5233,5237
ventricular|5238,5249
ejection|5250,5258
<EOL>|5258,5259
fraction|5259,5267
is|5268,5270
66|5271,5273
%|5274,5275
.|5275,5276
Left|5277,5281
ventricular|5282,5293
cardiac|5294,5301
index|5302,5307
is|5308,5310
normal|5311,5317
(|5318,5319
>|5319,5320
2.5|5320,5323
<EOL>|5324,5325
L|5325,5326
/|5326,5327
min|5327,5330
/|5330,5331
m2|5331,5333
)|5333,5334
.|5334,5335
No|5336,5338
ventricular|5339,5350
septal|5351,5357
defect|5358,5364
is|5365,5367
<EOL>|5367,5368
seen|5368,5372
.|5372,5373
Normal|5374,5380
right|5381,5386
ventricular|5387,5398
cavity|5399,5405
size|5406,5410
with|5411,5415
normal|5416,5422
free|5423,5427
wall|5428,5432
<EOL>|5433,5434
motion|5434,5440
.|5440,5441
There|5442,5447
is|5448,5450
abnormal|5451,5459
interventricular|5460,5476
<EOL>|5476,5477
septal|5477,5483
motion|5484,5490
.|5490,5491
The|5492,5495
aortic|5496,5502
sinus|5503,5508
diameter|5509,5517
is|5518,5520
normal|5521,5527
for|5528,5531
gender|5532,5538
<EOL>|5539,5540
with|5540,5544
normal|5545,5551
ascending|5552,5561
aorta|5562,5567
diameter|5568,5576
for|5577,5580
<EOL>|5580,5581
gender|5581,5587
.|5587,5588
The|5589,5592
aortic|5593,5599
arch|5600,5604
diameter|5605,5613
is|5614,5616
normal|5617,5623
.|5623,5624
There|5625,5630
is|5631,5633
no|5634,5636
evidence|5637,5645
<EOL>|5646,5647
for|5647,5650
an|5651,5653
aortic|5654,5660
arch|5661,5665
coarctation|5666,5677
.|5677,5678
The|5679,5682
aortic|5683,5689
<EOL>|5689,5690
valve|5690,5695
leaflets|5696,5704
(|5705,5706
?|5706,5707
#|5707,5708
)|5708,5709
appear|5710,5716
structurally|5717,5729
normal|5730,5736
.|5736,5737
There|5738,5743
is|5744,5746
no|5747,5749
<EOL>|5750,5751
aortic|5751,5757
valve|5758,5763
stenosis|5764,5772
.|5772,5773
There|5774,5779
is|5780,5782
no|5783,5785
aortic|5786,5792
<EOL>|5792,5793
regurgitation|5793,5806
.|5806,5807
The|5808,5811
mitral|5812,5818
valve|5819,5824
is|5825,5827
not|5828,5831
well|5832,5836
visualized|5837,5847
.|5847,5848
The|5849,5852
<EOL>|5853,5854
tricuspid|5854,5863
valve|5864,5869
is|5870,5872
not|5873,5876
well|5877,5881
seen|5882,5886
.|5886,5887
The|5888,5891
pulmonary|5892,5901
<EOL>|5901,5902
artery|5902,5908
systolic|5909,5917
pressure|5918,5926
could|5927,5932
not|5933,5936
be|5937,5939
estimated|5940,5949
.|5949,5950
There|5951,5956
is|5957,5959
no|5960,5962
<EOL>|5963,5964
pericardial|5964,5975
effusion|5976,5984
.|5984,5985
<EOL>|5985,5986
<EOL>|5986,5987
MICRO|5987,5992
:|5992,5993
<EOL>|5993,5994
=|5994,5995
=|5995,5996
=|5996,5997
=|5997,5998
=|5998,5999
=|5999,6000
<EOL>|6000,6001
_|6001,6002
_|6002,6003
_|6003,6004
1|6005,6006
:|6006,6007
05|6007,6009
am|6010,6012
FLUID|6013,6018
,|6018,6019
OTHER|6019,6024
PERICARDIAL|6030,6041
FLUID|6042,6047
.|6047,6048
<EOL>|6049,6050
<EOL>|6050,6051
GRAM|6054,6058
STAIN|6059,6064
(|6065,6066
Final|6066,6071
_|6072,6073
_|6073,6074
_|6074,6075
:|6075,6076
<EOL>|6077,6078
4|6084,6085
+|6085,6086
(|6089,6090
>|6090,6091
10|6091,6093
per|6094,6097
1000X|6098,6103
FIELD|6104,6109
)|6109,6110
:|6110,6111
POLYMORPHONUCLEAR|6114,6131
<EOL>|6132,6133
LEUKOCYTES|6133,6143
.|6143,6144
<EOL>|6145,6146
NO|6152,6154
MICROORGANISMS|6155,6169
SEEN|6170,6174
.|6174,6175
<EOL>|6176,6177
This|6183,6187
is|6188,6190
a|6191,6192
concentrated|6193,6205
smear|6206,6211
made|6212,6216
by|6217,6219
cytospin|6220,6228
method|6229,6235
,|6235,6236
<EOL>|6237,6238
please|6238,6244
refer|6245,6250
to|6251,6253
<EOL>|6253,6254
hematology|6260,6270
for|6271,6274
a|6275,6276
quantitative|6277,6289
white|6290,6295
blood|6296,6301
cell|6302,6306
count|6307,6312
.|6312,6313
.|6313,6314
<EOL>|6315,6316
<EOL>|6316,6317
FLUID|6320,6325
CULTURE|6326,6333
(|6334,6335
Preliminary|6335,6346
)|6346,6347
:|6347,6348
<EOL>|6349,6350
Reported|6356,6364
to|6365,6367
and|6368,6371
read|6372,6376
back|6377,6381
by|6382,6384
_|6385,6386
_|6386,6387
_|6387,6388
_|6389,6390
_|6390,6391
_|6391,6392
<EOL>|6393,6394
1|6394,6395
:|6395,6396
53PM|6396,6400
.|6400,6401
<EOL>|6402,6403
STAPHYLOCOCCUS|6409,6423
,|6423,6424
COAGULASE|6425,6434
NEGATIVE.|6435,6444
1|6448,6449
COLONY|6450,6456
ON|6457,6459
1|6460,6461
<EOL>|6462,6463
PLATE|6463,6468
.|6468,6469
<EOL>|6470,6471
<EOL>|6471,6472
ANAEROBIC|6475,6484
CULTURE|6485,6492
(|6493,6494
Preliminary|6494,6505
)|6505,6506
:|6506,6507
NO|6511,6513
ANAEROBES|6514,6523
ISOLATED|6524,6532
.|6532,6533
<EOL>|6534,6535
<EOL>|6535,6536
FUNGAL|6539,6545
CULTURE|6546,6553
(|6554,6555
Preliminary|6555,6566
)|6566,6567
:|6567,6568
<EOL>|6569,6570
<EOL>|6570,6571
ACID|6574,6578
FAST|6579,6583
SMEAR|6584,6589
(|6590,6591
Final|6591,6596
_|6597,6598
_|6598,6599
_|6599,6600
:|6600,6601
<EOL>|6602,6603
NO|6609,6611
ACID|6612,6616
FAST|6617,6621
BACILLI|6622,6629
SEEN|6630,6634
ON|6635,6637
DIRECT|6638,6644
SMEAR|6645,6650
.|6650,6651
<EOL>|6652,6653
<EOL>|6653,6654
ACID|6657,6661
FAST|6662,6666
CULTURE|6667,6674
(|6675,6676
Preliminary|6676,6687
)|6687,6688
:|6688,6689
<EOL>|6690,6691
<EOL>|6691,6692
DISCHARGE|6692,6701
LABS|6702,6706
:|6706,6707
<EOL>|6707,6708
=|6708,6709
=|6709,6710
=|6710,6711
=|6711,6712
=|6712,6713
=|6713,6714
=|6714,6715
=|6715,6716
=|6716,6717
=|6717,6718
=|6718,6719
=|6719,6720
=|6720,6721
=|6721,6722
=|6722,6723
<EOL>|6723,6724
_|6724,6725
_|6725,6726
_|6726,6727
04|6728,6730
:|6730,6731
01AM|6731,6735
BLOOD|6736,6741
WBC|6742,6745
-|6745,6746
13|6746,6748
.|6748,6749
0|6749,6750
*|6750,6751
RBC|6752,6755
-|6755,6756
4|6756,6757
.|6757,6758
05|6758,6760
*|6760,6761
Hgb|6762,6765
-|6765,6766
12|6766,6768
.|6768,6769
3|6769,6770
*|6770,6771
Hct|6772,6775
-|6775,6776
37|6776,6778
.|6778,6779
3|6779,6780
*|6780,6781
<EOL>|6782,6783
MCV|6783,6786
-|6786,6787
92|6787,6789
MCH|6790,6793
-|6793,6794
30.4|6794,6798
MCHC|6799,6803
-|6803,6804
33.0|6804,6808
RDW|6809,6812
-|6812,6813
13.0|6813,6817
RDWSD|6818,6823
-|6823,6824
43.8|6824,6828
Plt|6829,6832
_|6833,6834
_|6834,6835
_|6835,6836
<EOL>|6836,6837
_|6837,6838
_|6838,6839
_|6839,6840
03|6841,6843
:|6843,6844
30PM|6844,6848
BLOOD|6849,6854
Glucose|6855,6862
-|6862,6863
115|6863,6866
*|6866,6867
UreaN|6868,6873
-|6873,6874
22|6874,6876
*|6876,6877
Creat|6878,6883
-|6883,6884
0.6|6884,6887
Na|6888,6890
-|6890,6891
138|6891,6894
<EOL>|6895,6896
K|6896,6897
-|6897,6898
4.1|6898,6901
Cl|6902,6904
-|6904,6905
100|6905,6908
HCO3|6909,6913
-|6913,6914
24|6914,6916
AnGap|6917,6922
-|6922,6923
14|6923,6925
<EOL>|6925,6926
_|6926,6927
_|6927,6928
_|6928,6929
04|6930,6932
:|6932,6933
01AM|6933,6937
BLOOD|6938,6943
ALT|6944,6947
-|6947,6948
43|6948,6950
*|6950,6951
AST|6952,6955
-|6955,6956
27|6956,6958
AlkPhos|6959,6966
-|6966,6967
99|6967,6969
TotBili|6970,6977
-|6977,6978
0.5|6978,6981
<EOL>|6981,6982
_|6982,6983
_|6983,6984
_|6984,6985
03|6986,6988
:|6988,6989
30PM|6989,6993
BLOOD|6994,6999
Calcium|7000,7007
-|7007,7008
8|7008,7009
.|7009,7010
2|7010,7011
*|7011,7012
Phos|7013,7017
-|7017,7018
2.9|7018,7021
Mg|7022,7024
-|7024,7025
1.9|7025,7028
<EOL>|7028,7029
_|7029,7030
_|7030,7031
_|7031,7032
10|7033,7035
:|7035,7036
57PM|7036,7040
BLOOD|7041,7046
proBNP|7047,7053
-|7053,7054
110|7054,7057
<EOL>|7057,7058
_|7058,7059
_|7059,7060
_|7060,7061
03|7062,7064
:|7064,7065
29AM|7065,7069
BLOOD|7070,7075
TSH|7076,7079
-|7079,7080
0.93|7080,7084
<EOL>|7084,7085
_|7085,7086
_|7086,7087
_|7087,7088
11|7089,7091
:|7091,7092
04AM|7092,7096
BLOOD|7097,7102
_|7103,7104
_|7104,7105
_|7105,7106
pO2|7107,7110
-|7110,7111
82|7111,7113
*|7113,7114
pCO2|7115,7119
-|7119,7120
42|7120,7122
pH|7123,7125
-|7125,7126
7|7126,7127
.|7127,7128
34|7128,7130
*|7130,7131
<EOL>|7132,7133
calTCO2|7133,7140
-|7140,7141
24|7141,7143
Base|7144,7148
XS|7149,7151
-|7151,7152
-|7152,7153
2|7153,7154
<EOL>|7154,7155
<EOL>|7156,7157
SUMMARY|7180,7187
:|7187,7188
<EOL>|7189,7190
=|7190,7191
=|7191,7192
=|7192,7193
=|7193,7194
=|7194,7195
=|7195,7196
=|7196,7197
=|7197,7198
=|7198,7199
=|7199,7200
=|7200,7201
=|7201,7202
=|7202,7203
=|7203,7204
=|7204,7205
=|7205,7206
=|7206,7207
=|7207,7208
=|7208,7209
=|7209,7210
=|7210,7211
<EOL>|7212,7213
_|7213,7214
_|7214,7215
_|7215,7216
male|7217,7221
with|7222,7226
rheumatoid|7227,7237
arthritis|7238,7247
,|7247,7248
DMARD|7249,7254
holiday|7255,7262
,|7262,7263
and|7264,7267
<EOL>|7267,7268
recent|7268,7274
,|7274,7275
brief|7276,7281
hospitalization|7282,7297
for|7298,7301
presumptive|7302,7313
pericarditis|7314,7326
,|7326,7327
<EOL>|7327,7328
returned|7328,7336
to|7337,7339
outside|7340,7347
hospital|7348,7356
with|7357,7361
pericardial|7362,7373
effusion|7374,7382
with|7383,7387
<EOL>|7388,7389
possible|7389,7397
tamponade|7398,7407
physiology|7408,7418
now|7419,7422
post-bedside|7423,7435
<EOL>|7436,7437
pericardiocentesis|7437,7455
prior|7456,7461
to|7462,7464
transfer|7465,7473
,|7473,7474
with|7475,7479
persistent|7480,7490
<EOL>|7491,7492
pericardial|7492,7503
effusion|7504,7512
now|7513,7516
s|7517,7518
/|7518,7519
p|7519,7520
drain|7521,7526
placement|7527,7536
with|7537,7541
course|7542,7548
<EOL>|7549,7550
complicated|7550,7561
by|7562,7564
acute|7565,7570
hypercapneic|7571,7583
respiratory|7584,7595
distress|7596,7604
.|7604,7605
<EOL>|7606,7607
<EOL>|7607,7608
#|7608,7609
CORONARIES|7609,7619
:|7619,7620
unknown|7621,7628
.|7628,7629
<EOL>|7629,7630
#|7630,7631
PUMP|7631,7635
:|7635,7636
normal|7637,7643
biventricular|7644,7657
structure|7658,7667
and|7668,7671
function|7672,7680
.|7680,7681
<EOL>|7682,7683
#|7683,7684
RHYTHM|7684,7690
:|7690,7691
NSR|7692,7695
.|7695,7696
pAF|7697,7700
_|7701,7702
_|7702,7703
_|7703,7704
<EOL>|7704,7705
<EOL>|7705,7706
TRANSITIONAL|7706,7718
ISSUES|7719,7725
:|7725,7726
<EOL>|7726,7727
=|7727,7728
=|7728,7729
=|7729,7730
=|7730,7731
=|7731,7732
=|7732,7733
=|7733,7734
=|7734,7735
=|7735,7736
=|7736,7737
=|7737,7738
=|7738,7739
=|7739,7740
=|7740,7741
=|7741,7742
=|7742,7743
=|7743,7744
=|7744,7745
=|7745,7746
=|7746,7747
<EOL>|7747,7748
[|7748,7749
]|7749,7750
He|7751,7753
was|7754,7757
discharged|7758,7768
on|7769,7771
ibuprofen|7772,7781
600mg|7782,7787
TID|7788,7791
and|7792,7795
colchicine|7796,7806
0.6|7807,7810
mg|7810,7812
<EOL>|7813,7814
BID|7814,7817
for|7818,7821
his|7822,7825
inflammatory|7826,7838
pericarditis|7839,7851
.|7851,7852
He|7853,7855
should|7856,7862
continue|7863,7871
<EOL>|7872,7873
colchicine|7873,7883
for|7884,7887
3|7888,7889
months|7890,7896
.|7896,7897
He|7898,7900
should|7901,7907
have|7908,7912
his|7913,7916
ibuprofen|7917,7926
tapered|7927,7934
<EOL>|7935,7936
weekly|7936,7942
following|7943,7952
resolution|7953,7963
of|7964,7966
his|7967,7970
symptoms|7971,7979
over|7980,7984
3|7985,7986
weeks|7987,7992
to|7993,7995
<EOL>|7996,7997
reduce|7997,8003
the|8004,8007
risk|8008,8012
of|8013,8015
recurrence|8016,8026
.|8026,8027
<EOL>|8028,8029
[|8029,8030
]|8030,8031
He|8032,8034
was|8035,8038
discharged|8039,8049
on|8050,8052
a|8053,8054
PPI|8055,8058
and|8059,8062
should|8063,8069
continue|8070,8078
this|8079,8083
while|8084,8089
on|8090,8092
<EOL>|8093,8094
ibuprofen|8094,8103
.|8103,8104
<EOL>|8105,8106
[|8106,8107
]|8107,8108
Strongly|8109,8117
recommend|8118,8127
that|8128,8132
patient|8133,8140
receive|8141,8148
outpatient|8149,8159
PFTs|8160,8164
given|8165,8170
<EOL>|8171,8172
high|8172,8176
suspicion|8177,8186
for|8187,8190
baseline|8191,8199
obstructive|8200,8211
/|8211,8212
restrictive|8212,8223
pulmonary|8224,8233
<EOL>|8234,8235
disease|8235,8242
<EOL>|8243,8244
[|8244,8245
]|8245,8246
Patient|8247,8254
developed|8255,8264
paroxysmal|8265,8275
afib|8276,8280
with|8281,8285
RVR|8286,8289
during|8290,8296
this|8297,8301
<EOL>|8302,8303
admission|8303,8312
which|8313,8318
is|8319,8321
a|8322,8323
new|8324,8327
diagnosis|8328,8337
.|8337,8338
CHADSVASC|8339,8348
2|8349,8350
for|8351,8354
hypertension|8355,8367
<EOL>|8368,8369
and|8369,8372
diabetes|8373,8381
.|8381,8382
Anticoagulation|8383,8398
was|8399,8402
not|8403,8406
started|8407,8414
during|8415,8421
this|8422,8426
<EOL>|8427,8428
admission|8428,8437
given|8438,8443
that|8444,8448
he|8449,8451
was|8452,8455
felt|8456,8460
to|8461,8463
have|8464,8468
relatively|8469,8479
low|8480,8483
risk|8484,8488
for|8489,8492
<EOL>|8493,8494
CVA|8494,8497
,|8497,8498
however|8499,8506
please|8507,8513
make|8514,8518
a|8519,8520
note|8521,8525
of|8526,8528
this|8529,8533
new|8534,8537
diagnosis|8538,8547
and|8548,8551
<EOL>|8552,8553
reassess|8553,8561
need|8562,8566
for|8567,8570
anticoagulation|8571,8586
as|8587,8589
medically|8590,8599
appropriate|8600,8611
.|8611,8612
<EOL>|8613,8614
[|8614,8615
]|8615,8616
He|8617,8619
was|8620,8623
newly|8624,8629
diagnosed|8630,8639
with|8640,8644
DM|8645,8647
(|8648,8649
HbA1c|8649,8654
7.9|8655,8658
at|8659,8661
_|8662,8663
_|8663,8664
_|8664,8665
<EOL>|8666,8667
and|8667,8670
will|8671,8675
be|8676,8678
discharged|8679,8689
on|8690,8692
metformin|8693,8702
500|8703,8706
BID|8707,8710
.|8710,8711
Will|8712,8716
require|8717,8724
<EOL>|8725,8726
outpatient|8726,8736
follow|8737,8743
-|8743,8744
up|8744,8746
for|8747,8750
this|8751,8755
and|8756,8759
can|8760,8763
consider|8764,8772
uptitration|8773,8784
in|8785,8787
<EOL>|8788,8789
the|8789,8792
outpatient|8793,8803
setting|8804,8811
.|8811,8812
<EOL>|8813,8814
[|8814,8815
]|8815,8816
Please|8817,8823
reassess|8824,8832
need|8833,8837
for|8838,8841
diuretic|8842,8850
in|8851,8853
the|8854,8857
outpatient|8858,8868
setting|8869,8876
.|8876,8877
<EOL>|8878,8879
He|8879,8881
had|8882,8885
no|8886,8888
echocardiographic|8889,8906
evidence|8907,8915
of|8916,8918
heart|8919,8924
failure|8925,8932
during|8933,8939
<EOL>|8940,8941
this|8941,8945
admission|8946,8955
so|8956,8958
was|8959,8962
not|8963,8966
discharged|8967,8977
on|8978,8980
diuretics|8981,8990
.|8990,8991
<EOL>|8992,8993
<EOL>|8993,8994
New|8994,8997
medications|8998,9009
:|9009,9010
<EOL>|9010,9011
Metformin|9011,9020
500mg|9021,9026
BID|9027,9030
<EOL>|9030,9031
Metoprolol|9031,9041
XL|9042,9044
50mg|9045,9049
QD|9050,9052
<EOL>|9053,9054
Omeprazole|9054,9064
20mg|9065,9069
QD|9070,9072
<EOL>|9073,9074
<EOL>|9074,9075
Continued|9075,9084
medications|9085,9096
:|9096,9097
<EOL>|9097,9098
Atorvastatin|9098,9110
10mg|9111,9115
QPM|9116,9119
<EOL>|9119,9120
Colchicine|9120,9130
0.6|9131,9134
mg|9134,9136
BID|9137,9140
<EOL>|9140,9141
Ibuprofen|9141,9150
600mg|9151,9156
TID|9157,9160
<EOL>|9160,9161
Folic|9161,9166
acid|9167,9171
1mg|9172,9175
PO|9176,9178
QD|9179,9181
<EOL>|9181,9182
Sertraline|9182,9192
100mg|9193,9198
PO|9199,9201
QD|9202,9204
<EOL>|9204,9205
<EOL>|9205,9206
Stopped|9206,9213
medications|9214,9225
:|9225,9226
<EOL>|9227,9228
Methotrexate|9228,9240
20mg|9241,9245
PO|9246,9248
<EOL>|9248,9249
Famotidine|9249,9259
20mg|9260,9264
QD|9265,9267
<EOL>|9267,9268
<EOL>|9268,9269
ACUTE|9269,9274
ISSUES|9275,9281
:|9281,9282
<EOL>|9283,9284
=|9284,9285
=|9285,9286
=|9286,9287
=|9287,9288
=|9288,9289
=|9289,9290
=|9290,9291
=|9291,9292
=|9292,9293
=|9293,9294
=|9294,9295
=|9295,9296
=|9296,9297
<EOL>|9297,9298
#|9298,9299
)|9299,9300
Acute|9301,9306
pericarditis|9307,9319
<EOL>|9319,9320
#|9320,9321
)|9321,9322
Cardiac|9323,9330
tamponade|9331,9340
,|9340,9341
now|9342,9345
s|9346,9347
/|9347,9348
p|9348,9349
pericardiocentesis|9350,9368
and|9369,9372
drain|9373,9378
<EOL>|9378,9379
placement|9379,9388
<EOL>|9389,9390
He|9390,9392
presented|9393,9402
with|9403,9407
inflammatory|9408,9420
pericarditis|9421,9433
of|9434,9436
probable|9437,9445
viral|9446,9451
<EOL>|9452,9453
nature|9453,9459
in|9460,9462
the|9463,9466
context|9467,9474
of|9475,9477
viral|9478,9483
-|9483,9484
like|9484,9488
prodrome|9489,9497
versus|9498,9504
rheumatic|9505,9514
<EOL>|9515,9516
pericarditis|9516,9528
,|9528,9529
given|9530,9535
serologic|9536,9545
positive|9546,9554
active|9555,9561
disease|9562,9569
in|9570,9572
the|9573,9576
<EOL>|9577,9578
absence|9578,9585
of|9586,9588
DMARD|9589,9594
.|9594,9595
Pericardial|9596,9607
fluid|9608,9613
cultures|9614,9622
from|9623,9627
_|9628,9629
_|9629,9630
_|9630,9631
<EOL>|9632,9633
negative|9633,9641
,|9641,9642
cultures|9643,9651
here|9652,9656
with|9657,9661
1|9662,9663
colony|9664,9670
on|9671,9673
1|9674,9675
plate|9676,9681
of|9682,9684
coag|9685,9689
<EOL>|9690,9691
negative|9691,9699
staph|9700,9705
felt|9706,9710
to|9711,9713
be|9714,9716
contaminant|9717,9728
,|9728,9729
negative|9730,9738
acid|9739,9743
fast|9744,9748
smear|9749,9754
.|9754,9755
<EOL>|9756,9757
No|9757,9759
biochemical|9760,9771
evidence|9772,9780
of|9781,9783
myocardial|9784,9794
injury|9795,9801
on|9802,9804
admission|9805,9814
,|9814,9815
<EOL>|9816,9817
unlikely|9817,9825
to|9826,9828
have|9829,9833
concurrent|9834,9844
myocarditis|9845,9856
or|9857,9859
cardiac|9860,9867
event|9868,9873
<EOL>|9874,9875
sequelae|9875,9883
.|9883,9884
At|9885,9887
_|9888,9889
_|9889,9890
_|9890,9891
was|9892,9895
initially|9896,9905
noted|9906,9911
to|9912,9914
have|9915,9919
SBPs|9920,9924
in|9925,9927
<EOL>|9928,9929
the|9929,9932
_|9933,9934
_|9934,9935
_|9935,9936
and|9937,9940
received|9941,9949
fluid|9950,9955
resuscitation|9956,9969
and|9970,9973
pericardiocentesis|9974,9992
<EOL>|9993,9994
given|9994,9999
concern|10000,10007
for|10008,10011
tamponade|10012,10021
physiology|10022,10032
.|10032,10033
Hemodynamics|10034,10046
<EOL>|10047,10048
subsequently|10048,10060
stabilized|10061,10071
and|10072,10075
remained|10076,10084
so|10085,10087
throughout|10088,10098
the|10099,10102
duration|10103,10111
<EOL>|10112,10113
of|10113,10115
his|10116,10119
admission|10120,10129
here|10130,10134
.|10134,10135
TTE|10136,10139
on|10140,10142
_|10143,10144
_|10144,10145
_|10145,10146
showed|10147,10153
no|10154,10156
pericardial|10157,10168
<EOL>|10169,10170
effusion|10170,10178
.|10178,10179
Pericardial|10180,10191
drain|10192,10197
was|10198,10201
initially|10202,10211
left|10212,10216
to|10217,10219
gravity|10220,10227
due|10228,10231
to|10232,10234
<EOL>|10235,10236
continued|10236,10245
output|10246,10252
,|10252,10253
and|10254,10257
was|10258,10261
removed|10262,10269
_|10270,10271
_|10271,10272
_|10272,10273
.|10273,10274
He|10275,10277
was|10278,10281
treated|10282,10289
with|10290,10294
<EOL>|10295,10296
colchicine|10296,10306
0.6|10307,10310
mg|10310,10312
BID|10313,10316
which|10317,10322
he|10323,10325
will|10326,10330
continue|10331,10339
for|10340,10343
3|10344,10345
months|10346,10352
after|10353,10358
<EOL>|10359,10360
discharge|10360,10369
.|10369,10370
He|10371,10373
also|10374,10378
received|10379,10387
ibuprofen|10388,10397
600mg|10398,10403
PO|10404,10406
TID|10407,10410
and|10411,10414
will|10415,10419
be|10420,10422
<EOL>|10423,10424
discharged|10424,10434
on|10435,10437
a|10438,10439
slow|10440,10444
taper|10445,10450
;|10450,10451
he|10452,10454
received|10455,10463
PPI|10464,10467
while|10468,10473
receiving|10474,10483
<EOL>|10484,10485
NSAIDs|10485,10491
.|10491,10492
<EOL>|10493,10494
<EOL>|10494,10495
#|10495,10496
)|10496,10497
Acute|10498,10503
hypercapnic|10504,10515
respiratory|10516,10527
failure|10528,10535
-|10536,10537
resolving|10538,10547
<EOL>|10547,10548
Probable|10548,10556
flash|10557,10562
pulmonary|10563,10572
edema|10573,10578
from|10579,10583
rapid|10584,10589
large|10590,10595
-|10595,10596
volume|10596,10602
fluid|10603,10608
<EOL>|10609,10610
administration|10610,10624
on|10625,10627
tamponade|10628,10637
,|10637,10638
as|10639,10641
evidenced|10642,10651
by|10652,10654
radiographic|10655,10667
<EOL>|10668,10669
pulmonary|10669,10678
edema|10679,10684
.|10684,10685
Earlier|10686,10693
echocardiogram|10694,10708
otherwise|10709,10718
not|10719,10722
suggestive|10723,10733
<EOL>|10734,10735
of|10735,10737
ventricular|10738,10749
dysfunction|10750,10761
and|10762,10765
BNP|10766,10769
is|10770,10772
within|10773,10779
normal|10780,10786
limits.|10787,10794
TTE|10795,10798
<EOL>|10799,10800
on|10800,10802
_|10803,10804
_|10804,10805
_|10805,10806
was|10807,10810
without|10811,10818
evidence|10819,10827
of|10828,10830
cardiac|10831,10838
etiology|10839,10847
for|10848,10851
his|10852,10855
<EOL>|10856,10857
pulmonary|10857,10866
edema|10867,10872
/|10872,10873
respiratory|10873,10884
failure|10885,10892
.|10892,10893
<EOL>|10893,10894
Patient|10894,10901
likely|10902,10908
has|10909,10912
unappreciated|10913,10926
restrictive|10927,10938
pulmonary|10939,10948
<EOL>|10949,10950
physiology|10950,10960
.|10960,10961
Additionally|10962,10974
,|10974,10975
no|10976,10978
emphysematous|10979,10992
changes|10993,11000
noted|11001,11006
on|11007,11009
CT|11010,11012
<EOL>|11013,11014
one|11014,11017
week|11018,11022
ago|11023,11026
,|11026,11027
but|11028,11031
<EOL>|11031,11032
background|11032,11042
obstructive|11043,11054
defect|11055,11061
is|11062,11064
conceivable|11065,11076
,|11076,11077
given|11078,11083
compelling|11084,11094
<EOL>|11094,11095
smoking|11095,11102
history|11103,11110
.|11110,11111
He|11112,11114
had|11115,11118
a|11119,11120
negative|11121,11129
CTA|11130,11133
one|11134,11137
week|11138,11142
prior|11143,11148
to|11149,11151
<EOL>|11152,11153
admission|11153,11162
.|11162,11163
Patient|11164,11171
had|11172,11175
leukocytosis|11176,11188
on|11189,11191
admission|11192,11201
without|11202,11209
clear|11210,11215
<EOL>|11216,11217
radiographic|11217,11229
consolidation|11230,11243
suggestive|11244,11254
of|11255,11257
pneumonia|11258,11267
-|11268,11269
one|11270,11273
dose|11274,11278
of|11279,11281
<EOL>|11282,11283
empiric|11283,11290
azithromycin|11291,11303
was|11304,11307
given|11308,11313
overnight|11314,11323
and|11324,11327
discontinued|11328,11340
on|11341,11343
<EOL>|11344,11345
_|11345,11346
_|11346,11347
_|11347,11348
.|11348,11349
He|11350,11352
received|11353,11361
IV|11362,11364
diuresis|11365,11373
with|11374,11378
significant|11379,11390
improvement|11391,11402
in|11403,11405
<EOL>|11406,11407
his|11407,11410
respiratory|11411,11422
status|11423,11429
.|11429,11430
O2|11431,11433
weaned|11434,11440
_|11441,11442
_|11442,11443
_|11443,11444
morning|11445,11452
.|11452,11453
He|11454,11456
was|11457,11460
breathing|11461,11470
<EOL>|11471,11472
comfortably|11472,11483
on|11484,11486
RA|11487,11489
at|11490,11492
the|11493,11496
time|11497,11501
of|11502,11504
discharge|11505,11514
with|11515,11519
ambulatory|11520,11530
<EOL>|11531,11532
saturations|11532,11543
>|11544,11545
90|11545,11547
%|11547,11548
.|11548,11549
<EOL>|11550,11551
<EOL>|11551,11552
#|11552,11553
)|11553,11554
Paroxysmal|11555,11565
AFib|11566,11570
,|11570,11571
new|11572,11575
diagnosis|11576,11585
<EOL>|11586,11587
Patient|11587,11594
went|11595,11599
into|11600,11604
Afib|11605,11609
with|11610,11614
RVR|11615,11618
on|11619,11621
_|11622,11623
_|11623,11624
_|11624,11625
,|11625,11626
and|11627,11630
subsequently|11631,11643
<EOL>|11644,11645
received|11645,11653
metoprolol|11654,11664
.|11664,11665
He|11666,11668
subsequently|11669,11681
flipped|11682,11689
back|11690,11694
into|11695,11699
NSR|11700,11703
.|11703,11704
His|11705,11708
<EOL>|11709,11710
CHADsVASC|11710,11719
=|11720,11721
2|11722,11723
(|11724,11725
DM|11725,11727
,|11727,11728
HTN|11729,11732
)|11732,11733
.|11733,11734
Anticoagulation|11735,11750
was|11751,11754
discussed|11755,11764
but|11765,11768
<EOL>|11769,11770
ultimately|11770,11780
deferred|11781,11789
at|11790,11792
the|11793,11796
time|11797,11801
of|11802,11804
discharge|11805,11814
given|11815,11820
the|11821,11824
patient|11825,11832
's|11832,11834
<EOL>|11835,11836
lower|11836,11841
overall|11842,11849
risk|11850,11854
for|11855,11858
CVA|11859,11862
and|11863,11866
concerns|11867,11875
regarding|11876,11885
medication|11886,11896
<EOL>|11897,11898
adherence|11898,11907
/|11907,11908
cost|11908,11912
.|11912,11913
He|11914,11916
was|11917,11920
discharged|11921,11931
on|11932,11934
metoprolol|11935,11945
.|11945,11946
He|11947,11949
should|11950,11956
have|11957,11961
<EOL>|11962,11963
his|11963,11966
need|11967,11971
for|11972,11975
anticoagulation|11976,11991
reassessed|11992,12002
as|12003,12005
an|12006,12008
outpatient|12009,12019
as|12020,12022
<EOL>|12023,12024
medically|12024,12033
appropriate|12034,12045
.|12045,12046
<EOL>|12047,12048
<EOL>|12048,12049
#|12049,12050
)|12050,12051
Type|12052,12056
II|12057,12059
diabetes|12060,12068
:|12068,12069
<EOL>|12070,12071
He|12071,12073
was|12074,12077
newly|12078,12083
diagnosed|12084,12093
with|12094,12098
DM|12099,12101
with|12102,12106
a|12107,12108
A1C|12109,12112
of|12113,12115
7.9|12116,12119
%|12119,12120
during|12121,12127
this|12128,12132
<EOL>|12133,12134
admission|12134,12143
.|12143,12144
He|12145,12147
was|12148,12151
maintained|12152,12162
on|12163,12165
an|12166,12168
insulin|12169,12176
sliding|12177,12184
scale|12185,12190
during|12191,12197
<EOL>|12198,12199
this|12199,12203
admission|12204,12213
and|12214,12217
will|12218,12222
be|12223,12225
discharged|12226,12236
on|12237,12239
metformin|12240,12249
500mg|12250,12255
BID|12256,12259
.|12259,12260
<EOL>|12261,12262
<EOL>|12262,12263
CHRONIC|12263,12270
/|12270,12271
STABLE|12271,12277
ISSUES|12278,12284
:|12284,12285
<EOL>|12285,12286
=|12286,12287
=|12287,12288
=|12288,12289
=|12289,12290
=|12290,12291
=|12291,12292
=|12292,12293
=|12293,12294
=|12294,12295
=|12295,12296
=|12296,12297
=|12297,12298
=|12298,12299
=|12299,12300
=|12300,12301
=|12301,12302
=|12302,12303
=|12303,12304
=|12304,12305
=|12305,12306
<EOL>|12306,12307
#|12307,12308
)|12308,12309
Rheumatoid|12310,12320
arthritis|12321,12330
:|12330,12331
<EOL>|12332,12333
RF|12333,12335
and|12336,12339
anti-CCP|12340,12348
positive|12349,12357
per|12358,12361
outpatient|12362,12372
rheumatology|12373,12385
.|12385,12386
Not|12387,12390
<EOL>|12390,12391
currently|12391,12400
endorsing|12401,12410
sx|12411,12413
suggestive|12414,12424
of|12425,12427
RA|12428,12430
flare|12431,12436
.|12436,12437
Per|12438,12441
discussion|12442,12452
<EOL>|12452,12453
with|12453,12457
OP|12458,12460
rheumatologist|12461,12475
,|12475,12476
deferred|12477,12485
restarting|12486,12496
MTX|12497,12500
and|12501,12504
/|12504,12505
or|12505,12507
other|12508,12513
<EOL>|12513,12514
DMARD|12514,12519
until|12520,12525
outpatient|12526,12536
.|12536,12537
<EOL>|12537,12538
<EOL>|12538,12539
#|12539,12540
)|12540,12541
HTN|12542,12545
<EOL>|12545,12546
His|12546,12549
home|12550,12554
BP|12555,12557
meds|12558,12562
were|12563,12567
held|12568,12572
initially|12573,12582
due|12583,12586
to|12587,12589
soft|12590,12594
BPs|12595,12598
and|12599,12602
were|12603,12607
<EOL>|12608,12609
stopped|12609,12616
at|12617,12619
the|12620,12623
time|12624,12628
of|12629,12631
discharge|12632,12641
as|12642,12644
he|12645,12647
remained|12648,12656
normotensive|12657,12669
.|12669,12670
<EOL>|12671,12672
<EOL>|12672,12673
CORE|12673,12677
MEASURES|12678,12686
:|12686,12687
<EOL>|12688,12689
=|12689,12690
=|12690,12691
=|12691,12692
=|12692,12693
=|12693,12694
=|12694,12695
=|12695,12696
=|12696,12697
=|12697,12698
=|12698,12699
=|12699,12700
=|12700,12701
=|12701,12702
=|12702,12703
<EOL>|12704,12705
#|12705,12706
CODE|12706,12710
:|12710,12711
DNR|12712,12715
/|12715,12716
DNI|12716,12719
.|12719,12720
<EOL>|12720,12721
#|12721,12722
CONTACT|12722,12729
/|12729,12730
HCP|12730,12733
:|12733,12734
_|12735,12736
_|12736,12737
_|12737,12738
,|12738,12739
ex-wife|12740,12747
(|12748,12749
_|12749,12750
_|12750,12751
_|12751,12752
)|12752,12753
<EOL>|12754,12755
<EOL>|12756,12757
Medications|12757,12768
on|12769,12771
Admission|12772,12781
:|12781,12782
<EOL>|12782,12783
The|12783,12786
Preadmission|12787,12799
Medication|12800,12810
list|12811,12815
is|12816,12818
accurate|12819,12827
and|12828,12831
complete|12832,12840
.|12840,12841
<EOL>|12841,12842
1.|12842,12844
Atorvastatin|12845,12857
10|12858,12860
mg|12861,12863
PO|12864,12866
QPM|12867,12870
<EOL>|12871,12872
2.|12872,12874
Colchicine|12875,12885
0.6|12886,12889
mg|12890,12892
PO|12893,12895
BID|12896,12899
<EOL>|12900,12901
3.|12901,12903
Ibuprofen|12904,12913
600|12914,12917
mg|12918,12920
PO|12921,12923
TID|12924,12927
<EOL>|12928,12929
4.|12929,12931
Famotidine|12932,12942
20|12943,12945
mg|12946,12948
PO|12949,12951
DAILY|12952,12957
<EOL>|12958,12959
5.|12959,12961
lisinopril|12962,12972
-|12972,12973
hydrochlorothiazide|12973,12992
_|12993,12994
_|12994,12995
_|12995,12996
mg|12997,12999
oral|13000,13004
DAILY|13005,13010
<EOL>|13011,13012
6.|13012,13014
Methotrexate|13015,13027
20|13028,13030
mg|13031,13033
PO|13034,13036
1X|13037,13039
/|13039,13040
WEEK|13040,13044
(|13045,13046
_|13046,13047
_|13047,13048
_|13048,13049
)|13049,13050
<EOL>|13051,13052
7.|13052,13054
Sertraline|13055,13065
100|13066,13069
mg|13070,13072
PO|13073,13075
DAILY|13076,13081
<EOL>|13082,13083
8.|13083,13085
FoLIC|13086,13091
Acid|13092,13096
1|13097,13098
mg|13099,13101
PO|13102,13104
DAILY|13105,13110
<EOL>|13111,13112
<EOL>|13112,13113
<EOL>|13114,13115
Discharge|13115,13124
Medications|13125,13136
:|13136,13137
<EOL>|13137,13138
1.|13138,13140
Albuterol|13142,13151
Inhaler|13152,13159
2|13160,13161
PUFF|13162,13166
IH|13167,13169
Q6H|13170,13173
:|13173,13174
PRN|13174,13177
wheezing|13178,13186
,|13186,13187
shortness|13188,13197
of|13198,13200
<EOL>|13201,13202
breath|13202,13208
<EOL>|13209,13210
RX|13210,13212
*|13213,13214
albuterol|13214,13223
sulfate|13224,13231
[|13232,13233
ProAir|13233,13239
HFA|13240,13243
]|13243,13244
90|13245,13247
mcg|13248,13251
2|13252,13253
puffs|13254,13259
ih|13260,13262
every|13263,13268
6|13269,13270
<EOL>|13271,13272
hours|13272,13277
as|13278,13280
needed|13281,13287
Disp|13288,13292
#|13293,13294
*|13294,13295
1|13295,13296
Inhaler|13297,13304
Refills|13305,13312
:|13312,13313
*|13313,13314
0|13314,13315
<EOL>|13316,13317
2.|13317,13319
MetFORMIN|13321,13330
(|13331,13332
Glucophage|13332,13342
)|13342,13343
500|13344,13347
mg|13348,13350
PO|13351,13353
BID|13354,13357
<EOL>|13358,13359
RX|13359,13361
*|13362,13363
metformin|13363,13372
500|13373,13376
mg|13377,13379
1|13380,13381
tablet|13382,13388
(|13388,13389
s|13389,13390
)|13390,13391
by|13392,13394
mouth|13395,13400
Twice|13401,13406
a|13407,13408
day|13409,13412
Disp|13413,13417
#|13418,13419
*|13419,13420
60|13420,13422
<EOL>|13423,13424
Tablet|13424,13430
Refills|13431,13438
:|13438,13439
*|13439,13440
2|13440,13441
<EOL>|13442,13443
3.|13443,13445
Metoprolol|13447,13457
Succinate|13458,13467
XL|13468,13470
50|13471,13473
mg|13474,13476
PO|13477,13479
DAILY|13480,13485
<EOL>|13486,13487
RX|13487,13489
*|13490,13491
metoprolol|13491,13501
succinate|13502,13511
50|13512,13514
mg|13515,13517
1|13518,13519
tablet|13520,13526
(|13526,13527
s|13527,13528
)|13528,13529
by|13530,13532
mouth|13533,13538
Daily|13539,13544
Disp|13545,13549
<EOL>|13550,13551
#|13551,13552
*|13552,13553
30|13553,13555
Tablet|13556,13562
Refills|13563,13570
:|13570,13571
*|13571,13572
2|13572,13573
<EOL>|13574,13575
4.|13575,13577
Omeprazole|13579,13589
20|13590,13592
mg|13593,13595
PO|13596,13598
DAILY|13599,13604
<EOL>|13605,13606
RX|13606,13608
*|13609,13610
omeprazole|13610,13620
20|13621,13623
mg|13624,13626
1|13627,13628
capsule|13629,13636
(|13636,13637
s|13637,13638
)|13638,13639
by|13640,13642
mouth|13643,13648
Daily|13649,13654
Disp|13655,13659
#|13660,13661
*|13661,13662
30|13662,13664
<EOL>|13665,13666
Capsule|13666,13673
Refills|13674,13681
:|13681,13682
*|13682,13683
2|13683,13684
<EOL>|13685,13686
5.|13686,13688
Atorvastatin|13690,13702
10|13703,13705
mg|13706,13708
PO|13709,13711
QPM|13712,13715
<EOL>|13717,13718
6.|13718,13720
Colchicine|13722,13732
0.6|13733,13736
mg|13737,13739
PO|13740,13742
BID|13743,13746
<EOL>|13747,13748
RX|13748,13750
*|13751,13752
colchicine|13752,13762
0.6|13763,13766
mg|13767,13769
1|13770,13771
capsule|13772,13779
(|13779,13780
s|13780,13781
)|13781,13782
by|13783,13785
mouth|13786,13791
Twice|13792,13797
a|13798,13799
day|13800,13803
Disp|13804,13808
<EOL>|13809,13810
#|13810,13811
*|13811,13812
60|13812,13814
Capsule|13815,13822
Refills|13823,13830
:|13830,13831
*|13831,13832
2|13832,13833
<EOL>|13834,13835
7.|13835,13837
FoLIC|13839,13844
Acid|13845,13849
1|13850,13851
mg|13852,13854
PO|13855,13857
DAILY|13858,13863
<EOL>|13865,13866
8.|13866,13868
Ibuprofen|13870,13879
600|13880,13883
mg|13884,13886
PO|13887,13889
TID|13890,13893
<EOL>|13895,13896
9.|13896,13898
Sertraline|13900,13910
100|13911,13914
mg|13915,13917
PO|13918,13920
DAILY|13921,13926
<EOL>|13928,13929
10.|13929,13932
HELD|13933,13937
-|13937,13938
lisinopril|13939,13949
-|13949,13950
hydrochlorothiazide|13950,13969
_|13970,13971
_|13971,13972
_|13972,13973
mg|13974,13976
oral|13977,13981
DAILY|13982,13987
<EOL>|13989,13990
This|13990,13994
medication|13995,14005
was|14006,14009
held|14010,14014
.|14014,14015
Do|14016,14018
not|14019,14022
restart|14023,14030
<EOL>|14031,14032
lisinopril|14032,14042
-|14042,14043
hydrochlorothiazide|14043,14062
until|14063,14068
instructed|14069,14079
by|14080,14082
your|14083,14087
primary|14088,14095
<EOL>|14096,14097
care|14097,14101
doctor|14102,14108
or|14109,14111
cardiologist|14112,14124
<EOL>|14124,14125
11|14125,14127
.|14127,14128
HELD|14129,14133
-|14133,14134
Methotrexate|14135,14147
20|14148,14150
mg|14151,14153
PO|14154,14156
1X|14157,14159
/|14159,14160
WEEK|14160,14164
(|14165,14166
_|14166,14167
_|14167,14168
_|14168,14169
)|14169,14170
This|14172,14176
medication|14177,14187
<EOL>|14188,14189
was|14189,14192
held|14193,14197
.|14197,14198
Do|14199,14201
not|14202,14205
restart|14206,14213
Methotrexate|14214,14226
until|14227,14232
a|14233,14234
doctor|14235,14241
tells|14242,14247
you|14248,14251
<EOL>|14252,14253
to|14253,14255
<EOL>|14255,14256
<EOL>|14256,14257
<EOL>|14258,14259
Discharge|14259,14268
Disposition|14269,14280
:|14280,14281
<EOL>|14281,14282
Home|14282,14286
<EOL>|14286,14287
<EOL>|14288,14289
Discharge|14289,14298
Diagnosis|14299,14308
:|14308,14309
<EOL>|14309,14310
Primary|14310,14317
Diagnosis|14318,14327
:|14327,14328
inflammatory|14329,14341
pericarditis|14342,14354
<EOL>|14354,14355
Secondary|14355,14364
Diagnosis|14365,14374
:|14374,14375
rheumatoid|14376,14386
arthritis|14387,14396
<EOL>|14397,14398
<EOL>|14398,14399
<EOL>|14400,14401
Mental|14422,14428
Status|14429,14435
:|14435,14436
Clear|14437,14442
and|14443,14446
coherent|14447,14455
.|14455,14456
<EOL>|14456,14457
Level|14457,14462
of|14463,14465
Consciousness|14466,14479
:|14479,14480
Alert|14481,14486
and|14487,14490
interactive|14491,14502
.|14502,14503
<EOL>|14503,14504
Activity|14504,14512
Status|14513,14519
:|14519,14520
Ambulatory|14521,14531
-|14532,14533
Independent|14534,14545
.|14545,14546
<EOL>|14546,14547
<EOL>|14547,14548
<EOL>|14549,14550
Dear|14574,14578
Mr.|14579,14582
_|14583,14584
_|14584,14585
_|14585,14586
,|14586,14587
<EOL>|14589,14590
<EOL>|14591,14592
WHY|14592,14595
WERE|14596,14600
YOU|14601,14604
ADMITTED|14605,14613
TO|14614,14616
THE|14617,14620
HOSPITAL|14621,14629
?|14629,14630
<EOL>|14632,14633
-|14633,14634
You|14635,14638
were|14639,14643
admitted|14644,14652
to|14653,14655
the|14656,14659
hospital|14660,14668
with|14669,14673
chest|14674,14679
pain|14680,14684
.|14684,14685
<EOL>|14686,14687
<EOL>|14688,14689
WHAT|14689,14693
WAS|14694,14697
DONE|14698,14702
WHILE|14703,14708
YOU|14709,14712
WERE|14713,14717
IN|14718,14720
THE|14721,14724
HOSPITAL|14725,14733
?|14733,14734
<EOL>|14736,14737
-|14737,14738
You|14740,14743
were|14744,14748
found|14749,14754
to|14755,14757
have|14758,14762
inflammation|14763,14775
and|14776,14779
a|14780,14781
build|14782,14787
up|14788,14790
of|14791,14793
fluid|14794,14799
<EOL>|14800,14801
in|14801,14803
the|14804,14807
lining|14808,14814
of|14815,14817
the|14818,14821
heart|14822,14827
.|14827,14828
<EOL>|14828,14829
-|14829,14830
You|14831,14834
had|14835,14838
a|14839,14840
procedure|14841,14850
to|14851,14853
remove|14854,14860
the|14861,14864
fluid|14865,14870
from|14871,14875
the|14876,14879
lining|14880,14886
of|14887,14889
the|14890,14893
<EOL>|14894,14895
heart|14895,14900
and|14901,14904
a|14905,14906
temporary|14907,14916
drain|14917,14922
placed|14923,14929
.|14929,14930
This|14931,14935
was|14936,14939
removed|14940,14947
before|14948,14954
you|14955,14958
<EOL>|14959,14960
left|14960,14964
the|14965,14968
hospital|14969,14977
.|14977,14978
<EOL>|14979,14980
-|14980,14981
You|14982,14985
received|14986,14994
medication|14995,15005
to|15006,15008
help|15009,15013
you|15014,15017
pee|15018,15021
off|15022,15025
the|15026,15029
excess|15030,15036
fluid|15037,15042
<EOL>|15043,15044
in|15044,15046
your|15047,15051
body|15052,15056
.|15056,15057
<EOL>|15058,15059
-|15059,15060
You|15061,15064
developed|15065,15074
an|15075,15077
abnormal|15078,15086
heart|15087,15092
rhythm|15093,15099
(|15100,15101
afib|15101,15105
)|15105,15106
while|15107,15112
in|15113,15115
the|15116,15119
<EOL>|15120,15121
hospital|15121,15129
.|15129,15130
You|15131,15134
were|15135,15139
started|15140,15147
on|15148,15150
a|15151,15152
new|15153,15156
medication|15157,15167
for|15168,15171
this|15172,15176
<EOL>|15177,15178
(|15178,15179
metoprolol|15179,15189
)|15189,15190
.|15190,15191
<EOL>|15191,15192
-|15192,15193
You|15194,15197
were|15198,15202
diagnosed|15203,15212
with|15213,15217
diabetes|15218,15226
during|15227,15233
this|15234,15238
admission|15239,15248
.|15248,15249
You|15250,15253
<EOL>|15254,15255
were|15255,15259
started|15260,15267
on|15268,15270
a|15271,15272
new|15273,15276
medication|15277,15287
for|15288,15291
this|15292,15296
(|15297,15298
metformin|15298,15307
)|15307,15308
.|15308,15309
<EOL>|15310,15311
<EOL>|15312,15313
WHAT|15313,15317
DO|15318,15320
YOU|15321,15324
NEED|15325,15329
TO|15330,15332
DO|15333,15335
WHEN|15336,15340
YOU|15341,15344
LEAVE|15345,15350
THE|15351,15354
HOSPITAL|15355,15363
?|15363,15364
<EOL>|15366,15367
-|15367,15368
Take|15369,15373
all|15374,15377
of|15378,15380
your|15381,15385
medications|15386,15397
as|15398,15400
prescribed|15401,15411
(|15412,15413
listed|15413,15419
below|15420,15425
)|15425,15426
<EOL>|15428,15429
-|15429,15430
Follow|15431,15437
up|15438,15440
with|15441,15445
your|15446,15450
doctors|15451,15458
as|15459,15461
listed|15462,15468
below|15469,15474
<EOL>|15476,15477
-|15477,15478
Weigh|15479,15484
yourself|15485,15493
every|15494,15499
morning|15500,15507
,|15507,15508
seek|15509,15513
medical|15514,15521
attention|15522,15531
if|15532,15534
your|15535,15539
<EOL>|15540,15541
weight|15541,15547
goes|15548,15552
up|15553,15555
more|15556,15560
than|15561,15565
3|15566,15567
lbs|15568,15571
.|15571,15572
<EOL>|15574,15575
-|15575,15576
Seek|15577,15581
medical|15582,15589
attention|15590,15599
if|15600,15602
you|15603,15606
have|15607,15611
new|15612,15615
or|15616,15618
concerning|15619,15629
symptoms|15630,15638
<EOL>|15639,15640
or|15640,15642
you|15643,15646
develop|15647,15654
swelling|15655,15663
in|15664,15666
your|15667,15671
legs|15672,15676
,|15676,15677
abdominal|15678,15687
distention|15688,15698
,|15698,15699
or|15700,15702
<EOL>|15703,15704
shortness|15704,15713
of|15714,15716
breath|15717,15723
at|15724,15726
night|15727,15732
.|15732,15733
<EOL>|15735,15736
<EOL>|15736,15737
Please|15737,15743
see|15744,15747
below|15748,15753
for|15754,15757
more|15758,15762
information|15763,15774
on|15775,15777
your|15778,15782
hospitalization|15783,15798
.|15798,15799
<EOL>|15800,15801
It|15801,15803
was|15804,15807
a|15808,15809
pleasure|15810,15818
taking|15819,15825
part|15826,15830
in|15831,15833
your|15834,15838
care|15839,15843
here|15844,15848
at|15849,15851
_|15852,15853
_|15853,15854
_|15854,15855
!|15855,15856
<EOL>|15858,15859
<EOL>|15859,15860
We|15860,15862
wish|15863,15867
you|15868,15871
all|15872,15875
the|15876,15879
best|15880,15884
!|15884,15885
<EOL>|15887,15888
-|15889,15890
Your|15891,15895
_|15896,15897
_|15897,15898
_|15898,15899
Care|15900,15904
Team|15905,15909
<EOL>|15911,15912
<EOL>|15913,15914
Followup|15914,15922
Instructions|15923,15935
:|15935,15936
<EOL>|15936,15937
_|15937,15938
_|15938,15939
_|15939,15940
<EOL>|15940,15941

