 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Procedure|Health Care Activity|SIMPLE_SEGMENT|39,48|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|39,53|false|false|false|C2598112||Admission Date
Finding|Body Substance|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|73,82|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|73,82|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|73,87|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|105,110|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|129,132|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|129,132|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|140,147|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|140,147|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|149,157|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Attribute|Clinical Attribute|Allergies|181,190|false|false|false|C1717415||Allergies
Finding|Pathologic Function|Allergies|181,190|false|false|false|C0020517|Hypersensitivity|Allergies
Finding|Pathologic Function|Allergies|193,215|true|false|false|C0041755|Adverse reaction to drug|Adverse Drug Reactions
Drug|Pharmacologic Substance|Allergies|201,205|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|Drug
Finding|Finding|Allergies|201,205|false|false|false|C0740721|Drug problem|Drug
Finding|Pathologic Function|Allergies|201,215|true|false|false|C0041755|Adverse reaction to drug|Drug Reactions
Finding|Functional Concept|Allergies|218,227|false|false|false|C1999232|Attending (action)|Attending
Anatomy|Body Location or Region|Chief Complaint|253,256|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Chief Complaint|253,256|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Chief Complaint|253,256|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Finding|Classification|Chief Complaint|259,264|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|265,273|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|265,273|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|277,295|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|286,295|false|false|false|C0945766||Procedure
Event|Occupational Activity|Chief Complaint|286,295|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|286,295|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|286,295|false|false|false|C0184661|Interventional procedure|Procedure
Procedure|Diagnostic Procedure|Chief Complaint|297,300|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Finding|Idea or Concept|History of Present Illness|367,378|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|History of Present Illness|383,386|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|383,386|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|History of Present Illness|383,386|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|History of Present Illness|383,386|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|History of Present Illness|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|History of Present Illness|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|383,386|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|History of Present Illness|388,391|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|History of Present Illness|405,408|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|History of Present Illness|409,414|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|History of Present Illness|409,417|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|History of Present Illness|419,422|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|419,422|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|History of Present Illness|436,440|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|453,460|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|462,468|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|History of Present Illness|462,468|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Location or Region|History of Present Illness|485,490|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|History of Present Illness|485,490|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|485,499|false|false|false|C0230443|Structure of left lower leg|lower Left leg
Finding|Functional Concept|History of Present Illness|491,495|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|491,499|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|Left leg
Finding|Sign or Symptom|History of Present Illness|491,508|false|false|false|C2219779|numbness of left leg|Left leg numbness
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|496,499|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|History of Present Illness|496,508|false|true|false|C0857160|Numbness in leg|leg numbness
Finding|Finding|History of Present Illness|500,508|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|500,508|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|History of Present Illness|513,517|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|513,517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|513,517|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|548,556|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|548,556|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Disorder|Disease or Syndrome|History of Present Illness|579,582|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|History of Present Illness|579,582|false|false|false|C2346952|Bachelor of Education|bed
Attribute|Clinical Attribute|History of Present Illness|635,639|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|635,639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|635,639|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|640,648|false|false|false|C0026821|Muscle Cramp|cramping
Anatomy|Body Location or Region|History of Present Illness|667,671|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|667,671|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|697,701|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|History of Present Illness|697,701|false|false|false|C0555980|Foot problem|foot
Finding|Finding|History of Present Illness|737,744|false|false|false|C3888388|Usually|usually
Disorder|Disease or Syndrome|History of Present Illness|770,773|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|History of Present Illness|770,773|false|false|false|C2346952|Bachelor of Education|bed
Finding|Organism Function|History of Present Illness|785,793|false|false|false|C0015264|Exertion|exertion
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|806,809|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Finding|History of Present Illness|806,818|true|false|false|C0427068;C1836296|Monoparesis of lower limb;Muscle Weakness Lower Limb|leg weakness
Finding|Sign or Symptom|History of Present Illness|810,818|true|false|false|C0004093;C3714552|Asthenia;Weakness|weakness
Finding|Finding|History of Present Illness|827,831|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|History of Present Illness|827,831|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|History of Present Illness|827,831|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Finding|History of Present Illness|840,844|false|false|false|C1299581|Able (qualifier value)|able
Finding|Social Behavior|History of Present Illness|862,872|true|false|false|C0018896|Helping Behavior|assistance
Attribute|Clinical Attribute|History of Present Illness|884,888|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|884,888|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|884,888|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|History of Present Illness|893,901|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|893,901|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Finding|History of Present Illness|925,933|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|925,933|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Anatomy|Body Location or Region|History of Present Illness|949,953|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|949,953|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Location or Region|History of Present Illness|965,968|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|History of Present Illness|965,968|true|false|false|C2926618||DVT
Disorder|Disease or Syndrome|History of Present Illness|965,968|true|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|978,983|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Anatomy|Cell Component|History of Present Illness|978,983|false|false|false|C0037949;C2752558|Neuron spine;Vertebral column|spine
Finding|Finding|History of Present Illness|978,983|false|false|false|C0150920|Spine Problem|spine
Disorder|Injury or Poisoning|History of Present Illness|991,997|true|false|false|C1368081;C3263723;C3714660|Physical trauma;Trauma;Traumatic injury|trauma
Procedure|Health Care Activity|History of Present Illness|991,997|true|false|false|C0548346|Trauma assessment and care|trauma
Finding|Sign or Symptom|History of Present Illness|1002,1011|true|false|false|C0004604|Back Pain|back pain
Attribute|Clinical Attribute|History of Present Illness|1007,1011|true|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1007,1011|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1007,1011|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Disorder|Disease or Syndrome|History of Present Illness|1016,1028|true|false|false|C0021167|Incontinence|incontinence
Finding|Sign or Symptom|History of Present Illness|1034,1040|false|false|false|C0015967|Fever|fevers
Finding|Sign or Symptom|History of Present Illness|1041,1047|false|false|false|C0085593|Chills|chills
Finding|Finding|History of Present Illness|1052,1060|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1052,1060|true|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|History of Present Illness|1098,1106|false|false|false|C0018681|Headache|headache
Finding|Functional Concept|History of Present Illness|1108,1114|false|false|false|C0234621|Visual|visual
Finding|Finding|History of Present Illness|1108,1122|false|false|false|C0750280|Visual changes|visual changes
Finding|Functional Concept|History of Present Illness|1115,1122|false|false|false|C0392747|Changing|changes
Anatomy|Body Location or Region|History of Present Illness|1124,1129|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1124,1129|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1124,1134|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1124,1134|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1130,1134|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1130,1134|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1130,1134|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1130,1141|false|false|false|C0008031|Chest Pain|pain, chest
Anatomy|Body Location or Region|History of Present Illness|1136,1141|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1136,1141|false|false|false|C0741025|Chest problem|chest
Finding|Sign or Symptom|History of Present Illness|1136,1150|false|false|false|C0438716|Chest pressure|chest pressure
Finding|Finding|History of Present Illness|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|1142,1150|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|1142,1150|false|false|false|C0033095||pressure
Anatomy|Body Location or Region|History of Present Illness|1152,1157|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1152,1157|false|false|false|C0741025|Chest problem|chest
Finding|Finding|History of Present Illness|1159,1171|false|false|false|C0030252|Palpitations|palpitations
Attribute|Clinical Attribute|History of Present Illness|1173,1192|false|false|false|C2707305||shortness of breath
Finding|Sign or Symptom|History of Present Illness|1173,1192|false|false|false|C0013404|Dyspnea|shortness of breath
Finding|Body Substance|History of Present Illness|1186,1192|false|false|false|C0225386|Breath|breath
Anatomy|Body Location or Region|History of Present Illness|1193,1202|false|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1193,1207|false|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1203,1207|false|false|false|C2598155||pain
Finding|Functional Concept|History of Present Illness|1203,1207|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1203,1207|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1209,1216|false|false|false|C0013428|Dysuria|dysuria
Finding|Finding|History of Present Illness|1222,1230|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Finding|Sign or Symptom|History of Present Illness|1222,1230|false|false|false|C0011991;C2169706|Diarrhea;rectal discharge diarrhea (physical finding)|diarrhea
Disorder|Disease or Syndrome|Past Medical History|1259,1271|false|false|false|C0020538|Hypertensive disease|hypertension
Disorder|Disease or Syndrome|Past Medical History|1276,1284|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|diabetes
Disorder|Disease or Syndrome|Past Medical History|1292,1295|false|false|false|C0001365;C0038454|Acute ill-defined cerebrovascular disease;Cerebrovascular accident|CVA
Drug|Pharmacologic Substance|Past Medical History|1292,1295|false|false|false|C5779650|Cyclophosphamide/Doxorubicin/Vincristine|CVA
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1297,1307|false|false|false|C0007765|Cerebellum|cerebellar
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1308,1317|false|false|false|C0001629;C0025148;C1550278|Adrenal Medulla;Medulla Oblongata;Medullary - body parts|medullary
Disorder|Disease or Syndrome|Past Medical History|1318,1324|false|false|false|C0038454|Cerebrovascular accident|stroke
Finding|Finding|Past Medical History|1318,1324|false|false|false|C5977286|Stroke (heart beat)|stroke
Disorder|Disease or Syndrome|Past Medical History|1336,1339|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Past Medical History|1336,1339|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Past Medical History|1336,1339|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Past Medical History|1336,1339|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Past Medical History|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Past Medical History|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Past Medical History|1336,1339|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Past Medical History|1357,1360|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Disorder|Disease or Syndrome|Past Medical History|1392,1419|false|false|false|C0085096;C1704436|Peripheral Arterial Diseases;Peripheral Vascular Diseases|peripheral arterial disease
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1403,1411|false|false|false|C0003842|Arteries|arterial
Disorder|Disease or Syndrome|Past Medical History|1403,1419|false|false|false|C0852949|Arteriopathic disease|arterial disease
Disorder|Disease or Syndrome|Past Medical History|1412,1419|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Past Medical History|1421,1433|false|true|false|C0021775|Intermittent Claudication|claudication
Finding|Finding|Past Medical History|1421,1433|false|true|false|C0311395;C1456822|Claudication (finding);Lameness|claudication
Anatomy|Body Part, Organ, or Organ Component|Past Medical History|1448,1456|false|false|false|C0005847|Blood Vessel|vascular
Attribute|Clinical Attribute|Past Medical History|1483,1488|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Past Medical History|1483,1491|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Past Medical History|1492,1495|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Drug|Biomedical or Dental Material|Past Medical History|1497,1505|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Past Medical History|1497,1505|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Disease or Syndrome|Past Medical History|1519,1523|false|false|false|C0017168|Gastroesophageal reflux disease|GERD
Disorder|Disease or Syndrome|Past Medical History|1524,1534|false|false|false|C0014852|Esophageal Diseases|esophageal
Disorder|Disease or Syndrome|Past Medical History|1524,1540|false|false|false|C0267081|Terminal esophageal web|esophageal rings
Event|Activity|Family Medical History|1594,1598|false|false|false|C1947906|Sorting|sort
Finding|Cell Function|Family Medical History|1594,1598|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Finding|Mental Process|Family Medical History|1594,1598|false|false|false|C0237886;C0700314|Sorting (Cognition);Sorting - Cell Movement|sort
Disorder|Neoplastic Process|Family Medical History|1602,1608|false|false|false|C0006826|Malignant Neoplasms|cancer
Finding|Conceptual Entity|Family Medical History|1610,1616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Finding|Idea or Concept|Family Medical History|1610,1616|false|false|false|C1546503;C1547005;C2348513|Father - courtesy title;Indirect exposure mechanism - Father;Relationship - Father|Father
Anatomy|Body Location or Region|Family Medical History|1641,1645|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1641,1645|false|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|Family Medical History|1641,1645|false|false|false|C0024115|Lung diseases|lung
Finding|Finding|Family Medical History|1641,1645|false|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|Family Medical History|1641,1653|false|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|Family Medical History|1646,1653|false|false|false|C0012634|Disease|disease
Finding|Idea or Concept|Family Medical History|1656,1662|false|false|false|C1546508|Relationship - Mother|Mother
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Immunologic Factor|Family Medical History|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Drug|Pharmacologic Substance|Family Medical History|1689,1696|false|false|false|C1548502;C3541433|Unknown - Vaccines administered;unknown vaccine or immune globulin|unknown
Finding|Finding|Family Medical History|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Functional Concept|Family Medical History|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Idea or Concept|Family Medical History|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Intellectual Product|Family Medical History|1689,1696|false|false|false|C1546837;C1546841;C1547283;C1547294;C1547306;C1547312;C1548543;C1548550;C1549064;C1549105;C1549115;C1556120;C1556121;C1556122;C1556123;C1556124;C1556125;C1556126;C1556127;C1556128;C1556129;C1556130;C1556131;C1556132;C1556133;C1556134;C1556135;C1556136;C1556137;C1561529;C1609613;C3244284|Marital Status - Unknown;Unknown - Administrative Gender;Unknown - CWE statuses;Unknown - Contact Role;Unknown - Container status;Unknown - Employment Status;Unknown - Escort Required;Unknown - Event Expected;Unknown - Event reason;Unknown - Expanded yes/no indicator;Unknown - Immunization Registry Status;Unknown - Job Status;Unknown - Living Arrangement;Unknown - Living Dependency;Unknown - Living Will Code;Unknown - Notify Clergy Code;Unknown - Organ Donor Code;Unknown - Patient Class;Unknown - Patient Condition Code;Unknown - Patient Outcome;Unknown - Patient_s Relationship to Insured;Unknown - Precaution Code;Unknown - Production Class Code;Unknown - Recreational Drug Use Code;Unknown - Relationship;Unknown - Religion;Unknown - Special Program Code;Unknown - Transport Arranged;Unknown - mode of arrival code;Unknown - publishing section;Unknown Publicity Code;unknown - NullFlavor|unknown
Finding|Conceptual Entity|Family Medical History|1697,1702|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Finding|Functional Concept|Family Medical History|1697,1702|false|false|false|C0015127;C1524003|Etiology aspects;Science of Etiology|cause
Disorder|Disease or Syndrome|Family Medical History|1715,1718|true|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Family Medical History|1715,1718|true|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Family Medical History|1715,1718|true|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Family Medical History|1715,1718|true|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Family Medical History|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Family Medical History|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Family Medical History|1715,1718|true|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Finding|Pathologic Function|Family Medical History|1722,1742|true|false|false|C0085298|Sudden Cardiac Death|sudden cardiac death
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|1729,1736|false|false|false|C0018787|Heart|cardiac
Finding|Intellectual Product|Family Medical History|1729,1736|false|false|false|C1314974|Cardiac attachment|cardiac
Finding|Pathologic Function|Family Medical History|1729,1742|true|false|false|C0376297|Cardiac Death|cardiac death
Finding|Finding|Family Medical History|1737,1742|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Idea or Concept|Family Medical History|1737,1742|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Organism Function|Family Medical History|1737,1742|false|false|false|C0011065;C1306577;C1546949|Cessation of life;Death (finding);Event Consequence - Death|death
Finding|Conceptual Entity|Family Medical History|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Functional Concept|Family Medical History|1759,1766|true|false|false|C0019665;C0262512;C0262926;C1705255;C2004062|Concept History;Historical aspects qualifier;History of present illness (finding);History of previous events;Medical History|history
Finding|Finding|Family Medical History|1759,1769|true|false|false|C0262926|Medical History|history of
Disorder|Neoplastic Process|Family Medical History|1771,1777|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Health Care Activity|General Exam|1796,1805|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Finding|Finding|General Exam|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|1806,1814|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|1806,1814|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|1806,1819|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|1806,1819|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|General Exam|1815,1819|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|1815,1819|false|false|false|C0582103|Medical Examination|EXAM
Finding|Classification|General Exam|1866,1873|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|1866,1873|false|false|false|C3812897|General medical service|General
Finding|Mental Process|General Exam|1875,1883|false|false|false|C2987187|Pleasant|Pleasant
Finding|Mental Process|General Exam|1884,1890|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|1884,1890|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|General Exam|1902,1905|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|1902,1905|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|General Exam|1931,1934|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|1931,1934|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|1931,1934|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|1931,1934|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|1938,1943|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|1945,1951|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|1945,1951|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|1945,1951|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|1952,1961|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|1963,1966|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|1963,1966|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|1968,1978|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|1979,1984|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|General Exam|1992,1997|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|General Exam|2000,2004|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|2000,2004|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|2000,2004|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|General Exam|2006,2012|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|2014,2017|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Activity|General Exam|2046,2050|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|2046,2050|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|2055,2061|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2055,2061|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|General Exam|2082,2089|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|General Exam|2091,2095|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2108,2113|false|false|false|C0024109|Lung|Lungs
Finding|Finding|General Exam|2133,2141|false|false|false|C0034642;C0240859|Basilar Rales;Rales|crackles
Drug|Organic Chemical|General Exam|2156,2161|false|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|General Exam|2156,2161|false|false|false|C3815497|Cough (guaifenesin)|cough
Finding|Sign or Symptom|General Exam|2156,2161|false|false|false|C0010200|Coughing|cough
Anatomy|Body Location or Region|General Exam|2165,2172|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2165,2172|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|2165,2172|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2174,2179|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|2174,2187|false|false|false|C0426650|Obese abdomen|obese abdomen
Anatomy|Body Location or Region|General Exam|2180,2187|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|2180,2187|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|2180,2187|false|false|false|C0941288|Abdomen problem|abdomen
Disorder|Disease or Syndrome|General Exam|2189,2193|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|General Exam|2237,2245|false|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|General Exam|2249,2252|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|2249,2252|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|2254,2258|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2254,2258|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2260,2264|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|2278,2284|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|2278,2284|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|2278,2284|false|false|false|C0034107|Pulse taking|pulses
Finding|Functional Concept|General Exam|2286,2291|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|2286,2296|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|General Exam|2292,2296|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|2292,2296|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|General Exam|2292,2305|false|false|false|C0238882|Swollen calf|calf swelling
Finding|Finding|General Exam|2297,2305|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|2297,2305|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|General Exam|2320,2324|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|2320,2329|false|false|false|C0489800|Posterior part of left leg|left calf
Anatomy|Body Location or Region|General Exam|2325,2329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|2325,2329|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|General Exam|2325,2338|false|false|false|C0238882|Swollen calf|calf swelling
Finding|Finding|General Exam|2330,2338|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|2330,2338|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|General Exam|2343,2347|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|2343,2347|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|General Exam|2343,2358|true|false|false|C0238883|CALF TENDERNESS|calf tenderness
Finding|Mental Process|General Exam|2348,2358|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|2348,2358|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Procedure|Diagnostic Procedure|General Exam|2362,2371|false|false|false|C0030247|Palpation|palpation
Anatomy|Body Part, Organ, or Organ Component|General Exam|2380,2388|false|false|false|C0222007|Structure of nail of toe|toenails
Disorder|Disease or Syndrome|General Exam|2390,2398|false|false|false|C0043345|Xeroderma|dry skin
Drug|Pharmacologic Substance|General Exam|2390,2398|false|false|false|C0720057|Dry Skin brand of emollient|dry skin
Finding|Sign or Symptom|General Exam|2390,2398|false|false|false|C0151908|Dry skin|dry skin
Anatomy|Body System|General Exam|2394,2398|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|2394,2398|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|2394,2398|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Part, Organ, or Organ Component|General Exam|2405,2409|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Anatomy|Body Part, Organ, or Organ Component|General Exam|2411,2417|false|false|false|C0018534|Hallux structure|Hallux
Disorder|Acquired Abnormality|General Exam|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Anatomical Abnormality|General Exam|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Congenital Abnormality|General Exam|2411,2424|false|false|false|C0018536;C0158458;C0265656|Acquired hallux valgus;Congenital hallux valgus;Hallux Valgus|Hallux valgus
Disorder|Anatomical Abnormality|General Exam|2418,2424|false|false|false|C0042282|Valgus deformity|valgus
Finding|Finding|General Exam|2444,2450|false|false|false|C1554187|Gender Status - Intact|intact
Finding|Idea or Concept|General Exam|2456,2464|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|General Exam|2471,2476|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|2471,2476|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|2471,2488|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|2477,2488|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Finding|General Exam|2506,2515|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|2506,2515|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|2506,2515|false|false|false|C2229507|sensory exam|sensation
Finding|Body Substance|General Exam|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|2519,2528|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|2519,2528|false|false|false|C0030685|Patient Discharge|DISCHARGE
Finding|Finding|General Exam|2529,2537|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2529,2537|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2529,2537|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2529,2542|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2529,2542|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Finding|Functional Concept|General Exam|2538,2542|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2538,2542|false|false|false|C0582103|Medical Examination|EXAM
Attribute|Clinical Attribute|General Exam|2593,2597|false|false|false|C2317096|Saturation of Peripheral Oxygen|SpO2
Finding|Classification|General Exam|2620,2627|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|2620,2627|false|false|false|C3812897|General medical service|General
Finding|Mental Process|General Exam|2629,2637|false|false|false|C2987187|Pleasant|Pleasant
Finding|Mental Process|General Exam|2638,2644|false|false|false|C0001721|Affect (mental function)|affect
Procedure|Health Care Activity|General Exam|2638,2644|false|false|false|C2237113|assessment of affect|affect
Disorder|Disease or Syndrome|General Exam|2656,2659|false|false|false|C3159311|BORNHOLM EYE DISEASE|bed
Finding|Intellectual Product|General Exam|2656,2659|false|false|false|C2346952|Bachelor of Education|bed
Disorder|Disease or Syndrome|General Exam|2685,2688|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Disorder|Neoplastic Process|General Exam|2685,2688|false|false|false|C0205748;C0338473;C1850380|Dysplastic Nevus;NEUTROPHIL ACTIN DYSFUNCTION;Neuroaxonal Dystrophies|NAD
Drug|Biologically Active Substance|General Exam|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Drug|Pharmacologic Substance|General Exam|2685,2688|false|false|false|C0027270;C0621630|adenosine 5'-(alpha-thio)diphospho-5'-ribofuranosylnicotinamide;nicotinamide adenine dinucleotide (NAD)|NAD
Finding|Finding|General Exam|2685,2688|false|false|false|C2051415|patient appears in no acute distress (physical finding)|NAD
Anatomy|Body Location or Region|General Exam|2692,2697|false|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|2699,2705|false|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|2699,2705|false|false|false|C0036412|Scleral Diseases|Sclera
Procedure|Health Care Activity|General Exam|2699,2705|false|false|false|C2228481|examination of sclera|Sclera
Finding|Finding|General Exam|2706,2715|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|2717,2720|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|2717,2720|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|2722,2732|false|false|false|C0521367|Oropharyngeal|oropharynx
Finding|Idea or Concept|General Exam|2733,2738|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Finding|General Exam|2746,2751|false|false|false|C1642390|Pupil equal round and reacting to light|PERRL
Anatomy|Body Location or Region|General Exam|2754,2758|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|2754,2758|false|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|2754,2758|false|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Finding|Functional Concept|General Exam|2760,2766|false|false|false|C0332254|Supple|Supple
Finding|Finding|General Exam|2768,2771|false|false|false|C0428897|Jugular venous pressure|JVP
Event|Activity|General Exam|2800,2804|false|false|false|C0871208|Rating (action)|rate
Finding|Idea or Concept|General Exam|2800,2804|false|false|false|C1549480|Amount type - Rate|rate
Finding|Finding|General Exam|2809,2815|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2809,2815|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Finding|General Exam|2836,2843|true|false|false|C0018808|Heart murmur|murmurs
Finding|Finding|General Exam|2845,2849|true|false|false|C0232267|Pericardial friction rub|rubs
Anatomy|Body Part, Organ, or Organ Component|General Exam|2862,2867|false|false|false|C0024109|Lung|Lungs
Finding|Idea or Concept|General Exam|2869,2874|false|false|false|C1550016|Remote control command - Clear|clear
Procedure|Diagnostic Procedure|General Exam|2878,2890|false|false|false|C0004339|Auscultation|auscultation
Finding|Sign or Symptom|General Exam|2913,2920|true|false|false|C0043144|Wheezing|wheezes
Anatomy|Body Location or Region|General Exam|2932,2939|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|2932,2939|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|2932,2939|false|false|false|C0941288|Abdomen problem|Abdomen
Disorder|Disease or Syndrome|General Exam|2941,2946|false|false|false|C0028754|Obesity|obese
Finding|Finding|General Exam|2941,2954|false|false|false|C0426650|Obese abdomen|obese abdomen
Anatomy|Body Location or Region|General Exam|2947,2954|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|abdomen
Disorder|Neoplastic Process|General Exam|2947,2954|false|false|false|C0153662|Malignant neoplasm of abdomen|abdomen
Finding|Finding|General Exam|2947,2954|false|false|false|C0941288|Abdomen problem|abdomen
Disorder|Disease or Syndrome|General Exam|2956,2960|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Finding|Finding|General Exam|3004,3012|false|false|false|C0427198|Protective muscle spasm|guarding
Disorder|Congenital Abnormality|General Exam|3016,3019|false|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Finding|Gene or Genome|General Exam|3016,3019|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Finding|Finding|General Exam|3021,3025|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|3021,3025|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|3027,3031|false|false|false|C5575035|Well (answer to question)|well
Drug|Food|General Exam|3054,3060|false|false|false|C5890763||pulses
Finding|Physiologic Function|General Exam|3054,3060|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3054,3060|false|false|false|C0034107|Pulse taking|pulses
Attribute|Clinical Attribute|General Exam|3090,3095|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|General Exam|3090,3095|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|General Exam|3090,3095|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|General Exam|3090,3095|false|false|false|C0034107|Pulse taking|pulse
Attribute|Clinical Attribute|General Exam|3119,3124|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|General Exam|3119,3124|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|General Exam|3119,3124|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|General Exam|3119,3124|false|false|false|C0034107|Pulse taking|pulse
Finding|Conceptual Entity|General Exam|3136,3142|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Organ or Tissue Function|General Exam|3136,3148|false|false|false|C0232142||radial pulse
Procedure|Health Care Activity|General Exam|3136,3148|false|false|false|C2363059|examination of radial pulses|radial pulse
Attribute|Clinical Attribute|General Exam|3143,3148|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|General Exam|3143,3148|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|General Exam|3143,3148|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|General Exam|3143,3148|false|false|false|C0034107|Pulse taking|pulse
Finding|Finding|General Exam|3143,3151|false|false|false|C5238854|Pulse Wave Normal|pulse 2+
Finding|Conceptual Entity|General Exam|3155,3161|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Organ or Tissue Function|General Exam|3155,3167|false|false|false|C0232142||radial pulse
Procedure|Health Care Activity|General Exam|3155,3167|false|false|false|C2363059|examination of radial pulses|radial pulse
Attribute|Clinical Attribute|General Exam|3162,3167|false|false|false|C0232117|Pulse Rate|pulse
Finding|Physiologic Function|General Exam|3162,3167|false|false|false|C0391850|Physiologic pulse|pulse
Phenomenon|Phenomenon or Process|General Exam|3162,3167|false|false|false|C1947910|Pulse phenomenon|pulse
Procedure|Health Care Activity|General Exam|3162,3167|false|false|false|C0034107|Pulse taking|pulse
Finding|Finding|General Exam|3162,3170|false|false|false|C5238852|Pulse Wave Decreased|pulse 1+
Finding|Intellectual Product|General Exam|3172,3176|false|false|false|C1547225|Mild Severity of Illness Code|mild
Finding|Functional Concept|General Exam|3177,3182|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|3177,3187|false|false|false|C0489801|Posterior part of right leg|right calf
Anatomy|Body Location or Region|General Exam|3183,3187|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|3183,3187|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|General Exam|3183,3196|false|false|false|C0238882|Swollen calf|calf swelling
Finding|Finding|General Exam|3188,3196|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|3188,3196|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Functional Concept|General Exam|3211,3215|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|3211,3220|false|false|false|C0489800|Posterior part of left leg|left calf
Anatomy|Body Location or Region|General Exam|3216,3220|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|3216,3220|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Finding|General Exam|3216,3229|false|false|false|C0238882|Swollen calf|calf swelling
Finding|Finding|General Exam|3221,3229|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|3221,3229|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Anatomy|Body Location or Region|General Exam|3234,3238|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Anatomy|Body Part, Organ, or Organ Component|General Exam|3234,3238|false|false|false|C0230445;C1305418|Structure of calf of leg|calf
Finding|Sign or Symptom|General Exam|3234,3249|true|false|false|C0238883|CALF TENDERNESS|calf tenderness
Finding|Mental Process|General Exam|3239,3249|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3239,3249|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Procedure|Diagnostic Procedure|General Exam|3254,3263|false|false|false|C0030247|Palpation|palpation
Attribute|Clinical Attribute|General Exam|3268,3272|true|false|false|C2598155||pain
Finding|Functional Concept|General Exam|3268,3272|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|3268,3272|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Procedure|Diagnostic Procedure|General Exam|3276,3285|false|false|false|C0030247|Palpation|palpation
Finding|Functional Concept|General Exam|3289,3293|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3313,3317|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|General Exam|3313,3317|false|false|false|C0555980|Foot problem|foot
Disorder|Acquired Abnormality|General Exam|3321,3328|false|false|false|C0376154|Skin callus|callous
Finding|Finding|General Exam|3329,3336|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|3329,3336|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Functional Concept|General Exam|3340,3344|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|3353,3357|false|false|false|C0016504;C4299097|Foot;Lower extremity>Foot|foot
Finding|Finding|General Exam|3353,3357|false|false|false|C0555980|Foot problem|foot
Finding|Finding|General Exam|3359,3373|false|false|false|C4540337|Thick toenails|Thick toenails
Anatomy|Body Part, Organ, or Organ Component|General Exam|3365,3373|false|false|false|C0222007|Structure of nail of toe|toenails
Disorder|Disease or Syndrome|General Exam|3375,3383|false|false|false|C0043345|Xeroderma|dry skin
Drug|Pharmacologic Substance|General Exam|3375,3383|false|false|false|C0720057|Dry Skin brand of emollient|dry skin
Finding|Sign or Symptom|General Exam|3375,3383|false|false|false|C0151908|Dry skin|dry skin
Anatomy|Body System|General Exam|3379,3383|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|General Exam|3379,3383|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|General Exam|3379,3383|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|General Exam|3379,3383|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|General Exam|3379,3383|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Anatomy|Body Part, Organ, or Organ Component|General Exam|3391,3395|false|false|false|C0040357;C4299090|Lower extremity>Toes;Toes|toes
Finding|Functional Concept|General Exam|3408,3417|false|false|false|C0702114|indurated|indurated
Anatomy|Body Part, Organ, or Organ Component|General Exam|3418,3422|false|false|false|C1550235|Cord - Body Parts|cord
Disorder|Disease or Syndrome|General Exam|3418,3422|false|false|false|C3489532|Cone-Rod Dystrophy 2|cord
Finding|Functional Concept|General Exam|3426,3430|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|General Exam|3426,3448|false|false|false|C0694648|left antecubital fossa|left antecubital fossa
Anatomy|Body Part, Organ, or Organ Component|General Exam|3431,3442|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|General Exam|3431,3448|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|General Exam|3443,3448|false|false|false|C0836913|Fossa|fossa
Attribute|Clinical Attribute|General Exam|3457,3462|false|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3457,3462|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3457,3462|false|false|false|C0718338|Alert brand of caffeine|alert
Finding|Finding|General Exam|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3457,3462|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Finding|General Exam|3467,3475|false|false|false|C1961028|Oriented to place|oriented
Finding|Finding|General Exam|3490,3496|false|false|false|C1554187|Gender Status - Intact|intact
Drug|Organic Chemical|General Exam|3502,3505|false|false|false|C0939812|Ruta graveolens preparation|RUE
Drug|Pharmacologic Substance|General Exam|3502,3505|false|false|false|C0939812|Ruta graveolens preparation|RUE
Finding|Idea or Concept|General Exam|3512,3520|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Part, Organ, or Organ Component|General Exam|3530,3533|false|false|false|C0019552;C0022122;C0228391;C4299095|Bone structure of ischium;Hip structure;Lower extremity>Hip;Structure of habenulopeduncular tract|hip
Drug|Amino Acid, Peptide, or Protein|General Exam|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Biologically Active Substance|General Exam|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Drug|Pharmacologic Substance|General Exam|3530,3533|false|false|false|C0529134;C1430701;C1505163;C1654726|HHIP protein, human;RPL29 protein, human;ST13 protein, human;heme iron polypeptide|hip
Finding|Gene or Genome|General Exam|3530,3533|false|false|false|C1335638;C1337104;C1423009;C1538823;C1704840;C1709823;C3538851;C4284725|HHIP gene;HHIP wt Allele;REG3A gene;REG3A wt Allele;RPL29 gene;RPL29 wt Allele;ST13 gene;ST13 wt Allele|hip
Procedure|Therapeutic or Preventive Procedure|General Exam|3530,3533|false|false|false|C1292890|Procedure on hip|hip
Anatomy|Body Location or Region|General Exam|3534,3540|false|false|false|C1879367|Flexor (Anatomical coordinate)|flexor
Finding|Idea or Concept|General Exam|3541,3549|false|false|false|C0808080|Strength (attribute)|strength
Anatomy|Body Location or Region|General Exam|3565,3572|false|false|false|C0230463;C0442036|Plantar (qualifier value);Sole of Foot|plantar
Attribute|Clinical Attribute|General Exam|3574,3581|false|false|false|C1525443|W flexion|flexion
Finding|Organ or Tissue Function|General Exam|3574,3581|false|false|false|C0231452||flexion
Anatomy|Body Location or Region|General Exam|3595,3600|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|3595,3600|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|3595,3612|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|General Exam|3601,3612|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Finding|Functional Concept|General Exam|3622,3627|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Anatomy|Body Location or Region|General Exam|3628,3633|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|3628,3633|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|3635,3644|false|false|false|C0015385|Limb structure|extremity
Finding|Mental Process|General Exam|3663,3668|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|General Exam|3663,3668|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|General Exam|3663,3668|false|false|false|C0152054|Therapeutic Touch|touch
Finding|Organ or Tissue Function|General Exam|3663,3678|false|false|false|C0702221|Touch sensation|touch sensation
Finding|Finding|General Exam|3669,3678|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Finding|Organ or Tissue Function|General Exam|3669,3678|false|false|false|C0036658;C0542538|Observation of Sensation;Sensory perception|sensation
Procedure|Health Care Activity|General Exam|3669,3678|false|false|false|C2229507|sensory exam|sensation
Anatomy|Body Part, Organ, or Organ Component|General Exam|3682,3693|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Procedure|Health Care Activity|General Exam|3730,3739|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Lab|Laboratory or Test Result|General Exam|3740,3744|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3759,3764|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3759,3764|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3765,3768|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3773,3776|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3773,3776|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3773,3776|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3783,3786|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3783,3786|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3783,3786|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3783,3786|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3792,3795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3792,3795|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3803,3806|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|3803,3806|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3803,3806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3803,3806|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3810,3813|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3810,3813|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|3810,3813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3810,3813|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3810,3813|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3819,3823|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|3850,3853|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3870,3875|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|3870,3875|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3888,3894|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3901,3906|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3912,3915|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|3912,3915|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|4014,4019|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4014,4019|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4024,4027|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|General Exam|4024,4027|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4049,4054|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4049,4054|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4049,4062|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4049,4062|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4049,4062|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4055,4062|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4055,4062|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4055,4062|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|General Exam|4055,4062|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4055,4062|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|General Exam|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4110,4114|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4110,4114|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4140,4145|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4140,4145|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Amino Acid, Peptide, or Protein|General Exam|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Biologically Active Substance|General Exam|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Hormone|General Exam|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Drug|Pharmacologic Substance|General Exam|4171,4174|false|false|false|C0040162;C1702088;C3540580;C4521441|IL5 protein, human;Thyrotropin-Releasing Hormone, human;Tocotrienol-rich Fraction;thyrotropin-releasing hormone|TRF
Finding|Gene or Genome|General Exam|4171,4174|false|false|false|C1334121;C1336604;C1705002|IL5 gene;TERF1 gene;TERF1 wt Allele|TRF
Lab|Laboratory or Test Result|General Exam|4190,4194|false|false|false|C0587081|Laboratory test finding|LABS
Finding|Finding|General Exam|4195,4202|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4195,4202|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Drug|Amino Acid, Peptide, or Protein|General Exam|4222,4227|false|false|false|C2316467|Packed red blood cells|pRBCs
Drug|Pharmacologic Substance|General Exam|4222,4227|false|false|false|C2316467|Packed red blood cells|pRBCs
Procedure|Health Care Activity|General Exam|4231,4240|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Disease or Syndrome|General Exam|4256,4261|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4256,4261|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4262,4265|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4270,4273|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4270,4273|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4270,4273|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4280,4283|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4280,4283|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4280,4283|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4280,4283|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4289,4292|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4289,4292|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4300,4303|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4300,4303|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4300,4303|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4300,4303|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4307,4310|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4307,4310|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4307,4310|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4307,4310|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4307,4310|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4316,4320|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4347,4350|false|false|false|C0201617|Primed lymphocyte test|Plt
Finding|Gene or Genome|General Exam|4368,4373|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Food|General Exam|4385,4391|false|false|false|C0009237|Coffee|coffee
Finding|Finding|General Exam|4385,4405|false|false|false|C0278002;C1510416|Coffee ground vomiting;Vomit contains coffee grounds (finding)|coffee ground emesis
Finding|Sign or Symptom|General Exam|4385,4405|false|false|false|C0278002;C1510416|Coffee ground vomiting;Vomit contains coffee grounds (finding)|coffee ground emesis
Finding|Body Substance|General Exam|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|General Exam|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|General Exam|4399,4405|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Disorder|Disease or Syndrome|General Exam|4419,4424|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4419,4424|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4425,4428|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4433,4436|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4433,4436|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4433,4436|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4443,4446|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4443,4446|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4443,4446|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4443,4446|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4452,4455|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4452,4455|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4463,4466|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4463,4466|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4463,4466|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4463,4466|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4470,4473|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4470,4473|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4470,4473|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4470,4473|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4470,4473|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4479,4483|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4510,4513|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4566,4571|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|General Exam|4566,4571|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4572,4575|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4580,4583|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4580,4583|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4580,4583|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4591,4594|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4591,4594|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4591,4594|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4591,4594|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4602,4605|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4602,4605|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4613,4616|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|General Exam|4613,4616|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4613,4616|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4613,4616|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4620,4623|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4620,4623|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|General Exam|4620,4623|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4620,4623|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4620,4623|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4629,4633|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|General Exam|4660,4663|false|false|false|C0201617|Primed lymphocyte test|Plt
Anatomy|Body Location or Region|General Exam|4683,4688|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|General Exam|4683,4688|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|General Exam|4683,4698|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|General Exam|4689,4698|false|false|false|C0015385|Limb structure|extremity
Procedure|Diagnostic Procedure|General Exam|4699,4706|false|false|false|C0554756|Doppler studies|doppler
Attribute|Clinical Attribute|Impression|4729,4733|false|false|false|C4318566|Deep Resection Margin|Deep
Disorder|Disease or Syndrome|Impression|4729,4751|false|false|false|C0149871|Deep Vein Thrombosis|Deep venous thrombosis
Anatomy|Body Part, Organ, or Organ Component|Impression|4734,4740|false|false|false|C0042449|Veins|venous
Finding|Finding|Impression|4734,4751|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|Impression|4734,4751|false|false|false|C0042487;C0517555|Venous Thrombosis;Venous thrombosis after immobility|venous thrombosis
Finding|Pathologic Function|Impression|4741,4751|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|Impression|4769,4778|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|Impression|4779,4785|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|Impression|4787,4792|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Impression|4787,4792|false|false|false|C0398102|Procedure on vein|veins
Finding|Functional Concept|Impression|4818,4823|false|false|false|C1552823|Table Cell Horizontal Align - right|right
Disorder|Anatomical Abnormality|Impression|4834,4838|false|false|false|C0010709|Cyst|cyst
Finding|Body Substance|Impression|4834,4838|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Finding|Intellectual Product|Impression|4834,4838|false|false|false|C1546594;C1550626|SpecimenType - Cyst|cyst
Procedure|Diagnostic Procedure|Impression|4842,4845|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Finding|Intellectual Product|Impression|4856,4862|false|false|false|C1561574|Amount class - Amount|amount
Drug|Biologically Active Substance|Impression|4866,4873|false|false|false|C0018927|Hematin|hematin
Drug|Organic Chemical|Impression|4866,4873|false|false|false|C0018927|Hematin|hematin
Finding|Idea or Concept|Impression|4882,4890|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|4882,4893|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Pathologic Function|Impression|4894,4904|true|false|false|C0041582;C3887532|Ulcer;Ulceration|ulceration
Finding|Pathologic Function|Impression|4916,4924|false|false|false|C0019080|Hemorrhage|bleeding
Anatomy|Body Part, Organ, or Organ Component|Impression|4954,4961|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Impression|4954,4961|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Impression|4954,4961|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|Impression|4954,4961|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Impression|4954,4961|false|false|false|C0872393|Procedure on stomach|stomach
Disorder|Disease or Syndrome|Impression|4997,5005|false|false|false|C0041834|Erythema|erythema
Finding|Pathologic Function|Impression|5023,5034|false|false|false|C0041582|Ulcer|ulcerations
Anatomy|Body Part, Organ, or Organ Component|Impression|5042,5049|false|false|false|C0038351;C3714551;C4266636|Abdomen>Stomach;Stomach;Stomach structure|stomach
Disorder|Disease or Syndrome|Impression|5042,5049|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Disorder|Neoplastic Process|Impression|5042,5049|false|false|false|C0038354;C0153943;C0154060;C0496905|Benign neoplasm of stomach;Carcinoma in situ of stomach;Neoplasm of uncertain or unknown behavior of stomach;Stomach Diseases|stomach
Finding|Finding|Impression|5042,5049|false|false|false|C0577027|Stomach problem|stomach
Procedure|Therapeutic or Preventive Procedure|Impression|5042,5049|false|false|false|C0872393|Procedure on stomach|stomach
Finding|Idea or Concept|Impression|5050,5060|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|5050,5065|false|false|false|C0332290|Consistent with|consistent with
Finding|Finding|Impression|5066,5072|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Finding|Intellectual Product|Impression|5066,5072|false|false|false|C0205082;C1547227;C1547231;C1561581;C5203119|Allergy Severity - Severe;Intensity and Distress 5;Severe (severity modifier);Severe - Severity of Illness Code;Severe - Triage Code|severe
Disorder|Disease or Syndrome|Impression|5074,5083|false|false|false|C0017152|Gastritis|gastritis
Finding|Pathologic Function|Impression|5095,5103|true|false|false|C0019080|Hemorrhage|bleeding
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5116,5122|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|Medium
Drug|Substance|Impression|5116,5122|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|Medium
Finding|Finding|Impression|5116,5122|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|Medium
Finding|Intellectual Product|Impression|5116,5122|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|Medium
Disorder|Acquired Abnormality|Impression|5123,5136|false|false|false|C3489393|Hiatal Hernia|hiatal hernia
Disorder|Anatomical Abnormality|Impression|5130,5136|false|false|false|C0019270|Hernia|hernia
Disorder|Disease or Syndrome|Impression|5137,5145|false|false|false|C0041834|Erythema|Erythema
Finding|Pathologic Function|Impression|5162,5173|false|false|false|C0041582|Ulcer|ulcerations
Anatomy|Body Part, Organ, or Organ Component|Impression|5181,5189|false|false|false|C0013303|Duodenum|duodenal
Anatomy|Body Part, Organ, or Organ Component|Impression|5181,5194|false|false|false|C0227300|Duodenal ampulla|duodenal bulb
Anatomy|Anatomical Structure|Impression|5190,5194|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Anatomy|Body Part, Organ, or Organ Component|Impression|5190,5194|false|false|false|C0025148;C1947952|Medulla Oblongata;anatomical bulb|bulb
Finding|Idea or Concept|Impression|5196,5206|false|false|false|C0332290|Consistent with|consistent
Finding|Idea or Concept|Impression|5196,5211|false|false|false|C0332290|Consistent with|consistent with
Disorder|Disease or Syndrome|Impression|5212,5222|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Disorder|Neoplastic Process|Impression|5212,5222|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Procedure|Diagnostic Procedure|Impression|5241,5244|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Finding|Idea or Concept|Impression|5254,5258|false|false|false|C1552020|Role Class - part|part
Anatomy|Body Part, Organ, or Organ Component|Impression|5266,5274|false|false|false|C0013303|Duodenum|duodenum
Disorder|Neoplastic Process|Impression|5266,5274|false|false|false|C0153426;C0496869|Benign neoplasm of duodenum;Malignant neoplasm of duodenum|duodenum
Finding|Functional Concept|Impression|5280,5284|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Impression|5280,5300|false|false|false|C0230330|Left upper extremity|Left upper extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|5285,5300|false|false|false|C1140618|Upper Extremity|upper extremity
Anatomy|Body Part, Organ, or Organ Component|Impression|5291,5300|false|false|false|C0015385|Limb structure|extremity
Finding|Functional Concept|Impression|5301,5311|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Impression|5301,5311|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Impression|5301,5311|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Finding|Idea or Concept|Impression|5333,5341|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5333,5344|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Attribute|Clinical Attribute|Impression|5345,5349|true|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Impression|5345,5354|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|Impression|5345,5365|true|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Impression|5350,5354|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Impression|5350,5365|true|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|Impression|5355,5365|true|false|false|C0040053|Thrombosis|thrombosis
Finding|Functional Concept|Impression|5373,5377|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Impression|5385,5394|false|false|false|C0015385|Limb structure|extremity
Finding|Finding|Impression|5401,5407|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Idea or Concept|Impression|5401,5407|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|Likely
Finding|Functional Concept|Impression|5408,5416|false|true|false|C0332253|Evolving|evolving
Finding|Pathologic Function|Impression|5417,5425|false|true|false|C0018944|Hematoma|hematoma
Finding|Functional Concept|Impression|5433,5437|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Location or Region|Impression|5433,5455|false|false|false|C0694648|left antecubital fossa|left antecubital fossa
Anatomy|Body Part, Organ, or Organ Component|Impression|5438,5449|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|Impression|5438,5455|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|Impression|5450,5455|false|false|false|C0836913|Fossa|fossa
Attribute|Clinical Attribute|Impression|5463,5470|false|false|false|C0881943||CT head
Procedure|Diagnostic Procedure|Impression|5463,5470|false|false|false|C0202691|CAT scan of head|CT head
Anatomy|Body Location or Region|Impression|5466,5470|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|Impression|5466,5470|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|Impression|5466,5470|false|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|Impression|5466,5470|false|false|false|C0876917|Procedure on head|head
Drug|Indicator, Reagent, or Diagnostic Aid|Impression|5475,5483|false|false|false|C0009924|Contrast Media|contrast
Finding|Intellectual Product|Impression|5484,5494|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Mental Process|Impression|5484,5494|false|false|false|C0489484;C0596764|EKG impression;impression (attitude)|IMPRESSION
Finding|Idea or Concept|Impression|5502,5510|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Impression|5502,5513|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|Impression|5514,5519|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Impression|5520,5530|true|false|false|C0021308|Infarction|infarction
Finding|Pathologic Function|Impression|5532,5542|false|false|false|C0019080|Hemorrhage|hemorrhage
Disorder|Injury or Poisoning|Impression|5545,5554|false|false|false|C0016658|Fracture|fractures
Finding|Finding|Impression|5545,5554|false|false|false|C4554413|Fractured|fractures
Finding|Body Substance|Impression|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|Impression|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|Impression|5558,5567|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|Impression|5558,5567|false|false|false|C0030685|Patient Discharge|DISCHARGE
Lab|Laboratory or Test Result|Impression|5568,5572|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|Impression|5586,5591|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5586,5591|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|Impression|5592,5595|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|Impression|5600,5603|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|Impression|5600,5603|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|Impression|5600,5603|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|Impression|5610,5613|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|Impression|5610,5613|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|Impression|5610,5613|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|Impression|5610,5613|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|Impression|5619,5622|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|Impression|5619,5622|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|Impression|5630,5633|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Lab|Laboratory or Test Result|Impression|5630,5633|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|Impression|5630,5633|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|Impression|5630,5633|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|Impression|5637,5640|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|Impression|5637,5640|false|false|false|C0600370|methacholine|MCH
Finding|Gene or Genome|Impression|5637,5640|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|Impression|5637,5640|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|Impression|5637,5640|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|Impression|5646,5650|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Procedure|Laboratory Procedure|Impression|5677,5680|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|5697,5702|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5697,5702|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|5703,5706|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|Impression|5723,5728|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5723,5728|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|5723,5736|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|Impression|5723,5736|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|Impression|5723,5736|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|Impression|5729,5736|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|Impression|5729,5736|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|Impression|5729,5736|false|false|false|C0017725|glucose|Glucose
Lab|Laboratory or Test Result|Impression|5729,5736|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|Impression|5729,5736|false|false|false|C0337438|Glucose measurement|Glucose
Drug|Inorganic Chemical|Impression|5783,5787|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|Impression|5783,5787|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|Impression|5783,5787|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|Impression|5810,5815|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5810,5815|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|Impression|5810,5823|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|Impression|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|Impression|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|Impression|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|Impression|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|Impression|5816,5823|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Finding|Physiologic Function|Impression|5816,5823|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|Impression|5816,5823|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|Impression|5856,5861|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Finding|Body Substance|Impression|5856,5861|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|Impression|5862,5866|false|false|false|C0013618|edetic acid|EDTA
Drug|Pharmacologic Substance|Impression|5862,5866|false|false|false|C0013618|edetic acid|EDTA
Finding|Classification|Hospital Course|5896,5906|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Idea or Concept|Hospital Course|5896,5906|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|Outpatient
Finding|Functional Concept|Hospital Course|5907,5916|false|false|false|C1138603|Provider|Providers
Finding|Idea or Concept|Hospital Course|5932,5943|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Hospital Course|5948,5951|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|5948,5951|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|5948,5951|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|5948,5951|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5948,5951|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|5953,5956|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Hospital Course|5970,5973|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Hospital Course|5974,5979|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|5974,5982|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Hospital Course|5984,5987|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|5984,5987|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|Hospital Course|6001,6005|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6019,6026|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6019,6033|false|false|false|C0015801;C4299099|Lower extremity>Femoral artery;Structure of femoral artery|femoral artery
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6027,6033|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|6027,6033|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Location or Region|Hospital Course|6050,6055|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|6050,6055|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6050,6064|false|false|false|C0230443|Structure of left lower leg|lower left leg
Finding|Functional Concept|Hospital Course|6056,6060|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6056,6064|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|left leg
Finding|Sign or Symptom|Hospital Course|6056,6073|false|false|false|C2219779|numbness of left leg|left leg numbness
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6061,6064|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|6061,6073|false|false|false|C0857160|Numbness in leg|leg numbness
Finding|Finding|Hospital Course|6065,6073|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Hospital Course|6065,6073|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|Hospital Course|6078,6082|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|6078,6082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|6078,6082|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Anatomy|Body Location or Region|Hospital Course|6120,6123|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|6120,6123|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|6120,6123|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Drug|Biologically Active Substance|Hospital Course|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|6149,6156|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Pathologic Function|Hospital Course|6175,6183|false|false|false|C0019080|Hemorrhage|bleeding
Event|Event|Hospital Course|6184,6190|false|false|false|C0441471|Event|events
Procedure|Diagnostic Procedure|Hospital Course|6244,6247|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Procedure|Health Care Activity|Hospital Course|6284,6293|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biologically Active Substance|Hospital Course|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|6299,6306|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Intellectual Product|Hospital Course|6328,6332|false|false|false|C1720594|Then - dosing instruction fragment|then
Drug|Food|Hospital Course|6354,6360|false|false|false|C0009237|Coffee|coffee
Finding|Body Substance|Hospital Course|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|6368,6374|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Attribute|Clinical Attribute|Hospital Course|6389,6395|false|false|false|C0489144||stools
Finding|Body Substance|Hospital Course|6389,6395|false|false|false|C0015733|Feces|stools
Disorder|Cell or Molecular Dysfunction|Hospital Course|6408,6416|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|6408,6416|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|6408,6416|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|Hospital Course|6436,6441|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|6436,6441|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Drug|Biomedical or Dental Material|Hospital Course|6455,6461|false|false|false|C1272938|Rectal Dosage Form|rectal
Finding|Finding|Hospital Course|6455,6461|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Finding|Functional Concept|Hospital Course|6455,6461|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|rectal
Finding|Functional Concept|Hospital Course|6463,6467|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|6463,6467|false|false|false|C0582103|Medical Examination|exam
Procedure|Diagnostic Procedure|Hospital Course|6482,6493|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|6482,6493|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Body Substance|Hospital Course|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6519,6526|false|true|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|6558,6562|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6558,6566|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6563,6566|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|6563,6566|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Hospital Course|6563,6566|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6563,6566|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Pathologic Function|Hospital Course|6567,6575|false|false|false|C0018944|Hematoma|hematoma
Drug|Biologically Active Substance|Hospital Course|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|6581,6588|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Intellectual Product|Hospital Course|6611,6615|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Pathologic Function|Hospital Course|6636,6644|false|false|false|C0018944|Hematoma|hematoma
Finding|Intellectual Product|Hospital Course|6661,6667|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Functional Concept|Hospital Course|6677,6681|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Finding|Conceptual Entity|Hospital Course|6682,6688|false|false|false|C0442038;C0920847|Circumpennate;Radial|radial
Finding|Finding|Hospital Course|6692,6696|false|false|false|C5575035|Well (answer to question)|well
Anatomy|Body Location or Region|Hospital Course|6710,6715|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|6710,6715|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6710,6725|false|false|false|C0023216|Lower Extremity|lower extremity
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6716,6725|false|false|false|C0015385|Limb structure|extremity
Drug|Food|Hospital Course|6743,6749|false|false|false|C5890763||pulses
Finding|Physiologic Function|Hospital Course|6743,6749|false|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|Hospital Course|6743,6749|false|false|false|C0034107|Pulse taking|pulses
Procedure|Health Care Activity|Hospital Course|6761,6770|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Intellectual Product|Hospital Course|6772,6782|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|Hematology
Procedure|Laboratory Procedure|Hospital Course|6772,6782|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|Hematology
Finding|Body Substance|Hospital Course|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|6808,6815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|6828,6832|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6828,6836|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|6833,6836|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|6833,6836|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Hospital Course|6833,6836|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6833,6836|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Pathologic Function|Hospital Course|6837,6845|false|false|false|C0018944|Hematoma|hematoma
Finding|Idea or Concept|Hospital Course|6895,6910|false|false|false|C0034866|Recommendation|recommendations
Drug|Organic Chemical|Hospital Course|6945,6953|false|false|false|C0699129|Coumadin|coumadin
Drug|Pharmacologic Substance|Hospital Course|6945,6953|false|false|false|C0699129|Coumadin|coumadin
Attribute|Clinical Attribute|Hospital Course|6962,6965|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|6962,6965|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|6962,6965|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Body Substance|Hospital Course|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|6969,6978|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|6969,6978|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7010,7015|false|false|false|C0034991|Rehabilitation therapy|rehab
Attribute|Clinical Attribute|Hospital Course|7063,7070|false|false|false|C3854081||problem
Finding|Finding|Hospital Course|7063,7070|false|false|false|C0033213|Problem|problem
Finding|Intellectual Product|Hospital Course|7086,7093|false|false|false|C1552616;C1706244|Summary (document);summary - ActRelationshipSubset|summary
Finding|Idea or Concept|Hospital Course|7099,7111|false|false|false|C1548597|Marketing basis - Transitional|transitional
Finding|Idea or Concept|Hospital Course|7248,7259|false|false|false|C0750502|Significant|significant
Disorder|Disease or Syndrome|Hospital Course|7264,7267|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|7264,7267|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|7264,7267|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|7264,7267|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7264,7267|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|7269,7272|false|false|false|C0020538|Hypertensive disease|HTN
Disorder|Disease or Syndrome|Hospital Course|7285,7288|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Hospital Course|7290,7295|false|false|false|C1300072|Tumor stage|stage
Finding|Intellectual Product|Hospital Course|7290,7298|false|false|false|C0441772|Stage level 4|stage IV
Disorder|Disease or Syndrome|Hospital Course|7300,7303|false|false|false|C0085096|Peripheral Vascular Diseases|PVD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7300,7303|false|false|false|C4521226|Pomalidomide/Bortezomib/Dexamethasone Regimen|PVD
Finding|Functional Concept|Hospital Course|7317,7321|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7322,7348|false|false|false|C0447106|Superficial femoral artery|superficial femoral artery
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7334,7341|false|false|false|C0015811|Femur|femoral
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7334,7348|false|false|false|C0015801;C4299099|Lower extremity>Femoral artery;Structure of femoral artery|femoral artery
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7342,7348|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|7342,7348|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body Location or Region|Hospital Course|7367,7372|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|7367,7372|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7367,7381|false|false|false|C0230443|Structure of left lower leg|lower Left leg
Finding|Functional Concept|Hospital Course|7373,7377|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7373,7381|false|false|false|C0230416;C0230443|Left lower extremity;Structure of left lower leg|Left leg
Finding|Sign or Symptom|Hospital Course|7373,7390|false|true|false|C2219779|numbness of left leg|Left leg numbness
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7378,7381|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Sign or Symptom|Hospital Course|7378,7390|false|false|false|C0857160|Numbness in leg|leg numbness
Finding|Finding|Hospital Course|7382,7390|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Finding|Sign or Symptom|Hospital Course|7382,7390|false|false|false|C0020580;C0028643|Hypesthesia;Numbness|numbness
Attribute|Clinical Attribute|Hospital Course|7395,7399|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|7395,7399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|7395,7399|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Functional Concept|Hospital Course|7431,7441|false|false|false|C0220934|Ultrasonic|ultrasound
Phenomenon|Natural Phenomenon or Process|Hospital Course|7431,7441|false|false|false|C0041621;C1456803|Ultrasonic Shockwave;Ultrasonics (sound)|ultrasound
Procedure|Diagnostic Procedure|Hospital Course|7431,7441|false|false|false|C0041618;C1315081|Ultrasonography;Urological ultrasound|ultrasound
Anatomy|Body Location or Region|Hospital Course|7452,7457|false|false|false|C1548802|Body Site Modifier - Lower|lower
Event|Activity|Hospital Course|7452,7457|false|false|false|C2003888|Lower (action)|lower
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7452,7469|false|false|false|C0023216|Lower Extremity|lower extremities
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7458,7469|false|false|false|C0015385;C0278454|All extremities;Limb structure|extremities
Disorder|Disease or Syndrome|Hospital Course|7489,7498|false|false|false|C0751438|Posterior pituitary disease|posterior
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7489,7511|false|false|false|C0226832|Structure of posterior tibial vein|posterior tibial veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7499,7505|false|false|false|C0040184|Bone structure of tibia|tibial
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7499,7511|false|false|false|C0447138|Tibial vein structure|tibial veins
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|7506,7511|false|false|false|C0042449|Veins|veins
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7506,7511|false|false|false|C0398102|Procedure on vein|veins
Anatomy|Body Location or Region|Hospital Course|7512,7515|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|7512,7515|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|7512,7515|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Disease or Syndrome|Hospital Course|7543,7547|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Finding|Intellectual Product|Hospital Course|7552,7560|false|false|false|C1315013|Clinical NEC (not elsewhere classified in LNC)|clinical
Finding|Finding|Hospital Course|7561,7566|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|Hospital Course|7561,7566|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Procedure|Health Care Activity|Hospital Course|7577,7586|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Disorder|Cell or Molecular Dysfunction|Hospital Course|7603,7611|false|false|false|C4727483|BRAF Gene Rearrangement|positive
Finding|Classification|Hospital Course|7603,7611|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Finding|Finding|Hospital Course|7603,7611|false|false|false|C1446409;C1514241;C2699078|Positive;Positive Finding;Rh Positive Blood Group|positive
Disorder|Disease or Syndrome|Hospital Course|7622,7626|false|false|false|C0151950|Deep thrombophlebitis|DVTs
Attribute|Clinical Attribute|Hospital Course|7637,7641|false|false|false|C2598155||Pain
Finding|Functional Concept|Hospital Course|7637,7641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|Hospital Course|7637,7641|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Finding|Hospital Course|7647,7655|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Hospital Course|7647,7655|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Finding|Hospital Course|7668,7683|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|7668,7683|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7668,7683|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Body Substance|Hospital Course|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|7685,7692|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|Hospital Course|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|7711,7718|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7727,7738|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Hospital Course|7727,7738|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Finding|Functional Concept|Hospital Course|7727,7738|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Hospital Course|7727,7738|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7727,7738|false|false|false|C0087111|Therapeutic procedure|therapeutic
Drug|Hazardous or Poisonous Substance|Hospital Course|7739,7747|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|7739,7747|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|7739,7747|false|false|false|C0043031|warfarin|warfarin
Attribute|Clinical Attribute|Hospital Course|7753,7756|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|7753,7756|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|7753,7756|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Attribute|Clinical Attribute|Hospital Course|7753,7761|false|false|false|C5142654|Coagulation tissue factor induced.INR goal|INR goal
Finding|Idea or Concept|Hospital Course|7757,7761|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|Hospital Course|7757,7761|false|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Functional Concept|Hospital Course|7767,7770|false|false|false|C0678226;C3146286|Due;Due to|Due
Finding|Idea or Concept|Hospital Course|7767,7770|false|false|false|C0678226;C3146286|Due;Due to|Due
Disorder|Neoplastic Process|Hospital Course|7804,7807|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Hospital Course|7804,7807|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|Hospital Course|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|7817,7824|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Finding|Intellectual Product|Hospital Course|7832,7842|false|false|false|C1547985|Diagnostic Service Section ID - Hematology|hematology
Procedure|Laboratory Procedure|Hospital Course|7832,7842|false|false|false|C0018941;C0200627;C2183233|Hematologic Tests;Hematology procedure;diagnostic service sources hematology (procedure)|hematology
Drug|Biologically Active Substance|Hospital Course|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|Hospital Course|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|Hospital Course|7902,7909|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|Hospital Course|7952,7963|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|7952,7963|false|false|false|C0070166|clopidogrel|Clopidogrel
Finding|Classification|Hospital Course|7980,7990|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|7980,7990|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Body Substance|Hospital Course|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8005,8012|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Attribute|Clinical Attribute|Hospital Course|8024,8027|false|false|false|C1114365||age
Drug|Biologically Active Substance|Hospital Course|8024,8027|false|false|false|C0162574|Glycation End Products, Advanced|age
Drug|Organic Chemical|Hospital Course|8024,8027|false|false|false|C0162574|Glycation End Products, Advanced|age
Disorder|Neoplastic Process|Hospital Course|8040,8046|false|false|false|C0006826|Malignant Neoplasms|cancer
Procedure|Diagnostic Procedure|Hospital Course|8040,8056|false|false|false|C0199230|Screening for cancer|cancer screening
Finding|Finding|Hospital Course|8047,8056|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|Hospital Course|8047,8056|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|Hospital Course|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|Hospital Course|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|Hospital Course|8047,8056|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Diagnostic Procedure|Hospital Course|8067,8078|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|8067,8078|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Finding|Hospital Course|8084,8093|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|Hospital Course|8084,8093|false|false|false|C0024671|Mammography|mammogram
Finding|Body Substance|Hospital Course|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8095,8102|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|Hospital Course|8137,8152|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|8137,8152|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8137,8152|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Occupational Activity|Hospital Course|8153,8163|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|8153,8163|false|false|false|C0376636|Disease Management|management
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8184,8195|false|false|false|C0851145|on warfarin|on warfarin
Drug|Hazardous or Poisonous Substance|Hospital Course|8187,8195|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|8187,8195|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|8187,8195|false|false|false|C0043031|warfarin|warfarin
Procedure|Diagnostic Procedure|Hospital Course|8224,8232|false|false|false|C0203057|Upper gastrointestinal tract series|Upper GI
Finding|Pathologic Function|Hospital Course|8224,8238|false|false|false|C0041909|Upper gastrointestinal hemorrhage|Upper GI bleed
Finding|Pathologic Function|Hospital Course|8230,8238|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|8233,8238|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|Hospital Course|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8240,8247|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Gene or Genome|Hospital Course|8268,8273|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Drug|Food|Hospital Course|8274,8280|false|false|false|C0009237|Coffee|coffee
Finding|Body Substance|Hospital Course|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Physiologic Function|Hospital Course|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Finding|Sign or Symptom|Hospital Course|8289,8295|false|false|false|C0042963;C0042965;C2825053|Emesis [PE];Vomiting;Vomitus|emesis
Drug|Biologically Active Substance|Hospital Course|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8305,8312|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Disorder|Neoplastic Process|Hospital Course|8323,8326|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Hospital Course|8323,8326|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8347,8352|false|false|false|C2316467|Packed red blood cells|pRBCs
Drug|Pharmacologic Substance|Hospital Course|8347,8352|false|false|false|C2316467|Packed red blood cells|pRBCs
Procedure|Diagnostic Procedure|Hospital Course|8371,8374|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Disorder|Disease or Syndrome|Hospital Course|8382,8391|false|false|false|C0017152|Gastritis|gastritis
Disorder|Disease or Syndrome|Hospital Course|8409,8417|false|false|false|C0333307|Superficial ulcer|erosions
Finding|Pathologic Function|Hospital Course|8409,8417|false|false|false|C1959609|Erosion lesion|erosions
Finding|Pathologic Function|Hospital Course|8432,8440|true|false|false|C0019080|Hemorrhage|bleeding
Finding|Functional Concept|Hospital Course|8442,8452|false|false|false|C0444507|Incidental|Incidental
Finding|Finding|Hospital Course|8442,8460|false|false|false|C0743997|Incidental Findings|Incidental finding
Finding|Finding|Hospital Course|8453,8460|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Finding|Sign or Symptom|Hospital Course|8453,8460|false|false|false|C0037088;C0243095;C2825141|Experimental Finding;Finding;Signs and Symptoms|finding
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|8464,8470|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Drug|Substance|Hospital Course|8464,8470|false|false|false|C0010454;C1705217|Culture Media;Medium (Substance)|medium
Finding|Finding|Hospital Course|8464,8470|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Finding|Intellectual Product|Hospital Course|8464,8470|false|false|false|C0009458;C4522282;C4522283|A Medium Amount;A Medium Amount of Time;Communications Media|medium
Disorder|Acquired Abnormality|Hospital Course|8478,8491|false|false|false|C3489393|Hiatal Hernia|hiatal hernia
Disorder|Anatomical Abnormality|Hospital Course|8485,8491|false|false|false|C0019270|Hernia|hernia
Finding|Body Substance|Hospital Course|8493,8498|false|false|false|C0015733|Feces|Stool
Drug|Immunologic Factor|Hospital Course|8509,8516|false|false|false|C0003320|Antigens|antigen
Finding|Classification|Hospital Course|8521,8529|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|8521,8529|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|8521,8529|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|8558,8562|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Pharmacologic Substance|Hospital Course|8568,8571|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|8568,8571|false|false|false|C0871125|Prepulse Inhibition|PPI
Finding|Functional Concept|Hospital Course|8576,8580|false|false|false|C1552822|Table Cell Horizontal Align - left|Left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8581,8592|false|false|false|C1549091|Antecubital|antecubital
Finding|Pathologic Function|Hospital Course|8593,8601|false|false|false|C0018944|Hematoma|hematoma
Finding|Body Substance|Hospital Course|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8603,8610|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Gene or Genome|Hospital Course|8621,8626|false|false|false|C1416798;C5890938|LARGE1 gene;LARGE1 wt Allele|large
Finding|Functional Concept|Hospital Course|8627,8631|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|8633,8644|false|false|false|C1549091|Antecubital|antecubital
Finding|Pathologic Function|Hospital Course|8645,8653|false|true|false|C0018944|Hematoma|hematoma
Finding|Mental Process|Hospital Course|8657,8664|false|false|false|C0542559|contextual factors|setting
Finding|Finding|Hospital Course|8668,8678|false|false|false|C2183248|diagnostic service sources phlebotomy|phlebotomy
Procedure|Diagnostic Procedure|Hospital Course|8668,8678|false|false|false|C0031555;C0190979;C0684257|Phlebotomy, therapeutic (separate procedure);Venesection;Venous blood sampling|phlebotomy
Procedure|Therapeutic or Preventive Procedure|Hospital Course|8668,8678|false|false|false|C0031555;C0190979;C0684257|Phlebotomy, therapeutic (separate procedure);Venesection;Venous blood sampling|phlebotomy
Disorder|Neoplastic Process|Hospital Course|8683,8686|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Procedure|Laboratory Procedure|Hospital Course|8683,8686|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Drug|Biologically Active Substance|Hospital Course|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Organic Chemical|Hospital Course|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Drug|Pharmacologic Substance|Hospital Course|8697,8704|false|false|false|C0019134;C0770546|heparin;heparin, porcine|heparin
Disorder|Neoplastic Process|Hospital Course|8705,8708|false|false|false|C1135868|Gestational Trophoblastic Neoplasms|gtt
Drug|Biomedical or Dental Material|Hospital Course|8705,8708|false|false|false|C0991568|Drops - Drug Form|gtt
Procedure|Laboratory Procedure|Hospital Course|8705,8708|false|false|false|C0017741|Glucose tolerance test|gtt
Drug|Biologically Active Substance|Hospital Course|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Organic Chemical|Hospital Course|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Drug|Pharmacologic Substance|Hospital Course|8710,8717|false|false|false|C0019134;C0770546|heparin;heparin, porcine|Heparin
Finding|Pathologic Function|Hospital Course|8733,8741|false|false|false|C0018944|Hematoma|hematoma
Finding|Functional Concept|Hospital Course|8752,8758|false|false|false|C0205341;C1705914|Repeat;Repeat Object|Repeat
Finding|Intellectual Product|Hospital Course|8769,8775|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Intellectual Product|Hospital Course|8781,8786|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|Hospital Course|8790,8793|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Attribute|Clinical Attribute|Hospital Course|8794,8799|false|false|false|C1300072|Tumor stage|Stage
Finding|Intellectual Product|Hospital Course|8794,8802|false|false|false|C0441772|Stage level 4|Stage IV
Finding|Body Substance|Hospital Course|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|8804,8811|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Biologically Active Substance|Hospital Course|8817,8827|false|false|false|C0010294|creatinine|creatinine
Drug|Organic Chemical|Hospital Course|8817,8827|false|false|false|C0010294|creatinine|creatinine
Finding|Physiologic Function|Hospital Course|8817,8827|false|false|false|C4551889|Creatinine metabolic function|creatinine
Procedure|Laboratory Procedure|Hospital Course|8817,8827|false|false|false|C0201975|Creatinine measurement|creatinine
Procedure|Health Care Activity|Hospital Course|8839,8848|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Drug|Biomedical or Dental Material|Hospital Course|8854,8862|false|false|false|C0168634|BaseLine dental cement|baseline
Finding|Idea or Concept|Hospital Course|8854,8862|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Finding|Finding|Hospital Course|8886,8895|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Physiologic Function|Hospital Course|8886,8895|false|false|false|C1321013;C4520800|Hydration;Hydration status|hydration
Finding|Idea or Concept|Hospital Course|8897,8901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8897,8901|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8897,8901|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|8903,8908|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|8903,8908|false|false|false|C0699992|Lasix|lasix
Drug|Amino Acid, Peptide, or Protein|Hospital Course|8913,8923|false|false|false|C0065374|lisinopril|lisinopril
Drug|Pharmacologic Substance|Hospital Course|8913,8923|false|false|false|C0065374|lisinopril|lisinopril
Finding|Idea or Concept|Hospital Course|8945,8949|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|8945,8949|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|8945,8949|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|8950,8955|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|8950,8955|false|false|false|C0699992|Lasix|lasix
Finding|Body Substance|Hospital Course|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|8970,8979|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|8970,8979|false|false|false|C0030685|Patient Discharge|discharge
Disorder|Disease or Syndrome|Hospital Course|9010,9016|false|false|false|C0002871|Anemia|Anemia
Finding|Body Substance|Hospital Course|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|9018,9025|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Functional Concept|Hospital Course|9018,9029|false|false|false|C0332310|Has patient|Patient has
Disorder|Disease or Syndrome|Hospital Course|9041,9047|false|false|false|C0002871|Anemia|anemia
Drug|Biomedical or Dental Material|Hospital Course|9049,9055|false|false|false|C1272938|Rectal Dosage Form|Rectal
Finding|Finding|Hospital Course|9049,9055|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Finding|Functional Concept|Hospital Course|9049,9055|false|false|false|C1527425;C4521903|Rectal (intended site);Rectal Route of Administration|Rectal
Procedure|Diagnostic Procedure|Hospital Course|9049,9060|false|false|false|C0199900|Rectal examination|Rectal exam
Finding|Functional Concept|Hospital Course|9056,9060|false|false|false|C4284036|Exam|exam
Procedure|Health Care Activity|Hospital Course|9056,9060|false|false|false|C0582103|Medical Examination|exam
Drug|Indicator, Reagent, or Diagnostic Aid|Hospital Course|9072,9078|false|false|false|C0018302|guaiac|guaiac
Drug|Organic Chemical|Hospital Course|9072,9078|false|false|false|C0018302|guaiac|guaiac
Finding|Classification|Hospital Course|9079,9087|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|Hospital Course|9079,9087|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|Hospital Course|9079,9087|false|false|false|C5237010|Expression Negative|negative
Finding|Finding|Hospital Course|9121,9125|false|false|false|C5575035|Well (answer to question)|well
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Biologically Active Substance|Hospital Course|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Hormone|Hospital Course|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Drug|Pharmacologic Substance|Hospital Course|9130,9133|false|false|false|C0014822;C0357126;C2976467|EPO protein, human;Erythropoietin;epoetin alfa|EPO
Finding|Gene or Genome|Hospital Course|9130,9133|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|EPO
Finding|Intellectual Product|Hospital Course|9130,9133|false|false|false|C1366564;C1367459;C1414438;C1705819;C3496094|EPO gene;EPX gene;Exclusive Provider Organization Plan;TIMP1 gene;TIMP1 wt Allele|EPO
Finding|Conceptual Entity|Hospital Course|9135,9143|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Functional Concept|Hospital Course|9135,9143|false|false|false|C0015127;C1314792;C1524003|Etiology;Etiology aspects;Science of Etiology|Etiology
Finding|Finding|Hospital Course|9144,9150|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|9144,9150|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Drug|Organic Chemical|Hospital Course|9151,9158|false|false|false|C0163712|Relate - vinyl resin|related
Finding|Finding|Hospital Course|9151,9158|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Finding|Functional Concept|Hospital Course|9151,9158|false|false|false|C0445223;C1552599|Related (finding);Role Link Type - related|related
Disorder|Disease or Syndrome|Hospital Course|9173,9176|false|false|false|C1561643|Chronic Kidney Diseases|CKD
Finding|Pathologic Function|Hospital Course|9211,9219|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|9214,9219|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|Hospital Course|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9221,9228|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|9221,9232|false|false|false|C0332310|Has patient|patient has
Disorder|Disease or Syndrome|Hospital Course|9233,9242|false|false|false|C0017152|Gastritis|gastritis
Disorder|Disease or Syndrome|Hospital Course|9243,9253|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Disorder|Neoplastic Process|Hospital Course|9243,9253|false|false|false|C0013298;C1522057|Acute Enteritis of the Mouse Intestinal Tract;Duodenitis|duodenitis
Procedure|Diagnostic Procedure|Hospital Course|9258,9261|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Finding|Idea or Concept|Hospital Course|9269,9277|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|Hospital Course|9269,9280|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Pathologic Function|Hospital Course|9288,9296|true|false|false|C0019080|Hemorrhage|bleeding
Drug|Biologically Active Substance|Hospital Course|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Element, Ion, or Isotope|Hospital Course|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Drug|Pharmacologic Substance|Hospital Course|9298,9302|false|false|false|C0302583;C1166521;C3714701|Ferrum metallicum, Homeopathic preparation;Iron Drug Class;iron|Iron
Procedure|Laboratory Procedure|Hospital Course|9298,9302|false|false|false|C0337439|Iron measurement|Iron
Procedure|Laboratory Procedure|Hospital Course|9298,9310|false|false|false|C2079295|iron studies|Iron studies
Procedure|Research Activity|Hospital Course|9303,9310|false|false|false|C0947630|Scientific Study|studies
Finding|Idea or Concept|Hospital Course|9336,9340|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9336,9340|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9336,9340|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|9341,9351|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|9341,9351|false|false|false|C0016860|furosemide|furosemide
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9356,9366|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|9356,9366|false|false|false|C0065374|lisinopril|Lisinopril
Procedure|Health Care Activity|Hospital Course|9380,9389|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Pathologic Function|Hospital Course|9411,9419|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|9414,9419|false|false|false|C0019080|Hemorrhage|bleed
Drug|Organic Chemical|Hospital Course|9421,9431|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|9421,9431|false|false|false|C0054836|carvedilol|Carvedilol
Finding|Mental Process|Hospital Course|9459,9466|false|false|false|C0542559|contextual factors|setting
Finding|Idea or Concept|Hospital Course|9479,9484|false|false|false|C1552828|Table Frame - above|above
Drug|Organic Chemical|Hospital Course|9487,9497|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|Hospital Course|9487,9497|false|false|false|C0028066|nifedipine|Nifedipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9521,9524|false|false|false|C4546282|Body integrity dysphoria|bid
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9521,9524|false|false|false|C1530795|BID protein, human|bid
Drug|Biologically Active Substance|Hospital Course|9521,9524|false|false|false|C1530795|BID protein, human|bid
Finding|Gene or Genome|Hospital Course|9521,9524|false|false|false|C1332410|BID gene|bid
Drug|Organic Chemical|Hospital Course|9529,9534|false|false|false|C0699992|Lasix|lasix
Drug|Pharmacologic Substance|Hospital Course|9529,9534|false|false|false|C0699992|Lasix|lasix
Disorder|Disease or Syndrome|Hospital Course|9577,9580|false|false|false|C0010068;C0175816;C1956346|Cold Hemagglutinin Disease;Coronary Artery Disease;Coronary heart disease|CAD
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9577,9580|false|false|false|C1504769|DFFB protein, human|CAD
Drug|Enzyme|Hospital Course|9577,9580|false|false|false|C1504769|DFFB protein, human|CAD
Finding|Gene or Genome|Hospital Course|9577,9580|false|false|false|C1413078;C1413983;C1428349;C2239547;C3813548;C4284121|ACOD1 gene;B4GALNT2 gene;CAD gene;CALD1 wt Allele;DFFB gene;DFFB wt Allele|CAD
Procedure|Diagnostic Procedure|Hospital Course|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Research Activity|Hospital Course|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9577,9580|false|false|false|C0011905;C0170509;C0280573;C1707433|Collision-Induced Dissociation;Computer Assisted Diagnosis;CyADIC regimen;cytarabine/daunorubicin protocol|CAD
Disorder|Disease or Syndrome|Hospital Course|9598,9601|false|false|false|C0006430|Burning Mouth Syndrome|BMS
Anatomy|Body Location or Region|Hospital Course|9630,9633|false|false|false|C0449201|PER (body structure)|Per
Disorder|Disease or Syndrome|Hospital Course|9630,9633|false|false|false|C1861457|PROGRESSIVE ENCEPHALOMYELITIS WITH RIGIDITY|Per
Finding|Functional Concept|Hospital Course|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Gene or Genome|Hospital Course|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Finding|Intellectual Product|Hospital Course|9630,9633|false|false|false|C1418464;C1704764;C3273590;C4281991|Follow;PER1 gene;PER1 wt Allele;Per - dosing instruction fragment|Per
Procedure|Therapeutic or Preventive Procedure|Hospital Course|9635,9646|false|false|false|C0557061|Discussion (procedure)|discussions
Finding|Body Substance|Hospital Course|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|9661,9668|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Drug|Organic Chemical|Hospital Course|9686,9697|false|false|false|C0070166|clopidogrel|clopidogrel
Drug|Pharmacologic Substance|Hospital Course|9686,9697|false|false|false|C0070166|clopidogrel|clopidogrel
Finding|Pathologic Function|Hospital Course|9713,9721|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|9716,9721|false|false|false|C0019080|Hemorrhage|bleed
Finding|Functional Concept|Hospital Course|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Genetic Function|Hospital Course|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Finding|Mental Process|Hospital Course|9726,9736|false|false|false|C0589507;C1158830;C1704686|Initiation;Transcription Initiation|initiation
Drug|Hazardous or Poisonous Substance|Hospital Course|9740,9748|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|9740,9748|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Hospital Course|9740,9748|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Hospital Course|9751,9756|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|9751,9756|false|false|false|C0699992|Lasix|Lasix
Finding|Idea or Concept|Hospital Course|9775,9780|false|false|false|C1552828|Table Frame - above|above
Finding|Body Substance|Hospital Course|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|9799,9808|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|9799,9808|false|false|false|C0030685|Patient Discharge|discharge
Finding|Idea or Concept|Hospital Course|9825,9829|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9825,9829|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9825,9829|false|false|false|C1553498|home health encounter|Home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|9830,9833|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|Hospital Course|9830,9833|false|false|false|C1412553|ARSA gene|ASA
Drug|Organic Chemical|Hospital Course|9835,9841|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Drug|Pharmacologic Substance|Hospital Course|9835,9841|false|false|false|C0360714|Hydroxymethylglutaryl-CoA Reductase Inhibitors|statin
Finding|Gene or Genome|Hospital Course|9835,9841|false|false|false|C1414273|EEF1A2 gene|statin
Drug|Organic Chemical|Hospital Course|9847,9857|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|9847,9857|false|false|false|C0054836|carvedilol|carvedilol
Disorder|Disease or Syndrome|Hospital Course|9878,9881|false|false|false|C0020538|Hypertensive disease|HTN
Drug|Organic Chemical|Hospital Course|9883,9893|false|false|false|C0028066|nifedipine|Nifedipine
Drug|Pharmacologic Substance|Hospital Course|9883,9893|false|false|false|C0028066|nifedipine|Nifedipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9916,9919|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9916,9919|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9916,9919|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9916,9919|false|false|false|C1332410|BID gene|BID
Disorder|Mental or Behavioral Dysfunction|Hospital Course|9930,9933|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|9930,9933|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|9930,9933|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|9930,9933|false|false|false|C1332410|BID gene|BID
Finding|Pathologic Function|Hospital Course|9950,9958|false|false|false|C0019080|Hemorrhage|bleeding
Finding|Finding|Hospital Course|9950,9967|false|false|false|C1970394|Bleeding episodes|bleeding episodes
Disorder|Disease or Syndrome|Hospital Course|9979,9984|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Hospital Course|9979,9984|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Hospital Course|9979,9994|false|false|false|C1272641|Systemic arterial pressure|blood pressures
Finding|Finding|Hospital Course|9985,9994|false|false|false|C0460139|Pressure (finding)|pressures
Phenomenon|Phenomenon or Process|Hospital Course|9985,9994|false|false|false|C0033095||pressures
Finding|Idea or Concept|Hospital Course|9996,10000|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|Hospital Course|9996,10000|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|Hospital Course|9996,10000|false|false|false|C1553498|home health encounter|Home
Drug|Organic Chemical|Hospital Course|10002,10012|false|false|false|C0054836|carvedilol|carvedilol
Drug|Pharmacologic Substance|Hospital Course|10002,10012|false|false|false|C0054836|carvedilol|carvedilol
Finding|Body Substance|Hospital Course|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10024,10031|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|10034,10044|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10034,10044|false|false|false|C0028066|nifedipine|nifedipine
Finding|Intellectual Product|Hospital Course|10080,10085|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Hospital Course|10080,10091|false|false|false|C0333276|Acute hemorrhage|acute bleed
Finding|Pathologic Function|Hospital Course|10086,10091|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Space or Junction|Hospital Course|10096,10100|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Drug|Organic Chemical|Hospital Course|10112,10117|false|false|false|C0699992|Lasix|Lasix
Drug|Pharmacologic Substance|Hospital Course|10112,10117|false|false|false|C0699992|Lasix|Lasix
Disorder|Disease or Syndrome|Hospital Course|10163,10171|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Hospital Course|10163,10180|false|false|false|C0011849|Diabetes Mellitus|Diabetes Mellitus
Finding|Intellectual Product|Hospital Course|10182,10188|false|false|false|C1547311|Patient Condition Code - Stable|Stable
Finding|Idea or Concept|Hospital Course|10192,10196|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10192,10196|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10192,10196|false|false|false|C1553498|home health encounter|home
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|Hospital Course|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|Hospital Course|10212,10219|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Finding|Gene or Genome|Hospital Course|10212,10219|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|Hospital Course|10212,10219|false|false|false|C0202098|Insulin measurement|insulin
Finding|Idea or Concept|Hospital Course|10236,10248|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Finding|Body Substance|Hospital Course|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10263,10270|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Occupational Activity|Hospital Course|10289,10293|false|false|false|C0043227|Work|work
Procedure|Diagnostic Procedure|Hospital Course|10289,10296|false|false|false|C0750430|Work-up|work up
Finding|Finding|Hospital Course|10307,10316|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Finding|Functional Concept|Hospital Course|10307,10316|false|false|false|C0220909;C1305399;C1409616|Aspects of disease screening;Screening - procedure intent;Special screening finding|screening
Procedure|Diagnostic Procedure|Hospital Course|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Health Care Activity|Hospital Course|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Research Activity|Hospital Course|10307,10316|false|false|false|C0199230;C0220908;C1698960;C1710031;C1710032|Disease Screening;Screening;Screening for cancer;Screening procedure;research subject screening|screening
Procedure|Diagnostic Procedure|Hospital Course|10318,10329|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Procedure|Health Care Activity|Hospital Course|10318,10329|false|false|false|C0009378;C1548837|Consent Type - Colonoscopy;colonoscopy|colonoscopy
Finding|Finding|Hospital Course|10347,10356|false|false|false|C0260913|Encounter due to Screening for malignant neoplasm of breast|mammogram
Procedure|Diagnostic Procedure|Hospital Course|10347,10356|false|false|false|C0024671|Mammography|mammogram
Finding|Body Substance|Hospital Course|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10359,10366|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10394,10398|false|false|false|C1561540|Transaction counts and value totals - week|week
Finding|Finding|Hospital Course|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Hospital Course|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Hospital Course|10409,10413|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Drug|Pharmacologic Substance|Hospital Course|10420,10423|false|false|false|C0358591|Proton Pump Inhibitors|PPI
Finding|Physiologic Function|Hospital Course|10420,10423|false|false|false|C0871125|Prepulse Inhibition|PPI
Drug|Organic Chemical|Hospital Course|10438,10450|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Pharmacologic Substance|Hospital Course|10438,10450|false|false|false|C0081876|pantoprazole|pantoprazole
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10489,10492|false|false|false|C0082420|Endoglin, human|end
Drug|Immunologic Factor|Hospital Course|10489,10492|false|false|false|C0082420|Endoglin, human|end
Finding|Functional Concept|Hospital Course|10489,10492|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Finding|Gene or Genome|Hospital Course|10489,10492|false|false|false|C1366583;C1561490;C1704837|ENG gene;ENG wt Allele;end - ActRelationshipCheckpoint|end
Procedure|Diagnostic Procedure|Hospital Course|10506,10514|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|Hospital Course|10506,10520|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|Hospital Course|10512,10520|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|10515,10520|false|false|false|C0019080|Hemorrhage|bleed
Finding|Finding|Hospital Course|10521,10527|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|Hospital Course|10521,10527|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Disease or Syndrome|Hospital Course|10534,10543|false|false|false|C0017152|Gastritis|gastritis
Finding|Body Substance|Hospital Course|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10547,10554|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Disorder|Disease or Syndrome|Hospital Course|10557,10569|false|false|false|C0020538|Hypertensive disease|hypertension
Drug|Pharmacologic Substance|Hospital Course|10557,10581|false|false|false|C0684167|hypertensive agents|hypertension medications
Attribute|Clinical Attribute|Hospital Course|10570,10581|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Hospital Course|10570,10581|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Hospital Course|10570,10581|false|false|false|C4284232|Medications|medications
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10583,10593|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|10583,10593|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|10598,10608|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10598,10608|false|false|false|C0028066|nifedipine|nifedipine
Procedure|Diagnostic Procedure|Hospital Course|10628,10636|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|Hospital Course|10628,10642|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|Hospital Course|10634,10642|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|10637,10642|false|false|false|C0019080|Hemorrhage|bleed
Finding|Body Substance|Hospital Course|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10646,10653|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|10656,10666|false|false|false|C0016860|furosemide|furosemide
Drug|Pharmacologic Substance|Hospital Course|10656,10666|false|false|false|C0016860|furosemide|furosemide
Finding|Body Substance|Hospital Course|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10697,10704|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|10707,10717|false|false|false|C0028066|nifedipine|nifedipine
Drug|Pharmacologic Substance|Hospital Course|10707,10717|false|false|false|C0028066|nifedipine|nifedipine
Finding|Intellectual Product|Hospital Course|10752,10757|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Finding|Pathologic Function|Hospital Course|10759,10764|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Space or Junction|Hospital Course|10769,10773|false|false|false|C0228216|Structure of subparietal sulcus|SBPs
Finding|Body Substance|Hospital Course|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|Hospital Course|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|Hospital Course|10787,10794|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Drug|Organic Chemical|Hospital Course|10810,10818|false|false|false|C0699129|Coumadin|Coumadin
Drug|Pharmacologic Substance|Hospital Course|10810,10818|false|false|false|C0699129|Coumadin|Coumadin
Drug|Organic Chemical|Hospital Course|10820,10831|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|10820,10831|false|false|false|C0070166|clopidogrel|Clopidogrel
Anatomy|Body System|Hospital Course|10849,10859|false|false|false|C0007226|Cardiovascular system|cardiology
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Enzyme|Hospital Course|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Organic Chemical|Hospital Course|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Drug|Pharmacologic Substance|Hospital Course|10861,10864|false|false|false|C0004057;C3853627|Arylsulfatase A, human;aspirin|ASA
Finding|Gene or Genome|Hospital Course|10861,10864|false|false|false|C1412553|ARSA gene|ASA
Attribute|Clinical Attribute|Hospital Course|10894,10901|false|false|false|C2741676||address
Finding|Intellectual Product|Hospital Course|10894,10901|false|false|false|C0376649;C1442065;C1547327;C1578436;C1578437;C4319699|Address;Address (property);Address Data Type;Addresses (publication format);MDF Attribute Type - Address;Value type - Address|address
Finding|Body Substance|Hospital Course|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|10902,10909|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|10912,10916|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10912,10916|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10912,10916|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|10912,10928|false|false|false|C2242846|home environment (history)|home environment
Finding|Finding|Hospital Course|10933,10937|false|false|false|C0085639|Falls|fall
Finding|Finding|Hospital Course|10933,10942|false|false|false|C1268740|At increased risk for falls|fall risk
Finding|Idea or Concept|Hospital Course|10938,10942|false|false|false|C0035647|Risk|risk
Drug|Amino Acid, Peptide, or Protein|Hospital Course|10958,10962|false|false|false|C0077275|triptorelin|trip
Drug|Hormone|Hospital Course|10958,10962|false|false|false|C0077275|triptorelin|trip
Drug|Pharmacologic Substance|Hospital Course|10958,10962|false|false|false|C0077275|triptorelin|trip
Finding|Gene or Genome|Hospital Course|10958,10962|false|false|false|C1416921;C2239819;C2608049;C4085339|LRRFIP1 gene;PIK3IP1 gene;TRAIP gene;TRAIP wt Allele|trip
Phenomenon|Phenomenon or Process|Hospital Course|10958,10962|false|false|false|C0221188|Tripping|trip
Finding|Finding|Hospital Course|10964,10971|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Hospital Course|10967,10971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Hospital Course|10967,10971|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Hospital Course|10967,10971|false|false|false|C1553498|home health encounter|home
Finding|Finding|Hospital Course|10976,10979|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Hospital Course|10976,10979|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Finding|Hospital Course|10980,10995|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|10980,10995|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|10980,10995|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Finding|Body Substance|Hospital Course|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Hospital Course|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Hospital Course|11013,11020|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|Hospital Course|11013,11024|false|false|false|C0332310|Has patient|patient has
Finding|Classification|Hospital Course|11025,11035|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Hospital Course|11025,11035|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Finding|Hospital Course|11036,11051|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Finding|Physiologic Function|Hospital Course|11036,11051|false|false|false|C2919015;C3537050;C5887107|ANTICOAGULATION (finding);Anticoagulation function;Decreased Coagulation Activity [PE]|anticoagulation
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11036,11051|false|false|false|C0003281|Anticoagulation Therapy|anticoagulation
Event|Occupational Activity|Hospital Course|11067,11077|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Hospital Course|11067,11077|false|false|false|C0376636|Disease Management|management
Finding|Body Substance|Hospital Course|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|Hospital Course|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|Hospital Course|11083,11092|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|Hospital Course|11083,11092|false|false|false|C0030685|Patient Discharge|discharge
Procedure|Therapeutic or Preventive Procedure|Hospital Course|11098,11103|false|false|false|C0034991|Rehabilitation therapy|rehab
Attribute|Clinical Attribute|Hospital Course|11109,11120|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11109,11120|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|11109,11120|false|false|false|C4284232|Medications|Medications
Finding|Finding|Hospital Course|11109,11133|false|false|false|C1627937|Medications on admission|Medications on Admission
Procedure|Health Care Activity|Hospital Course|11124,11133|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|Hospital Course|11152,11162|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|Hospital Course|11152,11162|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|Hospital Course|11152,11167|false|false|false|C0746470|MEDICATION LIST|Medication list
Finding|Intellectual Product|Hospital Course|11163,11167|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Drug|Organic Chemical|Hospital Course|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|Hospital Course|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|Hospital Course|11184,11192|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Finding|Functional Concept|Hospital Course|11184,11192|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|Hospital Course|11184,11192|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11197,11207|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|11197,11207|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|11227,11238|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|11227,11238|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Organic Chemical|Hospital Course|11259,11271|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11259,11271|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|11289,11299|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|11289,11299|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11311,11314|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11311,11314|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11311,11314|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11311,11314|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11319,11330|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Hospital Course|11319,11330|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Hospital Course|11350,11360|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|11350,11360|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|Hospital Course|11380,11390|false|false|false|C0034665|ranitidine|Ranitidine
Drug|Pharmacologic Substance|Hospital Course|11380,11390|false|false|false|C0034665|ranitidine|Ranitidine
Finding|Gene or Genome|Hospital Course|11407,11410|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Pathologic Function|Hospital Course|11411,11417|false|false|false|C0232483|Reflux|reflux
Drug|Organic Chemical|Hospital Course|11422,11429|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|11422,11429|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|11449,11462|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|11465,11468|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|11483,11490|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|11483,11492|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|11483,11492|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Organic Chemical|Hospital Course|11516,11526|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|11516,11526|false|false|false|C0028066|nifedipine|NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11539,11542|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11539,11542|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11539,11542|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11539,11542|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11548,11561|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|11548,11561|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Hospital Course|11581,11584|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|11585,11590|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|11585,11590|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|11585,11595|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|11585,11595|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|11591,11595|false|true|false|C2598155||pain
Finding|Functional Concept|Hospital Course|11591,11595|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|11591,11595|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Daily or Recreational Activity|Hospital Course|11616,11622|false|false|false|C4048877|Dinner|Dinner
Finding|Body Substance|Hospital Course|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|11626,11635|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|11626,11635|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|11626,11647|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|Hospital Course|11636,11647|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|Hospital Course|11636,11647|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Finding|Intellectual Product|Hospital Course|11636,11647|false|false|false|C4284232|Medications|Medications
Drug|Organic Chemical|Hospital Course|11652,11663|false|false|false|C0002144|allopurinol|Allopurinol
Drug|Pharmacologic Substance|Hospital Course|11652,11663|false|false|false|C0002144|allopurinol|Allopurinol
Finding|Idea or Concept|Hospital Course|11686,11689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Finding|Intellectual Product|Hospital Course|11686,11689|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|DAY
Drug|Organic Chemical|Hospital Course|11694,11701|false|false|false|C0004057|aspirin|Aspirin
Drug|Pharmacologic Substance|Hospital Course|11694,11701|false|false|false|C0004057|aspirin|Aspirin
Drug|Organic Chemical|Hospital Course|11721,11733|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Pharmacologic Substance|Hospital Course|11721,11733|false|false|false|C0286651|atorvastatin|Atorvastatin
Drug|Organic Chemical|Hospital Course|11751,11761|false|false|false|C0054836|carvedilol|Carvedilol
Drug|Pharmacologic Substance|Hospital Course|11751,11761|false|false|false|C0054836|carvedilol|Carvedilol
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11773,11776|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11773,11776|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11773,11776|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11773,11776|false|false|false|C1332410|BID gene|BID
Finding|Daily or Recreational Activity|Hospital Course|11796,11802|false|false|false|C4048877|Dinner|Dinner
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11806,11816|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Pharmacologic Substance|Hospital Course|11806,11816|false|false|false|C0065374|lisinopril|Lisinopril
Drug|Organic Chemical|Hospital Course|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Pharmacologic Substance|Hospital Course|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Vitamin|Hospital Course|11836,11849|false|false|false|C0301532;C3714835|Multivitamin Drug Class;Multivitamin preparation|Multivitamins
Drug|Biomedical or Dental Material|Hospital Course|11852,11855|false|false|false|C0039225|Tablet Dosage Form|TAB
Drug|Organic Chemical|Hospital Course|11869,11879|false|false|false|C0028066|nifedipine|NIFEdipine
Drug|Pharmacologic Substance|Hospital Course|11869,11879|false|false|false|C0028066|nifedipine|NIFEdipine
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11892,11895|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11892,11895|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11892,11895|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11892,11895|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Pharmacologic Substance|Hospital Course|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Vitamin|Hospital Course|11900,11907|false|false|false|C0042890|Vitamins|Vitamin
Drug|Hormone|Hospital Course|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Organic Chemical|Hospital Course|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Pharmacologic Substance|Hospital Course|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Drug|Vitamin|Hospital Course|11900,11909|false|false|false|C0014695;C0042866;C2936842;C3537249;C3714503|D Vitamin;Vitamin D Drug Class;Vitamin D [EPC];ergocalciferol;vitamin D|Vitamin D
Procedure|Laboratory Procedure|Hospital Course|11900,11909|false|false|false|C0919758|Vitamin D measurement|Vitamin D
Drug|Organic Chemical|Hospital Course|11933,11941|false|false|false|C1692318|docusate|Docusate
Drug|Pharmacologic Substance|Hospital Course|11933,11941|false|false|false|C1692318|docusate|Docusate
Drug|Organic Chemical|Hospital Course|11933,11948|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Pharmacologic Substance|Hospital Course|11933,11948|false|false|false|C0243237|docusate sodium|Docusate Sodium
Drug|Biologically Active Substance|Hospital Course|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Element, Ion, or Isotope|Hospital Course|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Drug|Pharmacologic Substance|Hospital Course|11942,11948|false|false|false|C0037473;C3541959;C3714642|Sodium Drug Class;Sodium supplements;sodium|Sodium
Finding|Physiologic Function|Hospital Course|11942,11948|false|false|false|C4553025|Sodium metabolic function|Sodium
Procedure|Laboratory Procedure|Hospital Course|11942,11948|false|false|false|C0337443|Sodium measurement|Sodium
Disorder|Mental or Behavioral Dysfunction|Hospital Course|11959,11962|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|11959,11962|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|11959,11962|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|11959,11962|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|Hospital Course|11968,11978|false|false|false|C0060926|gabapentin|Gabapentin
Drug|Pharmacologic Substance|Hospital Course|11968,11978|false|false|false|C0060926|gabapentin|Gabapentin
Finding|Finding|Hospital Course|11993,12009|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Finding|Sign or Symptom|Hospital Course|11993,12009|false|false|false|C0027796;C3714625|Neuralgia;Neuropathic pain|neuropathic pain
Attribute|Clinical Attribute|Hospital Course|12005,12009|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|12005,12009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12005,12009|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12015,12027|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Hospital Course|12015,12027|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Organic Chemical|Hospital Course|12047,12052|false|false|false|C3489575|sennosides, USP|Senna
Drug|Pharmacologic Substance|Hospital Course|12047,12052|false|false|false|C3489575|sennosides, USP|Senna
Disorder|Mental or Behavioral Dysfunction|Hospital Course|12063,12066|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|Hospital Course|12063,12066|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|Hospital Course|12063,12066|false|false|false|C1530795|BID protein, human|BID
Finding|Gene or Genome|Hospital Course|12063,12066|false|false|false|C1332410|BID gene|BID
Finding|Sign or Symptom|Hospital Course|12067,12079|false|false|false|C0009806|Constipation|constipation
Drug|Hazardous or Poisonous Substance|Hospital Course|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Drug|Organic Chemical|Hospital Course|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Drug|Pharmacologic Substance|Hospital Course|12085,12093|false|false|false|C0043031|warfarin|Warfarin
Attribute|Clinical Attribute|Hospital Course|12138,12141|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Procedure|Laboratory Procedure|Hospital Course|12138,12141|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12138,12141|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Drug|Organic Chemical|Hospital Course|12147,12160|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Drug|Pharmacologic Substance|Hospital Course|12147,12160|false|false|false|C0017887|nitroglycerin|Nitroglycerin
Finding|Gene or Genome|Hospital Course|12180,12183|false|false|false|C1422467|CIAO3 gene|PRN
Anatomy|Body Location or Region|Hospital Course|12184,12189|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|Hospital Course|12184,12189|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|Hospital Course|12184,12194|false|false|false|C2926613||chest pain
Finding|Sign or Symptom|Hospital Course|12184,12194|false|false|false|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|Hospital Course|12190,12194|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|12190,12194|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12190,12194|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|Hospital Course|12200,12210|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|Hospital Course|12200,12210|false|false|false|C0016860|furosemide|Furosemide
Drug|Biomedical or Dental Material|Hospital Course|12231,12243|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|12231,12243|false|false|false|C0032487;C0137914;C0752345|Polyethylene;high-density polyethylene;polyethylenes|Polyethylene
Drug|Organic Chemical|Hospital Course|12231,12250|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Pharmacologic Substance|Hospital Course|12231,12250|false|false|false|C0032483|polyethylene glycols|Polyethylene Glycol
Drug|Hazardous or Poisonous Substance|Hospital Course|12244,12250|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|12244,12250|false|false|false|C0015083;C0017945;C0017951|Glycol;Glycols;ethylene glycol|Glycol
Drug|Organic Chemical|Hospital Course|12270,12283|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Drug|Pharmacologic Substance|Hospital Course|12270,12283|false|false|false|C0000970;C2917659|Acetaminophen [EPC];acetaminophen|Acetaminophen
Procedure|Laboratory Procedure|Hospital Course|12270,12283|false|false|false|C0373527|Acetaminophen measurement|Acetaminophen
Finding|Gene or Genome|Hospital Course|12302,12305|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|Hospital Course|12306,12310|false|false|false|C2598155||pain
Finding|Functional Concept|Hospital Course|12306,12310|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Hospital Course|12306,12310|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Finding|Hospital Course|12314,12319|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|Hospital Course|12314,12319|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Body Substance|Hospital Course|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12324,12333|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12324,12333|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|Hospital Course|12324,12345|false|false|false|C4019243||Discharge Disposition
Finding|Finding|Hospital Course|12324,12345|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|Hospital Course|12334,12345|false|false|false|C2926604||Disposition
Procedure|Health Care Activity|Hospital Course|12334,12345|false|false|false|C0184758|Patient disposition|Disposition
Finding|Finding|Hospital Course|12347,12355|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Finding|Functional Concept|Hospital Course|12347,12355|false|false|false|C0231448;C5781021|Extended (finding);Extension|Extended
Procedure|Health Care Activity|Hospital Course|12347,12360|false|false|false|C0023977|long-term care|Extended Care
Event|Activity|Hospital Course|12356,12360|false|false|false|C1947933|care activity|Care
Finding|Finding|Hospital Course|12356,12360|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|12356,12360|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Hospital Course|12363,12371|false|false|false|C4695111|ADMIN.FACILITY|Facility
Finding|Body Substance|Hospital Course|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|Hospital Course|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|Hospital Course|12379,12388|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|Hospital Course|12379,12388|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|Hospital Course|12379,12398|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|Hospital Course|12389,12398|false|false|false|C0945731||Diagnosis
Finding|Classification|Hospital Course|12389,12398|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|Hospital Course|12389,12398|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|Hospital Course|12389,12398|false|false|false|C0011900|Diagnosis|Diagnosis
Attribute|Clinical Attribute|Hospital Course|12409,12413|false|false|false|C4318566|Deep Resection Margin|Deep
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12409,12418|false|false|false|C0226514|Structure of deep vein|Deep vein
Disorder|Disease or Syndrome|Hospital Course|12409,12429|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|Deep vein thrombosis
Disorder|Disease or Syndrome|Hospital Course|12409,12435|false|false|false|C0149871|Deep Vein Thrombosis|Deep vein thrombosis (DVT)
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12414,12418|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Hospital Course|12414,12429|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|Hospital Course|12419,12429|false|false|false|C0040053|Thrombosis|thrombosis
Anatomy|Body Location or Region|Hospital Course|12431,12434|false|false|false|C5239664|area DVT|DVT
Attribute|Clinical Attribute|Hospital Course|12431,12434|false|false|false|C2926618||DVT
Disorder|Disease or Syndrome|Hospital Course|12431,12434|false|false|false|C0149871;C0151950|Deep Vein Thrombosis;Deep thrombophlebitis|DVT
Disorder|Neoplastic Process|Hospital Course|12437,12446|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Finding|Functional Concept|Hospital Course|12437,12446|false|false|false|C1522484|metastatic qualifier|Secondary
Procedure|Diagnostic Procedure|Hospital Course|12448,12456|false|false|false|C0203057|Upper gastrointestinal tract series|Upper GI
Finding|Pathologic Function|Hospital Course|12448,12462|false|false|false|C0041909|Upper gastrointestinal hemorrhage|Upper GI bleed
Finding|Pathologic Function|Hospital Course|12454,12462|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Hospital Course|12457,12462|false|false|false|C0019080|Hemorrhage|bleed
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12463,12468|false|false|false|C5779993|Left arm|L arm
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12465,12468|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Hospital Course|12465,12468|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Hospital Course|12465,12468|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Hospital Course|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Hospital Course|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12465,12468|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Pathologic Function|Hospital Course|12469,12477|false|false|false|C0018944|Hematoma|hematoma
Disorder|Disease or Syndrome|Hospital Course|12478,12506|false|false|false|C1510431|Superficial Thrombophlebitis|Superficial thrombophlebitis
Finding|Pathologic Function|Hospital Course|12490,12506|false|false|false|C0040046|Thrombophlebitis|thrombophlebitis
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12510,12521|false|false|false|C1549091|Antecubital|antecubital
Anatomy|Body Space or Junction|Hospital Course|12510,12527|false|false|false|C0446523|Antecubital Fossa|antecubital fossa
Anatomy|Body Space or Junction|Hospital Course|12522,12527|false|false|false|C0836913|Fossa|fossa
Finding|Intellectual Product|Hospital Course|12528,12535|false|false|false|C1547296|Chronic - Admission Level of Care Code|Chronic
Procedure|Health Care Activity|Hospital Course|12528,12535|false|false|false|C1555457|Provision of recurring care for chronic illness|Chronic
Disorder|Disease or Syndrome|Hospital Course|12528,12550|false|false|false|C1561643|Chronic Kidney Diseases|Chronic kidney disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12536,12542|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Hospital Course|12536,12542|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Finding|Sign or Symptom|Hospital Course|12536,12542|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Hospital Course|12536,12542|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Hospital Course|12536,12542|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Disease or Syndrome|Hospital Course|12536,12550|false|false|false|C0022658|Kidney Diseases|kidney disease
Disorder|Disease or Syndrome|Hospital Course|12543,12550|false|false|false|C0012634|Disease|disease
Attribute|Clinical Attribute|Hospital Course|12552,12557|false|true|false|C1300072|Tumor stage|Stage
Disorder|Disease or Syndrome|Hospital Course|12562,12589|false|false|false|C0085096|Peripheral Vascular Diseases|Peripheral vascular disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12573,12581|false|false|false|C0005847|Blood Vessel|vascular
Disorder|Disease or Syndrome|Hospital Course|12573,12589|false|false|false|C0042373|Vascular Diseases|vascular disease
Disorder|Disease or Syndrome|Hospital Course|12582,12589|false|false|false|C0012634|Disease|disease
Disorder|Disease or Syndrome|Hospital Course|12590,12598|false|false|false|C0011847;C0011849;C0011860|Diabetes;Diabetes Mellitus;Diabetes Mellitus, Non-Insulin-Dependent|Diabetes
Disorder|Disease or Syndrome|Hospital Course|12590,12607|false|false|false|C0011849|Diabetes Mellitus|Diabetes mellitus
Disorder|Disease or Syndrome|Hospital Course|12590,12615|false|false|false|C0011860|Diabetes Mellitus, Non-Insulin-Dependent|Diabetes mellitus type II
Finding|Gene or Genome|Hospital Course|12608,12612|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Finding|Intellectual Product|Hospital Course|12608,12612|false|false|false|C1420009;C1552651|SGCG gene;Type - ParameterizedDataType|type
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12616,12624|false|false|false|C0018787|Heart|Coronary
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12616,12631|false|false|false|C0205042|Coronary artery|Coronary artery
Disorder|Disease or Syndrome|Hospital Course|12616,12639|false|false|false|C0010054;C1956346|Coronary Arteriosclerosis;Coronary Artery Disease|Coronary artery disease
Anatomy|Body Part, Organ, or Organ Component|Hospital Course|12625,12631|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Anatomy|Body System|Hospital Course|12625,12631|false|false|false|C0003842;C0226004|Arterial system;Arteries|artery
Disorder|Disease or Syndrome|Hospital Course|12625,12639|false|false|false|C0852949|Arteriopathic disease|artery disease
Disorder|Disease or Syndrome|Hospital Course|12632,12639|false|false|false|C0012634|Disease|disease
Finding|Mental Process|Discharge Condition|12664,12670|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|12664,12677|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|12664,12677|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|12671,12677|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|12671,12677|false|false|false|C1546481|What subject filter - Status|Status
Finding|Idea or Concept|Discharge Condition|12679,12684|false|false|false|C1550016|Remote control command - Clear|Clear
Finding|Finding|Discharge Condition|12689,12697|false|false|false|C4068804|Coherent|coherent
Attribute|Clinical Attribute|Discharge Condition|12699,12721|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|12699,12721|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Finding|Finding|Discharge Condition|12708,12721|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|12708,12721|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|12723,12728|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|12723,12728|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|12723,12728|false|false|false|C0718338|Alert brand of caffeine|Alert
Finding|Finding|Discharge Condition|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|12723,12728|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|12733,12744|false|false|false|C1704675|Interaction|interactive
Finding|Gene or Genome|Discharge Instructions|12773,12777|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Finding|Intellectual Product|Discharge Instructions|12793,12801|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|12793,12801|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12848,12851|false|false|false|C0023216;C1140621|Leg;Lower Extremity|leg
Finding|Pathologic Function|Discharge Instructions|12848,12860|false|true|false|C0581394|Swelling of lower limb|leg swelling
Finding|Finding|Discharge Instructions|12852,12860|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|Discharge Instructions|12852,12860|false|false|false|C0013604;C0038999|Edema;Swelling|swelling
Attribute|Clinical Attribute|Discharge Instructions|12865,12869|false|false|false|C2598155||pain
Finding|Functional Concept|Discharge Instructions|12865,12869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|Discharge Instructions|12865,12869|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Indicator, Reagent, or Diagnostic Aid|Discharge Instructions|12871,12881|false|false|false|C0358514|Diagnostic agents|Diagnostic
Finding|Functional Concept|Discharge Instructions|12871,12881|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Finding|Intellectual Product|Discharge Instructions|12871,12881|false|false|false|C0348026;C1547424|Diagnostic;Location Service Code - Diagnostic|Diagnostic
Procedure|Diagnostic Procedure|Discharge Instructions|12871,12881|false|false|false|C0011900;C0430533|Diagnosis;Diagnostic dental procedure|Diagnostic
Procedure|Diagnostic Procedure|Discharge Instructions|12871,12887|false|false|false|C0086143|Diagnostic tests|Diagnostic tests
Finding|Intellectual Product|Discharge Instructions|12882,12887|false|false|false|C0392366|Tests (qualifier value)|tests
Procedure|Laboratory Procedure|Discharge Instructions|12882,12887|false|false|false|C0022885|Laboratory Procedures|tests
Attribute|Clinical Attribute|Discharge Instructions|12932,12936|false|false|false|C4318566|Deep Resection Margin|deep
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12932,12941|false|false|false|C0226514|Structure of deep vein|deep vein
Disorder|Disease or Syndrome|Discharge Instructions|12932,12952|false|false|false|C0149871;C0340708|Deep Vein Thrombosis;Deep vein thrombosis of lower limb|deep vein thrombosis
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12937,12941|false|false|false|C0042449|Veins|vein
Finding|Pathologic Function|Discharge Instructions|12937,12952|false|false|false|C0042487|Venous Thrombosis|vein thrombosis
Finding|Pathologic Function|Discharge Instructions|12942,12952|false|false|false|C0040053|Thrombosis|thrombosis
Disorder|Disease or Syndrome|Discharge Instructions|12954,12959|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|12954,12959|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|Discharge Instructions|12954,12965|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clots
Finding|Pathologic Function|Discharge Instructions|12960,12965|false|false|false|C0302148|Blood Clot|clots
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|12975,12979|false|false|false|C1140621|Leg|legs
Attribute|Clinical Attribute|Discharge Instructions|12975,12979|false|false|false|C5781420||legs
Disorder|Disease or Syndrome|Discharge Instructions|13003,13008|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|13003,13008|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Sign or Symptom|Discharge Instructions|13009,13017|false|false|false|C0851184|Thinning Weight Loss|thinning
Attribute|Clinical Attribute|Discharge Instructions|13018,13029|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|Discharge Instructions|13018,13029|false|false|false|C0013227|Pharmaceutical Preparations|medications
Finding|Intellectual Product|Discharge Instructions|13018,13029|false|false|false|C4284232|Medications|medications
Finding|Finding|Discharge Instructions|13054,13061|false|false|false|C4534363|At home|at home
Finding|Idea or Concept|Discharge Instructions|13057,13061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|Discharge Instructions|13057,13061|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|Discharge Instructions|13057,13061|false|false|false|C1553498|home health encounter|home
Procedure|Diagnostic Procedure|Discharge Instructions|13085,13093|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|Discharge Instructions|13085,13102|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleeding
Finding|Pathologic Function|Discharge Instructions|13091,13102|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleeding
Finding|Pathologic Function|Discharge Instructions|13094,13102|false|false|false|C0019080|Hemorrhage|bleeding
Drug|Pharmacologic Substance|Discharge Instructions|13158,13168|false|false|false|C0013227|Pharmaceutical Preparations|medication
Finding|Intellectual Product|Discharge Instructions|13158,13168|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|medication
Procedure|Diagnostic Procedure|Discharge Instructions|13191,13194|false|false|false|C0079304|Esophagogastroduodenoscopy|EGD
Finding|Functional Concept|Discharge Instructions|13212,13216|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13212,13220|false|false|false|C0230347;C5779993|Left arm;Left upper arm structure|left arm
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|13217,13220|false|false|false|C0446516;C1140618;C1269078|Upper Extremity;Upper arm|arm
Disorder|Anatomical Abnormality|Discharge Instructions|13217,13220|false|false|false|C3495676|Anorectal Malformations|arm
Finding|Gene or Genome|Discharge Instructions|13217,13220|false|false|false|C1824218;C3715044|AKR1A1 wt Allele;ARMC9 gene|arm
Procedure|Diagnostic Procedure|Discharge Instructions|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Research Activity|Discharge Instructions|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|13217,13220|false|false|false|C1522541;C4761640;C5400986|Axillary Reverse Mapping;Protocol Treatment Arm;Study Arm|arm
Finding|Pathologic Function|Discharge Instructions|13221,13229|false|false|false|C0018944|Hematoma|hematoma
Finding|Finding|Discharge Instructions|13234,13238|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|Discharge Instructions|13282,13285|false|false|false|C5939094|Own|own
Finding|Finding|Discharge Instructions|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Idea or Concept|Discharge Instructions|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Finding|Intellectual Product|Discharge Instructions|13291,13295|false|false|false|C1547403;C1548318;C2024467;C3541383;C5400024;C5575590|Data types - Time;Instructions for Use of the CPT Codebook - Time;Time (foundation metadata concept);Time - Instructions for Selecting a Level of Pathology Clinical Consultation Services;Value type - Time|time
Disorder|Disease or Syndrome|Discharge Instructions|13307,13312|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|13307,13312|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Pathologic Function|Discharge Instructions|13307,13318|false|false|false|C0087086;C0302148|Blood Clot;Thrombus|blood clots
Finding|Pathologic Function|Discharge Instructions|13313,13318|false|false|false|C0302148|Blood Clot|clots
Finding|Finding|Discharge Instructions|13342,13345|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Finding|Idea or Concept|Discharge Instructions|13342,13345|false|false|false|C1553390;C1578513|Act Status - new;Query Status Code - new|new
Drug|Pharmacologic Substance|Discharge Instructions|13346,13350|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Discharge Instructions|13346,13350|false|false|false|C0740721|Drug problem|drug
Drug|Hazardous or Poisonous Substance|Discharge Instructions|13359,13367|false|false|false|C0043031|warfarin|warfarin
Drug|Organic Chemical|Discharge Instructions|13359,13367|false|false|false|C0043031|warfarin|warfarin
Drug|Pharmacologic Substance|Discharge Instructions|13359,13367|false|false|false|C0043031|warfarin|warfarin
Disorder|Disease or Syndrome|Discharge Instructions|13396,13401|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Finding|Body Substance|Discharge Instructions|13396,13401|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Procedure|Diagnostic Procedure|Discharge Instructions|13442,13450|false|false|false|C0203057|Upper gastrointestinal tract series|upper GI
Finding|Pathologic Function|Discharge Instructions|13442,13456|false|false|false|C0041909|Upper gastrointestinal hemorrhage|upper GI bleed
Finding|Pathologic Function|Discharge Instructions|13448,13456|false|false|false|C0017181|Gastrointestinal Hemorrhage|GI bleed
Finding|Pathologic Function|Discharge Instructions|13451,13456|false|false|false|C0019080|Hemorrhage|bleed
Drug|Organic Chemical|Discharge Instructions|13479,13491|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Discharge Instructions|13479,13491|false|false|false|C0081876|pantoprazole|Pantoprazole
Drug|Pharmacologic Substance|Discharge Instructions|13533,13537|false|false|false|C0013227;C1254351|Pharmaceutical Preparations;Pharmacologic Substance|drug
Finding|Finding|Discharge Instructions|13533,13537|false|false|false|C0740721|Drug problem|drug
Finding|Classification|Discharge Instructions|13545,13555|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|Discharge Instructions|13545,13555|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|Discharge Instructions|13622,13633|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Pharmacologic Substance|Discharge Instructions|13622,13633|false|false|false|C0070166|clopidogrel|Clopidogrel
Drug|Organic Chemical|Discharge Instructions|13635,13641|false|false|false|C0633084|Plavix|Plavix
Drug|Pharmacologic Substance|Discharge Instructions|13635,13641|false|false|false|C0633084|Plavix|Plavix
Finding|Intellectual Product|Discharge Instructions|13695,13703|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|13695,13703|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|13711,13715|false|false|false|C1947933|care activity|care
Finding|Finding|Discharge Instructions|13711,13715|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|13711,13715|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Idea or Concept|Discharge Instructions|13732,13740|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Activity|Discharge Instructions|13771,13775|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|13771,13775|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|13771,13775|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|13771,13780|false|false|false|C4321316||Care Team
Finding|Finding|Discharge Instructions|13771,13780|false|false|false|C4321315|Care team|Care Team
Procedure|Health Care Activity|Discharge Instructions|13783,13791|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|13792,13804|false|false|false|C3263700||Instructions
Finding|Intellectual Product|Discharge Instructions|13792,13804|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

