 Semantic Group | Semantic Type | Section | Span | Negated | Uncertain | Generic | CUI | Preferred Text | Document Text 
Event|Event|SIMPLE_SEGMENT|2,6|false|false|false|||Name
Finding|Intellectual Product|SIMPLE_SEGMENT|2,6|false|false|false|C0027365;C1547383;C1554107|MDF Attribute Type - Name;Name;Person Name|Name
Event|Event|SIMPLE_SEGMENT|50,59|false|false|false|||Admission
Procedure|Health Care Activity|SIMPLE_SEGMENT|50,59|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Attribute|Clinical Attribute|SIMPLE_SEGMENT|50,64|false|false|false|C2598112||Admission Date
Event|Event|SIMPLE_SEGMENT|84,93|false|false|false|||Discharge
Finding|Body Substance|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|SIMPLE_SEGMENT|84,93|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|SIMPLE_SEGMENT|84,93|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|SIMPLE_SEGMENT|84,98|false|false|false|C2361122||Discharge Date
Finding|Finding|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Intellectual Product|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Finding|Organism Function|SIMPLE_SEGMENT|116,121|false|false|false|C0005615;C1148523;C1550722;C3245487;C4551887|Birth;Childbirth;Entity Name Part Qualifier - birth;Name Given at Birth;birth (history)|Birth
Attribute|Clinical Attribute|SIMPLE_SEGMENT|140,143|false|false|false|C0804628||Sex
Finding|Behavior|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Finding|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Gene or Genome|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Finding|Organism Function|SIMPLE_SEGMENT|140,143|false|false|false|C0009253;C0036864;C1314687;C1418662|Coitus;PLXNA3 gene;Sex Behavior|Sex
Event|Occupational Activity|SIMPLE_SEGMENT|151,158|false|false|false|C0557854|Services|Service
Finding|Idea or Concept|SIMPLE_SEGMENT|151,158|false|false|false|C3245478|ActInformationPrivacyReason - service|Service
Drug|Pharmacologic Substance|SIMPLE_SEGMENT|160,168|false|false|false|C0013227|Pharmaceutical Preparations|MEDICINE
Drug|Organic Chemical|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Drug|Pharmacologic Substance|Allergies|183,191|false|false|false|C0086787|Percocet|Percocet
Drug|Organic Chemical|Allergies|194,201|false|false|false|C0483514|Vicodin|Vicodin
Drug|Pharmacologic Substance|Allergies|194,201|false|false|false|C0483514|Vicodin|Vicodin
Event|Event|Allergies|204,213|false|false|false|||Attending
Finding|Functional Concept|Allergies|204,213|false|false|false|C1999232|Attending (action)|Attending
Event|Event|Chief Complaint|238,245|false|false|false|||altered
Finding|Mental Process|Chief Complaint|246,252|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|Chief Complaint|246,259|false|false|false|C0488568;C0488569||mental status
Finding|Finding|Chief Complaint|246,259|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|Chief Complaint|253,259|false|false|false|C5889824||status
Event|Event|Chief Complaint|253,259|false|false|false|||status
Finding|Idea or Concept|Chief Complaint|253,259|false|false|false|C1546481|What subject filter - Status|status
Finding|Classification|Chief Complaint|262,267|false|false|false|C4521762|United States Military Commissioned Officer O4 (qualifier value)|Major
Procedure|Health Care Activity|Chief Complaint|268,276|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|268,276|false|false|false|C0543467;C0587668|Operative Surgical Procedures;Surgical service|Surgical
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|280,298|false|false|false|C4048276|Invasive procedure|Invasive Procedure
Attribute|Clinical Attribute|Chief Complaint|289,298|false|false|false|C0945766||Procedure
Event|Event|Chief Complaint|289,298|false|false|false|||Procedure
Event|Occupational Activity|Chief Complaint|289,298|false|false|false|C1546467|Act Class - procedure|Procedure
Finding|Functional Concept|Chief Complaint|289,298|false|false|false|C2700391|Procedure (set of actions)|Procedure
Procedure|Therapeutic or Preventive Procedure|Chief Complaint|289,298|false|false|false|C0184661|Interventional procedure|Procedure
Disorder|Disease or Syndrome|History of Present Illness|365,368|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|History of Present Illness|365,368|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|History of Present Illness|365,368|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|History of Present Illness|365,368|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|History of Present Illness|365,368|false|false|false|||HIV
Event|Event|History of Present Illness|372,377|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|372,377|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|History of Present Illness|379,383|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|History of Present Illness|379,383|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|History of Present Illness|379,383|false|false|false|||COPD
Finding|Gene or Genome|History of Present Illness|379,383|false|false|false|C1412502|ARCN1 gene|COPD
Disorder|Disease or Syndrome|History of Present Illness|385,388|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|History of Present Illness|385,388|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|History of Present Illness|385,388|false|false|false|||HCV
Disorder|Disease or Syndrome|History of Present Illness|390,399|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|History of Present Illness|390,399|false|false|false|||cirrhosis
Event|Event|History of Present Illness|400,411|false|false|false|||complicated
Disorder|Disease or Syndrome|History of Present Illness|415,422|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|415,422|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|415,422|false|false|false|C5441966|Peritoneal Effusion|ascites
Anatomy|Body Location or Region|History of Present Illness|427,434|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|History of Present Illness|427,449|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|History of Present Illness|435,449|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|History of Present Illness|435,449|false|false|false|||encephalopathy
Event|Event|History of Present Illness|465,474|false|false|false|||presented
Event|Event|History of Present Illness|500,511|false|false|false|||hypotension
Finding|Finding|History of Present Illness|500,511|false|false|false|C0020649|Hypotension|hypotension
Event|Event|History of Present Illness|521,533|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|521,533|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Body Substance|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|541,548|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|History of Present Illness|541,552|false|false|false|C0332310|Has patient|patient has
Event|Event|History of Present Illness|557,568|false|false|false|||accelerated
Event|Event|History of Present Illness|569,583|false|false|false|||decompensation
Finding|Finding|History of Present Illness|569,583|false|false|false|C0231187|Decompensation|decompensation
Disorder|Disease or Syndrome|History of Present Illness|591,600|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|History of Present Illness|591,600|false|false|false|||cirrhosis
Finding|Idea or Concept|History of Present Illness|616,625|false|false|false|C1546960|Patient Outcome - Worsening|worsening
Disorder|Disease or Syndrome|History of Present Illness|626,633|false|false|false|C0003962|Ascites|ascites
Event|Event|History of Present Illness|626,633|false|false|false|||ascites
Finding|Pathologic Function|History of Present Illness|626,633|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|History of Present Illness|646,656|false|false|false|||maintained
Event|Event|History of Present Illness|674,686|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|674,686|false|false|false|C0034115|Paracentesis|paracentesis
Event|Event|History of Present Illness|711,718|false|false|false|C1883016|Activity Session|session
Finding|Conceptual Entity|History of Present Illness|711,718|false|false|false|C1883017|Session|session
Event|Event|History of Present Illness|719,728|false|false|false|||yesterday
Event|Event|History of Present Illness|743,754|false|false|false|||hypotension
Finding|Finding|History of Present Illness|743,754|false|false|false|C0020649|Hypotension|hypotension
Attribute|Clinical Attribute|History of Present Illness|758,761|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|758,761|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|History of Present Illness|758,761|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|History of Present Illness|758,761|false|false|false|||SBP
Finding|Gene or Genome|History of Present Illness|758,761|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|History of Present Illness|758,761|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|History of Present Illness|775,790|false|false|false|||lightheadedness
Finding|Sign or Symptom|History of Present Illness|775,790|false|false|false|C0220870|Lightheadedness|lightheadedness
Finding|Body Substance|History of Present Illness|801,808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|801,808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|801,808|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|826,832|false|false|false|||memory
Finding|Finding|History of Present Illness|826,832|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Intellectual Product|History of Present Illness|826,832|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Finding|Mental Process|History of Present Illness|826,832|false|false|false|C0025260;C0700327;C4282129|Memory;Memory G-code;Memory observations|memory
Event|Event|History of Present Illness|833,840|false|false|false|||started
Event|Event|History of Present Illness|848,853|false|false|false|||fuzzy
Finding|Finding|History of Present Illness|848,853|false|false|false|C0541974|Fuzzy head|fuzzy
Finding|Finding|History of Present Illness|874,878|true|true|false|C4281574|Much|much
Event|Event|History of Present Illness|879,891|true|false|false|||recollection
Event|Event|History of Present Illness|900,908|false|false|false|||happened
Finding|Intellectual Product|History of Present Illness|915,919|false|false|false|C1720594|Then - dosing instruction fragment|then
Finding|Classification|History of Present Illness|926,936|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|History of Present Illness|926,936|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|History of Present Illness|937,949|false|false|false|||hepatologist
Event|Event|History of Present Illness|950,953|false|false|false|||saw
Event|Event|History of Present Illness|962,973|false|false|false|||recommended
Event|Event|History of Present Illness|983,985|false|false|false|||go
Event|Event|History of Present Illness|1017,1026|false|false|false|||evaluated
Event|Event|History of Present Illness|1031,1037|false|false|false|||deemed
Event|Event|History of Present Illness|1047,1053|false|false|false|||stable
Finding|Intellectual Product|History of Present Illness|1047,1053|false|false|false|C1547311|Patient Condition Code - Stable|stable
Finding|Finding|History of Present Illness|1047,1068|false|false|false|C0428896|Stable blood pressure|stable blood pressure
Disorder|Disease or Syndrome|History of Present Illness|1054,1059|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|History of Present Illness|1054,1059|false|false|false|||blood
Finding|Body Substance|History of Present Illness|1054,1059|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|History of Present Illness|1054,1068|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|History of Present Illness|1054,1068|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|History of Present Illness|1054,1068|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|History of Present Illness|1060,1068|false|false|false|||pressure
Finding|Finding|History of Present Illness|1060,1068|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|History of Present Illness|1060,1068|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|History of Present Illness|1060,1068|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|History of Present Illness|1060,1068|false|false|false|C0033095||pressure
Event|Event|History of Present Illness|1078,1088|false|false|false|||discharged
Event|Event|History of Present Illness|1089,1093|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1089,1093|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1089,1093|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1089,1093|false|false|false|C1553498|home health encounter|home
Finding|Finding|History of Present Illness|1095,1102|false|false|false|C4534363|At home|At home
Event|Event|History of Present Illness|1098,1102|false|false|false|||home
Finding|Idea or Concept|History of Present Illness|1098,1102|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|History of Present Illness|1098,1102|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|History of Present Illness|1098,1102|false|false|false|C1553498|home health encounter|home
Event|Event|History of Present Illness|1113,1122|false|false|false|||worsening
Finding|Mental Process|History of Present Illness|1123,1129|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|History of Present Illness|1123,1136|false|false|false|C0488568;C0488569||mental status
Finding|Finding|History of Present Illness|1123,1136|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|History of Present Illness|1130,1136|false|false|false|C5889824||status
Event|Event|History of Present Illness|1130,1136|false|false|false|||status
Finding|Idea or Concept|History of Present Illness|1130,1136|false|false|false|C1546481|What subject filter - Status|status
Event|Event|History of Present Illness|1163,1172|false|false|false|||concerned
Event|Event|History of Present Illness|1183,1191|false|false|false|||returned
Finding|Idea or Concept|History of Present Illness|1216,1223|false|false|false|C1555582|Initial (abbreviation)|initial
Event|Event|History of Present Illness|1224,1230|false|false|false|||vitals
Finding|Body Substance|History of Present Illness|1266,1273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1266,1273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1266,1273|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|History of Present Illness|1283,1291|false|false|false|||oriented
Attribute|Clinical Attribute|History of Present Illness|1295,1301|false|false|false|C5890614||person
Event|Event|History of Present Illness|1295,1301|false|false|false|||person
Finding|Intellectual Product|History of Present Illness|1295,1301|false|false|false|C1522390|Person Info|person
Lab|Laboratory or Test Result|History of Present Illness|1307,1311|false|false|false|C0587081|Laboratory test finding|labs
Event|Event|History of Present Illness|1317,1324|false|false|false|||notable
Drug|Biomedical or Dental Material|History of Present Illness|1353,1361|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|History of Present Illness|1353,1361|false|false|false|||baseline
Finding|Idea or Concept|History of Present Illness|1353,1361|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Disorder|Neoplastic Process|History of Present Illness|1368,1371|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1368,1371|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|History of Present Illness|1368,1371|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|History of Present Illness|1368,1371|false|false|false|||ALT
Finding|Gene or Genome|History of Present Illness|1368,1371|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|History of Present Illness|1368,1371|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|History of Present Illness|1368,1371|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1368,1371|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|History of Present Illness|1377,1380|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|History of Present Illness|1377,1380|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|History of Present Illness|1377,1380|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|History of Present Illness|1377,1380|false|false|false|||AST
Finding|Gene or Genome|History of Present Illness|1377,1380|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1398,1401|false|false|false|C0023759|Lip structure|Lip
Disorder|Disease or Syndrome|History of Present Illness|1398,1401|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|Lip
Disorder|Neoplastic Process|History of Present Illness|1398,1401|false|false|false|C0153932;C0264511|Benign neoplasm of the lip;Lymphoid interstitial pneumonia|Lip
Finding|Gene or Genome|History of Present Illness|1398,1401|false|false|false|C1846919;C3889123|SMG1 gene;SMG1 wt Allele|Lip
Attribute|Clinical Attribute|History of Present Illness|1406,1409|false|false|false|C0368980|Coagulation tissue factor induced.INR|INR
Event|Event|History of Present Illness|1406,1409|false|false|false|||INR
Procedure|Laboratory Procedure|History of Present Illness|1406,1409|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1406,1409|false|false|false|C0525032;C1704538|Integrated Neuromusculoskeletal Release;International Normalized Ratio|INR
Finding|Idea or Concept|History of Present Illness|1415,1422|false|false|false|C1555582|Initial (abbreviation)|Initial
Event|Event|History of Present Illness|1423,1426|false|false|false|||EKG
Finding|Intellectual Product|History of Present Illness|1423,1426|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|History of Present Illness|1423,1426|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|History of Present Illness|1427,1433|false|false|false|||showed
Anatomy|Body Space or Junction|History of Present Illness|1434,1439|false|false|false|C0030471;C1305231|Nasal sinus;Sinus - general anatomical term|sinus
Disorder|Anatomical Abnormality|History of Present Illness|1434,1439|false|false|false|C0016169|pathologic fistula|sinus
Drug|Organic Chemical|History of Present Illness|1434,1439|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Drug|Pharmacologic Substance|History of Present Illness|1434,1439|false|false|false|C0723346|Sinus brand of acetaminophen-pseudoephedrine|sinus
Finding|Finding|History of Present Illness|1434,1446|false|false|false|C0232201;C2041122|Sinus rhythm|sinus rhythm
Event|Event|History of Present Illness|1440,1446|false|false|false|||rhythm
Finding|Finding|History of Present Illness|1440,1446|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|History of Present Illness|1440,1446|false|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Attribute|Clinical Attribute|History of Present Illness|1460,1467|false|false|false|C0429104||T waves
Finding|Finding|History of Present Illness|1460,1467|false|false|false|C0429103|T wave feature|T waves
Event|Event|History of Present Illness|1462,1467|false|false|false|||waves
Phenomenon|Natural Phenomenon or Process|History of Present Illness|1462,1467|false|false|false|C0678544||waves
Anatomy|Body Location or Region|History of Present Illness|1473,1477|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|History of Present Illness|1473,1477|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|History of Present Illness|1473,1477|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|History of Present Illness|1473,1477|true|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|History of Present Illness|1473,1480|true|false|false|C0202691|CAT scan of head|head CT
Event|Event|History of Present Illness|1478,1480|true|false|false|||CT
Event|Event|History of Present Illness|1485,1493|true|false|false|||negative
Finding|Classification|History of Present Illness|1485,1493|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|History of Present Illness|1485,1493|true|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|History of Present Illness|1485,1493|true|false|false|C5237010|Expression Negative|negative
Finding|Finding|History of Present Illness|1485,1497|true|false|false|C0205160|Negative|negative for
Event|Event|History of Present Illness|1502,1507|true|false|false|||acute
Finding|Intellectual Product|History of Present Illness|1502,1507|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|History of Present Illness|1509,1518|true|false|false|||processes
Drug|Antibiotic|History of Present Illness|1533,1544|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Organic Chemical|History of Present Illness|1533,1544|false|false|false|C0007561|ceftriaxone|ceftriaxone
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1553,1568|false|false|false|C0021641|Insulin|regular insulin
Drug|Hormone|History of Present Illness|1553,1568|false|false|false|C0021641|Insulin|regular insulin
Drug|Pharmacologic Substance|History of Present Illness|1553,1568|false|false|false|C0021641|Insulin|regular insulin
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1561,1568|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|History of Present Illness|1561,1568|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|History of Present Illness|1561,1568|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|History of Present Illness|1561,1568|false|false|false|||insulin
Finding|Gene or Genome|History of Present Illness|1561,1568|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|History of Present Illness|1561,1568|false|false|false|C0202098|Insulin measurement|insulin
Drug|Biologically Active Substance|History of Present Illness|1575,1582|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Element, Ion, or Isotope|History of Present Illness|1575,1582|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Inorganic Chemical|History of Present Illness|1575,1582|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Pharmacologic Substance|History of Present Illness|1575,1582|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Drug|Vitamin|History of Present Illness|1575,1582|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|calcium
Event|Event|History of Present Illness|1575,1582|false|false|false|||calcium
Finding|Physiologic Function|History of Present Illness|1575,1582|false|false|false|C4553026|Calcium metabolic function|calcium
Procedure|Laboratory Procedure|History of Present Illness|1575,1582|false|false|false|C0201925|Calcium measurement|calcium
Drug|Organic Chemical|History of Present Illness|1575,1592|false|false|false|C0006699|calcium gluconate|calcium gluconate
Drug|Pharmacologic Substance|History of Present Illness|1575,1592|false|false|false|C0006699|calcium gluconate|calcium gluconate
Drug|Biologically Active Substance|History of Present Illness|1583,1592|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Organic Chemical|History of Present Illness|1583,1592|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Drug|Pharmacologic Substance|History of Present Illness|1583,1592|false|false|false|C0017714;C0220836|Gluconates;gluconate|gluconate
Event|Event|History of Present Illness|1593,1595|false|false|false|||1g
Drug|Organic Chemical|History of Present Illness|1597,1606|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|History of Present Illness|1597,1606|false|false|false|C0022957|lactulose|lactulose
Event|Event|History of Present Illness|1597,1606|false|false|false|||lactulose
Drug|Amino Acid, Peptide, or Protein|History of Present Illness|1628,1635|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|History of Present Illness|1628,1635|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|History of Present Illness|1628,1635|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|History of Present Illness|1628,1635|false|false|false|||albumin
Finding|Gene or Genome|History of Present Illness|1628,1635|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|History of Present Illness|1628,1635|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|History of Present Illness|1628,1635|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|History of Present Illness|1642,1650|false|false|false|||transfer
Finding|Functional Concept|History of Present Illness|1642,1650|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Finding|Idea or Concept|History of Present Illness|1642,1650|false|false|false|C0348011;C1555583;C1705822;C3244299|ActClass - transfer;Transfer - product ownership;Transfer Technique|transfer
Procedure|Health Care Activity|History of Present Illness|1642,1650|false|false|false|C4706767|Transfer (immobility management)|transfer
Event|Event|History of Present Illness|1652,1658|false|false|false|||vitals
Event|Activity|History of Present Illness|1692,1699|false|false|false|C1706079||arrival
Event|Event|History of Present Illness|1692,1699|false|false|false|||arrival
Finding|Functional Concept|History of Present Illness|1692,1699|false|false|false|C1555577|arrival - ActRelationshipType|arrival
Event|Event|History of Present Illness|1708,1712|false|false|false|||MICU
Finding|Body Substance|History of Present Illness|1714,1721|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|History of Present Illness|1714,1721|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|History of Present Illness|1714,1721|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Attribute|Clinical Attribute|History of Present Illness|1731,1736|false|false|false|C5890168||alert
Drug|Organic Chemical|History of Present Illness|1731,1736|false|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|History of Present Illness|1731,1736|false|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|History of Present Illness|1731,1736|false|false|false|||alert
Finding|Finding|History of Present Illness|1731,1736|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|History of Present Illness|1731,1736|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|History of Present Illness|1731,1736|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|History of Present Illness|1741,1751|false|false|false|||conversant
Anatomy|Body Location or Region|History of Present Illness|1765,1774|true|false|false|C0000726|Abdomen|abdominal
Finding|Sign or Symptom|History of Present Illness|1765,1779|true|false|false|C0000737|Abdominal Pain|abdominal pain
Attribute|Clinical Attribute|History of Present Illness|1775,1779|true|false|false|C2598155||pain
Event|Event|History of Present Illness|1775,1779|true|false|false|||pain
Finding|Functional Concept|History of Present Illness|1775,1779|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1775,1779|true|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Attribute|Clinical Attribute|History of Present Illness|1781,1787|true|false|false|C4255480||nausea
Event|Event|History of Present Illness|1781,1787|true|false|false|||nausea
Finding|Sign or Symptom|History of Present Illness|1781,1787|true|false|false|C0027497|Nausea|nausea
Event|Event|History of Present Illness|1789,1797|true|false|false|||vomiting
Finding|Sign or Symptom|History of Present Illness|1789,1797|true|false|false|C0042963|Vomiting|vomiting
Anatomy|Body Location or Region|History of Present Illness|1799,1804|false|false|false|C0817096;C1527391|Anterior thoracic region;Chest|chest
Finding|Finding|History of Present Illness|1799,1804|false|false|false|C0741025|Chest problem|chest
Attribute|Clinical Attribute|History of Present Illness|1799,1809|false|false|true|C2926613||chest pain
Finding|Sign or Symptom|History of Present Illness|1799,1809|false|false|true|C0008031|Chest Pain|chest pain
Attribute|Clinical Attribute|History of Present Illness|1805,1809|false|true|false|C2598155||pain
Event|Event|History of Present Illness|1805,1809|false|false|false|||pain
Finding|Functional Concept|History of Present Illness|1805,1809|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|History of Present Illness|1805,1809|false|true|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Event|Event|History of Present Illness|1814,1824|false|false|false|||difficulty
Finding|Finding|History of Present Illness|1814,1824|false|false|false|C1299586|Has difficulty doing (qualifier value)|difficulty
Attribute|Clinical Attribute|History of Present Illness|1826,1835|false|false|false|C5885990||breathing
Event|Event|History of Present Illness|1826,1835|false|false|false|||breathing
Finding|Finding|History of Present Illness|1826,1835|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Organism Function|History of Present Illness|1826,1835|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Finding|Physiologic Function|History of Present Illness|1826,1835|false|false|false|C0004048;C0035203;C2015926|Inspiration (function);Respiration;outcomes otolaryngology breathing|breathing
Phenomenon|Biologic Function|History of Present Illness|1826,1835|false|false|false|C1160636|respiratory system process|breathing
Finding|Intellectual Product|History of Present Illness|1847,1854|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|History of Present Illness|1847,1854|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Finding|Sign or Symptom|History of Present Illness|1847,1860|true|false|false|C0010201|Chronic Cough|chronic cough
Drug|Organic Chemical|History of Present Illness|1855,1860|true|false|false|C3815497|Cough (guaifenesin)|cough
Drug|Pharmacologic Substance|History of Present Illness|1855,1860|true|false|false|C3815497|Cough (guaifenesin)|cough
Event|Event|History of Present Illness|1855,1860|true|false|false|||cough
Finding|Sign or Symptom|History of Present Illness|1855,1860|true|false|false|C0010200|Coughing|cough
Finding|Finding|History of Present Illness|1873,1877|true|false|false|C4281574|Much|much
Event|Event|History of Present Illness|1878,1885|true|false|false|||changed
Event|Event|History of Present Illness|1908,1913|true|false|false|||fever
Finding|Finding|History of Present Illness|1908,1913|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1908,1913|true|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|History of Present Illness|1908,1923|true|false|false|C5570922|Fever or chills|fever or chills
Event|Event|History of Present Illness|1917,1923|true|false|false|||chills
Finding|Sign or Symptom|History of Present Illness|1917,1923|true|false|false|C0085593|Chills|chills
Event|Event|History of Present Illness|1929,1936|false|false|false|||reports
Event|Event|History of Present Illness|1937,1943|false|false|false|||taking
Attribute|Clinical Attribute|History of Present Illness|1956,1967|false|false|false|C0802604;C2598133||medications
Drug|Pharmacologic Substance|History of Present Illness|1956,1967|false|false|false|C0013227|Pharmaceutical Preparations|medications
Event|Event|History of Present Illness|1956,1967|false|false|false|||medications
Finding|Intellectual Product|History of Present Illness|1956,1967|false|false|false|C4284232|Medications|medications
Drug|Organic Chemical|History of Present Illness|1979,1988|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|History of Present Illness|1979,1988|false|false|false|C0022957|lactulose|lactulose
Event|Event|History of Present Illness|1979,1988|false|false|false|||lactulose
Event|Event|History of Present Illness|2007,2012|false|false|false|||taste
Finding|Organ or Tissue Function|History of Present Illness|2007,2012|false|false|false|C0039336|Taste Perception|taste
Event|Event|History of Present Illness|2014,2024|false|false|false|||disgusting
Finding|Mental Process|History of Present Illness|2014,2024|false|false|false|C0683283|Disgust|disgusting
Disorder|Disease or Syndrome|Past Medical History|2054,2057|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|Past Medical History|2054,2057|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|Past Medical History|2054,2057|false|false|false|||HCV
Disorder|Disease or Syndrome|Past Medical History|2058,2067|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|Past Medical History|2058,2067|false|false|false|||Cirrhosis
Event|Event|Past Medical History|2069,2077|false|false|false|||genotype
Procedure|Laboratory Procedure|Past Medical History|2069,2077|false|false|false|C1285573|Genotype determination|genotype
Disorder|Disease or Syndrome|Past Medical History|2085,2088|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Past Medical History|2085,2088|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Past Medical History|2085,2088|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Past Medical History|2085,2088|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Past Medical History|2085,2088|false|false|false|||HIV
Event|Event|Past Medical History|2093,2098|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2093,2098|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Drug|Amino Acid, Peptide, or Protein|Past Medical History|2104,2107|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Biologically Active Substance|Past Medical History|2104,2107|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Immunologic Factor|Past Medical History|2104,2107|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Finding|Gene or Genome|Past Medical History|2104,2107|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Finding|Receptor|Past Medical History|2104,2107|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Procedure|Laboratory Procedure|Past Medical History|2104,2113|false|false|false|C0243009;C3541261|CD4 Count determination procedure;CD4 Expressing Cell Count|CD4 count
Event|Event|Past Medical History|2108,2113|false|false|false|||count
Disorder|Disease or Syndrome|Past Medical History|2123,2126|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|Past Medical History|2123,2126|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|Past Medical History|2123,2126|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|Past Medical History|2123,2126|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|Past Medical History|2123,2126|false|false|false|||HIV
Procedure|Laboratory Procedure|Past Medical History|2123,2137|false|false|false|C1168369|HIV viral load|HIV viral load
Finding|Functional Concept|Past Medical History|2127,2132|false|false|false|C0521026|Viral|viral
Finding|Finding|Past Medical History|2127,2137|false|false|false|C0376705|Viral Load result|viral load
Procedure|Laboratory Procedure|Past Medical History|2127,2137|false|false|false|C1261478|Viral load (procedure)|viral load
Event|Activity|Past Medical History|2133,2137|false|false|false|C1708715|Loading Technique|load
Event|Event|Past Medical History|2133,2137|false|false|false|||load
Finding|Idea or Concept|Past Medical History|2133,2137|false|false|false|C1550025|Load - Remote control command|load
Attribute|Clinical Attribute|Past Medical History|2139,2151|false|false|false|C3827727|Undetectable|undetectable
Disorder|Disease or Syndrome|Past Medical History|2156,2160|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|Past Medical History|2156,2160|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|Past Medical History|2156,2160|false|false|false|||COPD
Finding|Gene or Genome|Past Medical History|2156,2160|false|false|false|C1412502|ARCN1 gene|COPD
Anatomy|Body Location or Region|Past Medical History|2166,2169|false|false|false|C5239891|area PFt|PFT
Drug|Indicator, Reagent, or Diagnostic Aid|Past Medical History|2166,2169|false|false|false|C0053122|bentiromide|PFT
Drug|Pharmacologic Substance|Past Medical History|2166,2169|false|false|false|C0053122|bentiromide|PFT
Event|Event|Past Medical History|2166,2169|false|false|false|||PFT
Procedure|Diagnostic Procedure|Past Medical History|2166,2169|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Procedure|Therapeutic or Preventive Procedure|Past Medical History|2166,2169|false|false|false|C0024119;C0279232|Pulmonary function tests;fluorouracil/melphalan/tamoxifen|PFT
Event|Event|Past Medical History|2170,2176|false|false|false|||showed
Event|Event|Past Medical History|2177,2180|false|false|false|||FVC
Lab|Laboratory or Test Result|Past Medical History|2177,2180|false|false|false|C3714541|Forced Vital Capacity|FVC
Attribute|Clinical Attribute|Past Medical History|2193,2197|false|false|false|C0802965||FEV1
Event|Event|Past Medical History|2193,2197|false|false|false|||FEV1
Procedure|Diagnostic Procedure|Past Medical History|2193,2197|false|false|false|C0849974|Pulmonary Function Test/Forced Expiratory Volume 1|FEV1
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2233,2259|false|false|false|C0005586;C1839839;C1852197;C1970943;C1970945;C2700438;C2700439;C2700440|Bipolar Disorder;MAJOR AFFECTIVE DISORDER 1;MAJOR AFFECTIVE DISORDER 2;MAJOR AFFECTIVE DISORDER 4;MAJOR AFFECTIVE DISORDER 6;MAJOR AFFECTIVE DISORDER 7;MAJOR AFFECTIVE DISORDER 8;MAJOR AFFECTIVE DISORDER 9|Bipolar Affective Disorder
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2241,2259|false|false|false|C0525045|Mood Disorders|Affective Disorder
Disorder|Disease or Syndrome|Past Medical History|2251,2259|false|false|false|C0012634|Disease|Disorder
Event|Event|Past Medical History|2251,2259|false|false|false|||Disorder
Disorder|Disease or Syndrome|Past Medical History|2264,2268|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2264,2268|false|false|false|C0038436;C0878676|6-pyruvoyl-tetrahydropterin synthase deficiency;Post-Traumatic Stress Disorder|PTSD
Event|Event|Past Medical History|2264,2268|false|false|false|||PTSD
Disorder|Injury or Poisoning|Past Medical History|2279,2286|false|false|false|C0274659|Poisoning by cocaine|cocaine
Drug|Biomedical or Dental Material|Past Medical History|2279,2286|false|false|false|C0009170|cocaine|cocaine
Drug|Hazardous or Poisonous Substance|Past Medical History|2279,2286|false|false|false|C0009170|cocaine|cocaine
Drug|Organic Chemical|Past Medical History|2279,2286|false|false|false|C0009170|cocaine|cocaine
Drug|Pharmacologic Substance|Past Medical History|2279,2286|false|false|false|C0009170|cocaine|cocaine
Event|Event|Past Medical History|2279,2286|false|false|false|||cocaine
Procedure|Laboratory Procedure|Past Medical History|2279,2286|false|false|false|C0202362|Cocaine measurement|cocaine
Disorder|Injury or Poisoning|Past Medical History|2291,2297|false|false|false|C0161541|Poisoning by heroin|heroin
Drug|Hazardous or Poisonous Substance|Past Medical History|2291,2297|false|false|false|C0011892|heroin|heroin
Drug|Organic Chemical|Past Medical History|2291,2297|false|false|false|C0011892|heroin|heroin
Drug|Pharmacologic Substance|Past Medical History|2291,2297|false|false|false|C0011892|heroin|heroin
Event|Event|Past Medical History|2291,2297|false|false|false|||heroin
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2291,2303|false|false|false|C0600241|heroin abuse|heroin abuse
Disorder|Mental or Behavioral Dysfunction|Past Medical History|2298,2303|false|false|false|C0013146|Drug abuse|abuse
Event|Event|Past Medical History|2298,2303|false|false|false|||abuse
Event|Event|Past Medical History|2298,2303|false|false|false|C1546935|Abuse|abuse
Finding|Finding|Past Medical History|2298,2303|false|false|false|C0562381|Victim of abuse (finding)|abuse
Disorder|Neoplastic Process|Past Medical History|2311,2325|false|false|false|C0007114|Malignant neoplasm of skin|of skin cancer
Anatomy|Body System|Past Medical History|2314,2318|false|false|false|C1123023;C4520765|Skin;Skin, Human|skin
Disorder|Disease or Syndrome|Past Medical History|2314,2318|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Disorder|Neoplastic Process|Past Medical History|2314,2318|false|false|false|C0178298;C0496955|Neoplasm of uncertain or unknown behavior of skin;Skin and subcutaneous tissue disorders|skin
Finding|Body Substance|Past Medical History|2314,2318|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Finding|Intellectual Product|Past Medical History|2314,2318|false|false|false|C0444099;C1546781|Skin Specimen;Skin Specimen Source Code|skin
Disorder|Neoplastic Process|Past Medical History|2314,2325|false|false|false|C0007114|Malignant neoplasm of skin|skin cancer
Disorder|Neoplastic Process|Past Medical History|2319,2325|false|false|false|C0006826|Malignant Neoplasms|cancer
Event|Event|Past Medical History|2319,2325|false|false|false|||cancer
Finding|Body Substance|Past Medical History|2330,2337|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|Past Medical History|2330,2337|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|2330,2337|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|Past Medical History|2330,2344|false|false|false|C0747307|Patient-Reported|patient report
Attribute|Clinical Attribute|Past Medical History|2338,2344|false|false|false|C4255046||report
Event|Event|Past Medical History|2338,2344|false|false|false|||report
Finding|Intellectual Product|Past Medical History|2338,2344|false|false|false|C0684224|Report (document)|report
Procedure|Health Care Activity|Past Medical History|2338,2344|false|false|false|C0700287|Reporting|report
Event|Event|Family Medical History|2431,2438|true|false|false|||talking
Finding|Conceptual Entity|Family Medical History|2474,2481|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Finding|Idea or Concept|Family Medical History|2474,2481|false|false|false|C1546493;C1704648|Brother - courtesy title;Relationship - Brother|brother
Event|Event|Family Medical History|2498,2503|false|false|false|||touch
Finding|Mental Process|Family Medical History|2498,2503|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Finding|Organ or Tissue Function|Family Medical History|2498,2503|false|false|false|C0702221;C2350522|Touch Perception;Touch sensation|touch
Procedure|Therapeutic or Preventive Procedure|Family Medical History|2498,2503|false|false|false|C0152054|Therapeutic Touch|touch
Event|Event|Family Medical History|2514,2519|false|false|false|||lives
Event|Event|Family Medical History|2539,2544|true|false|false|||aware
Finding|Mental Process|Family Medical History|2539,2544|true|false|false|C0004448|Awareness|aware
Anatomy|Body Part, Organ, or Organ Component|Family Medical History|2564,2569|true|false|false|C0023884;C1278929;C4037986|Abdomen>Liver;Liver|liver
Disorder|Disease or Syndrome|Family Medical History|2564,2569|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Disorder|Neoplastic Process|Family Medical History|2564,2569|true|false|false|C0023895;C0496870|Benign neoplasm of liver;Liver diseases|liver
Drug|Organic Chemical|Family Medical History|2564,2569|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Pharmacologic Substance|Family Medical History|2564,2569|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Drug|Vitamin|Family Medical History|2564,2569|true|false|false|C0023899;C0721399|Liver brand of Vitamin B 12;liver extract|liver
Event|Event|Family Medical History|2564,2569|true|false|false|||liver
Finding|Finding|Family Medical History|2564,2569|true|false|false|C0577060|Liver problem|liver
Procedure|Health Care Activity|Family Medical History|2564,2569|true|false|false|C0872387|Procedures on liver|liver
Disorder|Disease or Syndrome|Family Medical History|2571,2578|true|false|false|C0012634|Disease|disease
Event|Event|Family Medical History|2571,2578|true|false|false|||disease
Drug|Amino Acid, Peptide, or Protein|Family Medical History|2582,2592|false|false|false|C3812393|ErbB Receptors|her family
Drug|Enzyme|Family Medical History|2582,2592|false|false|false|C3812393|ErbB Receptors|her family
Finding|Receptor|Family Medical History|2582,2592|false|false|false|C3812393|ErbB Receptors|her family
Finding|Classification|Family Medical History|2586,2592|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Conceptual Entity|Family Medical History|2586,2592|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Idea or Concept|Family Medical History|2586,2592|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Finding|Intellectual Product|Family Medical History|2586,2592|false|false|false|C1301584;C1546847;C1563343;C1704727;C2700055|Entity Name Part Type - family;Family (taxonomic);Family Collection;Last Name;Living Arrangement - Family|family
Procedure|Health Care Activity|General Exam|2613,2622|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|2623,2631|false|false|false|||PHYSICAL
Finding|Finding|General Exam|2623,2631|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|2623,2631|false|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|2623,2631|false|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|2623,2636|false|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|2623,2636|false|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|2632,2636|false|false|false|||EXAM
Finding|Functional Concept|General Exam|2632,2636|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|2632,2636|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|2694,2701|false|false|false|||GENERAL
Finding|Classification|General Exam|2694,2701|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|GENERAL
Procedure|Health Care Activity|General Exam|2694,2701|false|false|false|C3812897|General medical service|GENERAL
Attribute|Clinical Attribute|General Exam|2703,2708|true|false|false|C5890168||Alert
Drug|Organic Chemical|General Exam|2703,2708|true|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|General Exam|2703,2708|true|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|General Exam|2703,2708|true|false|false|||Alert
Finding|Finding|General Exam|2703,2708|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|General Exam|2703,2708|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|General Exam|2703,2708|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|General Exam|2710,2718|true|false|false|||oriented
Finding|Intellectual Product|General Exam|2723,2728|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|2729,2737|true|false|false|||distress
Finding|Finding|General Exam|2729,2737|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|2729,2737|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Part, Organ, or Organ Component|General Exam|2740,2745|true|false|false|C0024109|Lung|LUNGS
Event|Event|General Exam|2747,2756|false|false|false|||Decreased
Drug|Inorganic Chemical|General Exam|2757,2760|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Pharmacologic Substance|General Exam|2757,2760|false|false|false|C0001861;C3536832|Air (substance);air|air
Drug|Substance|General Exam|2757,2760|false|false|false|C0001861;C3536832|Air (substance);air|air
Finding|Finding|General Exam|2757,2760|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Gene or Genome|General Exam|2757,2760|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Finding|Intellectual Product|General Exam|2757,2760|false|false|false|C1140091;C1866503;C2681903|ACUTE INSULIN RESPONSE;AI/RHEUM;AIRN gene|air
Phenomenon|Natural Phenomenon or Process|General Exam|2757,2769|false|false|false|C0001868|Air Movements|air movement
Event|Event|General Exam|2761,2769|false|false|false|||movement
Finding|Organism Function|General Exam|2761,2769|false|false|false|C0026649|Movement|movement
Event|Event|General Exam|2778,2783|false|false|false|||sides
Event|Event|General Exam|2785,2794|false|false|false|||scattered
Finding|Organism Function|General Exam|2796,2806|false|false|false|C0231800|Expiration, Respiratory|expiratory
Finding|Sign or Symptom|General Exam|2796,2814|false|false|false|C0231875|Expiratory wheezing|expiratory wheezes
Event|Event|General Exam|2807,2814|false|false|false|||wheezes
Finding|Sign or Symptom|General Exam|2807,2814|false|false|false|C0043144|Wheezing|wheezes
Event|Activity|General Exam|2829,2833|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|2829,2833|false|false|false|||rate
Finding|Idea or Concept|General Exam|2829,2833|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|2838,2844|true|false|false|||rhythm
Finding|Finding|General Exam|2838,2844|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|2838,2844|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|2863,2870|true|false|false|||murmurs
Finding|Finding|General Exam|2863,2870|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|2872,2876|true|false|false|||rubs
Finding|Finding|General Exam|2872,2876|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|2879,2886|true|false|false|||gallops
Anatomy|Body Location or Region|General Exam|2889,2892|false|false|false|C0000726;C0449202|ABD (body structure);Abdomen|ABD
Disorder|Cell or Molecular Dysfunction|General Exam|2889,2892|false|false|false|C3811055|Absence of Biallelic TCRgamma Deletion|ABD
Event|Event|General Exam|2889,2892|false|false|false|||ABD
Disorder|Disease or Syndrome|General Exam|2894,2898|false|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|Soft
Event|Event|General Exam|2894,2898|false|false|false|||Soft
Event|Event|General Exam|2912,2921|false|false|false|||distended
Finding|Finding|General Exam|2912,2921|false|false|false|C0700124|Dilated|distended
Anatomy|Body Location or Region|General Exam|2923,2928|false|false|false|C0230171|Flank (surface region)|flank
Event|Event|General Exam|2929,2937|false|false|false|||dullness
Finding|Finding|General Exam|2929,2937|false|false|false|C0541911|Dullness|dullness
Anatomy|Body Part, Organ, or Organ Component|General Exam|2952,2957|false|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|2952,2964|false|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|2958,2964|false|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|2958,2964|false|false|false|C0037709||sounds
Finding|Finding|General Exam|2965,2972|false|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|2965,2972|false|false|false|C0150312;C0449450|Present;Presentation|present
Disorder|Congenital Abnormality|General Exam|2975,2978|false|false|false|C0015306|Hereditary Multiple Exostoses|EXT
Event|Event|General Exam|2975,2978|false|false|false|||EXT
Finding|Gene or Genome|General Exam|2975,2978|false|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|EXT
Event|Event|General Exam|2980,2984|false|false|false|||Warm
Finding|Finding|General Exam|2980,2984|false|false|false|C0582051|Feels warm|Warm
Phenomenon|Natural Phenomenon or Process|General Exam|2980,2984|false|false|false|C0687712|warming process|Warm
Finding|Finding|General Exam|2986,2990|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|2991,2999|true|false|false|||perfused
Drug|Food|General Exam|3004,3010|true|false|false|C5890763||pulses
Event|Event|General Exam|3004,3010|true|false|false|||pulses
Finding|Physiologic Function|General Exam|3004,3010|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3004,3010|true|false|false|C0034107|Pulse taking|pulses
Event|Event|General Exam|3015,3023|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3015,3023|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|3027,3032|true|false|false|C1717255||edema
Event|Event|General Exam|3027,3032|true|false|false|||edema
Finding|Pathologic Function|General Exam|3027,3032|true|false|false|C0013604|Edema|edema
Finding|Body Substance|General Exam|3036,3045|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|3036,3045|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|3036,3045|true|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|3036,3045|true|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|3046,3054|true|false|false|||PHYSICAL
Finding|Finding|General Exam|3046,3054|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Finding|Functional Concept|General Exam|3046,3054|true|false|false|C0205485;C1509143|Physical;physical examination (physical finding)|PHYSICAL
Procedure|Health Care Activity|General Exam|3046,3054|true|false|false|C0031809|Physical Examination|PHYSICAL
Finding|Finding|General Exam|3046,3059|true|false|false|C1509143|physical examination (physical finding)|PHYSICAL EXAM
Procedure|Health Care Activity|General Exam|3046,3059|true|false|false|C0031809|Physical Examination|PHYSICAL EXAM
Event|Event|General Exam|3055,3059|false|false|false|||EXAM
Finding|Functional Concept|General Exam|3055,3059|false|false|false|C4284036|Exam|EXAM
Procedure|Health Care Activity|General Exam|3055,3059|false|false|false|C0582103|Medical Examination|EXAM
Event|Event|General Exam|3121,3124|false|false|false|||7BM
Finding|Classification|General Exam|3128,3135|false|false|false|C4521767|United States Military Commissioned Officer O10 (qualifier value)|General
Procedure|Health Care Activity|General Exam|3128,3135|false|false|false|C3812897|General medical service|General
Finding|Sign or Symptom|General Exam|3137,3146|false|false|false|C0006625|Cachexia|Cachectic
Attribute|Clinical Attribute|General Exam|3164,3169|true|false|false|C5890168||alert
Drug|Organic Chemical|General Exam|3164,3169|true|false|false|C0718338|Alert brand of caffeine|alert
Drug|Pharmacologic Substance|General Exam|3164,3169|true|false|false|C0718338|Alert brand of caffeine|alert
Event|Event|General Exam|3164,3169|true|false|false|||alert
Finding|Finding|General Exam|3164,3169|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Functional Concept|General Exam|3164,3169|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Finding|Intellectual Product|General Exam|3164,3169|true|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|alert
Event|Event|General Exam|3171,3179|true|false|false|||oriented
Finding|Finding|General Exam|3171,3179|true|false|false|C1961028|Oriented to place|oriented
Event|Event|General Exam|3184,3189|true|false|false|||acute
Finding|Intellectual Product|General Exam|3184,3189|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|3191,3199|true|false|false|||distress
Finding|Finding|General Exam|3191,3199|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Finding|Mental Process|General Exam|3191,3199|true|false|false|C0231303;C0700361|Distress;Emotional distress|distress
Anatomy|Body Location or Region|General Exam|3202,3207|true|false|false|C1512338|HEENT|HEENT
Anatomy|Body Part, Organ, or Organ Component|General Exam|3209,3215|true|false|false|C0036410|Sclera|Sclera
Disorder|Disease or Syndrome|General Exam|3209,3215|true|false|false|C0036412|Scleral Diseases|Sclera
Event|Event|General Exam|3209,3215|true|false|false|||Sclera
Procedure|Health Care Activity|General Exam|3209,3215|true|false|false|C2228481|examination of sclera|Sclera
Event|Event|General Exam|3216,3225|false|false|false|||anicteric
Finding|Finding|General Exam|3216,3225|false|false|false|C0205180|Anicteric|anicteric
Anatomy|Body Part, Organ, or Organ Component|General Exam|3227,3230|false|false|false|C0694605|Medial part of medial mammillary nucleus|MMM
Disorder|Neoplastic Process|General Exam|3227,3230|false|false|false|C0026987|Myelofibrosis|MMM
Anatomy|Body Location or Region|General Exam|3232,3242|false|false|false|C0521367|Oropharyngeal|oropharynx
Event|Event|General Exam|3243,3248|false|false|false|||clear
Finding|Idea or Concept|General Exam|3243,3248|false|false|false|C1550016|Remote control command - Clear|clear
Finding|Intellectual Product|General Exam|3250,3254|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Finding|Sign or Symptom|General Exam|3250,3264|false|false|false|C0149758|Poor dentition|poor dentition
Anatomy|Body Part, Organ, or Organ Component|General Exam|3255,3264|false|false|false|C0011443;C0040426|Dentition;Tooth structure|dentition
Finding|Idea or Concept|General Exam|3271,3278|false|false|false|C1550516|Target Awareness - partial|partial
Event|Event|General Exam|3279,3287|true|false|false|||dentures
Finding|Finding|General Exam|3279,3287|true|false|false|C2266651|dentures (physical finding)|dentures
Procedure|Therapeutic or Preventive Procedure|General Exam|3279,3287|true|false|false|C2064697|dentures (treatment)|dentures
Anatomy|Body Location or Region|General Exam|3290,3294|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Anatomy|Cell Component|General Exam|3290,3294|true|false|false|C0027530;C3159206|Neck;dendritic spine neck|Neck
Finding|Finding|General Exam|3290,3294|true|false|false|C0684335;C0812434|Neck problem;Passive joint movement of neck (finding)|Neck
Event|Event|General Exam|3296,3302|true|false|false|||supple
Finding|Functional Concept|General Exam|3296,3302|true|false|false|C0332254|Supple|supple
Event|Event|General Exam|3304,3307|true|false|false|||JVP
Finding|Finding|General Exam|3304,3307|true|false|false|C0428897|Jugular venous pressure|JVP
Event|Event|General Exam|3312,3320|true|false|false|||elevated
Anatomy|Body Part, Organ, or Organ Component|General Exam|3325,3328|true|false|false|C0226032|Anterior descending branch of left coronary artery|LAD
Disorder|Disease or Syndrome|General Exam|3325,3328|true|false|false|C0398738;C5550999|Leukocyte adhesion deficiency;Leukocyte adhesion deficiency type 1|LAD
Event|Event|General Exam|3325,3328|true|false|false|||LAD
Finding|Gene or Genome|General Exam|3325,3328|true|false|false|C1414063;C1706333|DLD gene;ITGB2 wt Allele|LAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|3331,3336|true|false|false|C0024109|Lung|Lungs
Event|Event|General Exam|3338,3343|true|false|false|||Clear
Finding|Idea or Concept|General Exam|3338,3343|true|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|General Exam|3347,3359|true|false|false|||auscultation
Procedure|Diagnostic Procedure|General Exam|3347,3359|true|false|false|C0004339|Auscultation|auscultation
Event|Event|General Exam|3376,3383|true|false|false|||wheezes
Finding|Sign or Symptom|General Exam|3376,3383|true|false|false|C0043144|Wheezing|wheezes
Event|Event|General Exam|3385,3390|true|false|false|||rales
Finding|Finding|General Exam|3385,3390|true|false|false|C0034642;C0240859|Basilar Rales;Rales|rales
Event|Activity|General Exam|3414,3418|false|false|false|C0871208|Rating (action)|rate
Event|Event|General Exam|3414,3418|false|false|false|||rate
Finding|Idea or Concept|General Exam|3414,3418|false|false|false|C1549480|Amount type - Rate|rate
Event|Event|General Exam|3423,3429|true|false|false|||rhythm
Finding|Finding|General Exam|3423,3429|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Finding|Physiologic Function|General Exam|3423,3429|true|false|false|C0871269;C1523018|Rhythm;rhythmic process (biological)|rhythm
Event|Event|General Exam|3450,3457|true|false|false|||murmurs
Finding|Finding|General Exam|3450,3457|true|false|false|C0018808|Heart murmur|murmurs
Event|Event|General Exam|3459,3463|true|false|false|||rubs
Finding|Finding|General Exam|3459,3463|true|false|false|C0232267|Pericardial friction rub|rubs
Event|Event|General Exam|3466,3473|true|false|false|||gallops
Anatomy|Body Location or Region|General Exam|3476,3483|false|false|false|C0000726;C0230168|Abdomen;Abdominal Cavity|Abdomen
Disorder|Neoplastic Process|General Exam|3476,3483|false|false|false|C0153662|Malignant neoplasm of abdomen|Abdomen
Finding|Finding|General Exam|3476,3483|false|false|false|C0941288|Abdomen problem|Abdomen
Event|Event|General Exam|3492,3501|false|false|false|||distended
Finding|Finding|General Exam|3492,3501|false|false|false|C0700124|Dilated|distended
Anatomy|Body Part, Organ, or Organ Component|General Exam|3524,3529|true|false|false|C0021853|Intestines|bowel
Finding|Finding|General Exam|3524,3536|true|false|false|C0232693|Bowel sounds|bowel sounds
Event|Event|General Exam|3530,3536|true|false|false|||sounds
Phenomenon|Natural Phenomenon or Process|General Exam|3530,3536|true|false|false|C0037709||sounds
Event|Event|General Exam|3538,3545|true|false|false|||present
Finding|Finding|General Exam|3538,3545|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Idea or Concept|General Exam|3538,3545|true|false|false|C0150312;C0449450|Present;Presentation|present
Finding|Sign or Symptom|General Exam|3550,3568|true|false|false|C0234246|Rebound tenderness|rebound tenderness
Event|Event|General Exam|3558,3568|true|false|false|||tenderness
Finding|Mental Process|General Exam|3558,3568|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Finding|Sign or Symptom|General Exam|3558,3568|true|false|false|C0234233;C0684239|Emotional tenderness;Sore to touch|tenderness
Event|Event|General Exam|3572,3580|true|false|false|||guarding
Finding|Finding|General Exam|3572,3580|true|false|false|C0427198|Protective muscle spasm|guarding
Event|Event|General Exam|3590,3595|true|false|false|||foley
Disorder|Congenital Abnormality|General Exam|3598,3601|true|false|false|C0015306|Hereditary Multiple Exostoses|Ext
Event|Event|General Exam|3598,3601|true|false|false|||Ext
Finding|Gene or Genome|General Exam|3598,3601|true|false|false|C0694878;C1707871|EXT1 gene;EXT1 wt Allele|Ext
Event|Event|General Exam|3603,3607|true|false|false|||warm
Finding|Finding|General Exam|3603,3607|true|false|false|C0582051|Feels warm|warm
Phenomenon|Natural Phenomenon or Process|General Exam|3603,3607|true|false|false|C0687712|warming process|warm
Finding|Finding|General Exam|3609,3613|true|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|3614,3622|true|false|false|||perfused
Drug|Food|General Exam|3627,3633|true|false|false|C5890763||pulses
Event|Event|General Exam|3627,3633|true|false|false|||pulses
Finding|Physiologic Function|General Exam|3627,3633|true|false|false|C0391850|Physiologic pulse|pulses
Procedure|Health Care Activity|General Exam|3627,3633|true|false|false|C0034107|Pulse taking|pulses
Disorder|Anatomical Abnormality|General Exam|3638,3646|true|false|false|C0149651|Clubbing|clubbing
Event|Event|General Exam|3638,3646|true|false|false|||clubbing
Event|Event|General Exam|3648,3656|true|false|false|||cyanosis
Finding|Sign or Symptom|General Exam|3648,3656|true|false|false|C0010520|Cyanosis|cyanosis
Attribute|Clinical Attribute|General Exam|3661,3666|true|false|false|C1717255||edema
Event|Event|General Exam|3661,3666|true|false|false|||edema
Finding|Pathologic Function|General Exam|3661,3666|true|false|false|C0013604|Edema|edema
Event|Event|General Exam|3685,3694|true|false|false|||asterixis
Finding|Sign or Symptom|General Exam|3685,3694|true|false|false|C0232766|Asterixis|asterixis
Procedure|Health Care Activity|General Exam|3719,3728|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|ADMISSION
Event|Event|General Exam|3729,3733|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|3729,3733|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|3765,3770|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3765,3770|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3765,3770|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|3771,3774|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|3779,3782|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|3779,3782|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|3779,3782|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|3789,3792|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|3789,3792|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|3789,3792|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|3789,3792|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|3798,3801|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|3798,3801|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|3808,3811|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|3808,3811|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|3808,3811|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|3808,3811|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|3808,3811|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|3817,3820|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|3817,3820|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|3817,3820|false|false|false|||MCH
Finding|Gene or Genome|General Exam|3817,3820|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|3817,3820|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|3817,3820|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|3827,3831|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|3837,3840|false|false|false|||RDW
Procedure|Laboratory Procedure|General Exam|3847,3850|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|3867,3872|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3867,3872|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3867,3872|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Finding|Body Substance|General Exam|3885,3891|false|false|false|C0024202|Lymph|Lymphs
Drug|Antibiotic|General Exam|3898,3903|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Biomedical or Dental Material|General Exam|3898,3903|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Drug|Organic Chemical|General Exam|3898,3903|false|false|false|C0540173;C3275179|Mono-S;Monos|Monos
Disorder|Disease or Syndrome|General Exam|3909,3912|false|false|false|C0272192;C1836122|Familial eosinophilia;SARCOIDOSIS, EARLY-ONSET|Eos
Finding|Gene or Genome|General Exam|3909,3912|false|false|false|C1421861;C1538729|IKZF4 gene;PRSS33 gene|Eos
Disorder|Disease or Syndrome|General Exam|3938,3943|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3938,3943|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3938,3943|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|3948,3951|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|3948,3951|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|3948,3951|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|3973,3978|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|3973,3978|false|false|false|||BLOOD
Finding|Body Substance|General Exam|3973,3978|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|3973,3986|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|3973,3986|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|3973,3986|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|3979,3986|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|3979,3986|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|3979,3986|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|3979,3986|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|3979,3986|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|3979,3986|false|false|false|C0337438|Glucose measurement|Glucose
Disorder|Disease or Syndrome|General Exam|4064,4069|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4064,4069|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4064,4069|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4070,4073|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4070,4073|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4070,4073|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4070,4073|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4070,4073|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4070,4073|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4070,4073|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4070,4073|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4079,4082|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4079,4082|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4079,4082|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4079,4082|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4079,4082|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|4079,4082|false|false|false|||AST
Finding|Gene or Genome|General Exam|4079,4082|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4088,4095|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4088,4095|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4127,4132|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4127,4132|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4127,4132|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4127,4140|false|false|false|C0853248|Blood albumin|BLOOD Albumin
Drug|Amino Acid, Peptide, or Protein|General Exam|4133,4140|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Biologically Active Substance|General Exam|4133,4140|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Drug|Pharmacologic Substance|General Exam|4133,4140|false|false|false|C0001924;C5966160|Albumin;Albumins|Albumin
Event|Event|General Exam|4133,4140|false|false|false|||Albumin
Finding|Gene or Genome|General Exam|4133,4140|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Finding|Physiologic Function|General Exam|4133,4140|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|Albumin
Procedure|Laboratory Procedure|General Exam|4133,4140|false|false|false|C0201838|Albumin measurement|Albumin
Event|Event|General Exam|4146,4153|false|false|false|||IMAGING
Finding|Finding|General Exam|4146,4153|false|false|false|C0740845|Imaging problem|IMAGING
Procedure|Diagnostic Procedure|General Exam|4146,4153|false|false|false|C0011923;C0079595|Diagnostic Imaging;Imaging Techniques|IMAGING
Event|Event|General Exam|4154,4161|false|false|false|||STUDIES
Procedure|Research Activity|General Exam|4154,4161|false|false|false|C0947630|Scientific Study|STUDIES
Attribute|Clinical Attribute|General Exam|4184,4191|false|false|false|C0881943||CT HEAD
Procedure|Diagnostic Procedure|General Exam|4184,4191|false|false|false|C0202691|CAT scan of head|CT HEAD
Anatomy|Body Location or Region|General Exam|4187,4191|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Anatomy|Body Part, Organ, or Organ Component|General Exam|4187,4191|false|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|HEAD
Disorder|Disease or Syndrome|General Exam|4187,4191|false|false|false|C0362076|Problems with head|HEAD
Event|Event|General Exam|4187,4191|false|false|false|||HEAD
Procedure|Therapeutic or Preventive Procedure|General Exam|4187,4191|false|false|false|C0876917|Procedure on head|HEAD
Event|Event|General Exam|4196,4204|true|false|false|||evidence
Finding|Idea or Concept|General Exam|4196,4204|true|false|false|C3887511|Evidence|evidence
Finding|Functional Concept|General Exam|4196,4207|true|false|false|C0332120|Evidence of (contextual qualifier)|evidence of
Finding|Intellectual Product|General Exam|4208,4213|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Anatomy|Body Location or Region|General Exam|4214,4226|true|false|false|C0524466|Intracranial|intracranial
Finding|Functional Concept|General Exam|4214,4226|true|false|false|C1522213|Intracranial Route of Administration|intracranial
Anatomy|Body Part, Organ, or Organ Component|General Exam|4227,4234|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|4227,4234|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|General Exam|4227,4234|true|false|false|||process
Finding|Functional Concept|General Exam|4227,4234|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|4227,4234|true|false|false|C1522240|Process|process
Finding|Functional Concept|General Exam|4240,4244|false|false|false|C1552822|Table Cell Horizontal Align - left|left
Anatomy|Body Part, Organ, or Organ Component|General Exam|4240,4259|false|false|false|C0925567|Left zygomatic arch|left zygomatic arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|4245,4259|false|false|false|C0162485|Zygomatic Arch|zygomatic arch
Anatomy|Body Location or Region|General Exam|4255,4259|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Part, Organ, or Organ Component|General Exam|4255,4259|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Anatomy|Body Space or Junction|General Exam|4255,4259|false|false|false|C0003741;C0230467;C0741204|ARCH;Arch of foot;Structure of nucleus infundibularis hypothalami|arch
Finding|Finding|General Exam|4255,4259|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Finding|Gene or Genome|General Exam|4255,4259|false|false|false|C1538146;C4722404|Age-Related Clonal Hematopoiesis;ZBTB8OS gene|arch
Disorder|Anatomical Abnormality|General Exam|4260,4269|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Disorder|Congenital Abnormality|General Exam|4260,4269|false|false|false|C0000768;C0302142|Congenital Abnormality;Deformity|deformity
Event|Event|General Exam|4260,4269|false|false|false|||deformity
Finding|Finding|General Exam|4260,4269|false|false|false|C2117111||deformity
Finding|Finding|General Exam|4273,4281|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Finding|Idea or Concept|General Exam|4273,4281|true|false|false|C0332148;C0750492|Probable diagnosis;Probably|probably
Event|Event|General Exam|4282,4289|true|false|false|||chronic
Finding|Intellectual Product|General Exam|4282,4289|true|false|false|C1547296|Chronic - Admission Level of Care Code|chronic
Procedure|Health Care Activity|General Exam|4282,4289|true|false|false|C1555457|Provision of recurring care for chronic illness|chronic
Disorder|Disease or Syndrome|General Exam|4317,4321|true|false|false|C3542022|Short stature, onychodysplasia, facial dysmorphism, hypotrichosis syndrome|soft
Anatomy|Body Location or Region|General Exam|4317,4328|true|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Anatomy|Tissue|General Exam|4317,4328|true|false|false|C0225317;C4532079|Neck+Chest>Soft tissue;soft tissue|soft tissue
Disorder|Disease or Syndrome|General Exam|4317,4337|true|false|false|C0037580|Soft tissue swelling|soft tissue swelling
Anatomy|Tissue|General Exam|4322,4328|true|false|false|C0040300|Body tissue|tissue
Finding|Intellectual Product|General Exam|4322,4328|true|false|false|C1547928|Tissue Specimen Code|tissue
Event|Event|General Exam|4329,4337|true|false|false|||swelling
Finding|Finding|General Exam|4329,4337|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Finding|Pathologic Function|General Exam|4329,4337|true|false|false|C0013604;C0038999|Edema;Swelling|swelling
Event|Event|General Exam|4344,4347|false|false|false|||CXR
Procedure|Diagnostic Procedure|General Exam|4344,4347|false|false|false|C0039985|Plain chest X-ray|CXR
Finding|Intellectual Product|General Exam|4352,4357|true|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|acute
Event|Event|General Exam|4358,4371|true|false|false|||intrathoracic
Finding|Functional Concept|General Exam|4358,4371|true|false|false|C0595836|Intrathoracic Route of Administration|intrathoracic
Anatomy|Body Part, Organ, or Organ Component|General Exam|4372,4379|true|false|false|C1184743|bony process|process
Drug|Pharmacologic Substance|General Exam|4372,4379|true|false|false|C1951340|Process Pharmacologic Substance|process
Event|Event|General Exam|4372,4379|true|false|false|||process
Finding|Functional Concept|General Exam|4372,4379|true|false|false|C4521054|Process (qualifier value)|process
Phenomenon|Phenomenon or Process|General Exam|4372,4379|true|false|false|C1522240|Process|process
Finding|Body Substance|General Exam|4382,4391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Intellectual Product|General Exam|4382,4391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Finding|Sign or Symptom|General Exam|4382,4391|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|DISCHARGE
Procedure|Health Care Activity|General Exam|4382,4391|false|false|false|C0030685|Patient Discharge|DISCHARGE
Event|Event|General Exam|4392,4396|false|false|false|||LABS
Lab|Laboratory or Test Result|General Exam|4392,4396|false|false|false|C0587081|Laboratory test finding|LABS
Disorder|Disease or Syndrome|General Exam|4426,4431|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4426,4431|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4426,4431|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Anatomy|Cell|General Exam|4432,4435|false|false|false|C0023516|Leukocytes|WBC
Anatomy|Cell|General Exam|4440,4443|false|false|false|C0014792|Erythrocytes|RBC
Attribute|Clinical Attribute|General Exam|4440,4443|false|false|false|C1114281||RBC
Drug|Pharmacologic Substance|General Exam|4440,4443|false|false|false|C0014792|Erythrocytes|RBC
Drug|Amino Acid, Peptide, or Protein|General Exam|4450,4453|false|false|false|C0019046|Hemoglobin|Hgb
Drug|Biologically Active Substance|General Exam|4450,4453|false|false|false|C0019046|Hemoglobin|Hgb
Finding|Gene or Genome|General Exam|4450,4453|false|false|false|C1424337|CYGB gene|Hgb
Lab|Laboratory or Test Result|General Exam|4450,4453|false|false|false|C0019029|Hemoglobin concentration|Hgb
Procedure|Laboratory Procedure|General Exam|4460,4463|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Procedure|Therapeutic or Preventive Procedure|General Exam|4460,4463|false|false|false|C0018935;C0472699|Hematocrit Measurement;Hemopoietic stem cell transplant|Hct
Disorder|Virus|General Exam|4471,4474|false|false|false|C2304881|Merkel cell polyomavirus|MCV
Event|Event|General Exam|4471,4474|false|false|false|||MCV
Lab|Laboratory or Test Result|General Exam|4471,4474|false|false|false|C0524587|Mean Corpuscular Volume|MCV
Procedure|Laboratory Procedure|General Exam|4471,4474|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Procedure|Therapeutic or Preventive Procedure|General Exam|4471,4474|false|false|false|C0285131;C1948043|Cisplatin-Methotrexate-Vinblastine Regimen;Erythrocyte Mean Corpuscular Volume Measurement|MCV
Drug|Organic Chemical|General Exam|4480,4483|false|false|false|C0600370|methacholine|MCH
Drug|Pharmacologic Substance|General Exam|4480,4483|false|false|false|C0600370|methacholine|MCH
Event|Event|General Exam|4480,4483|false|false|false|||MCH
Finding|Gene or Genome|General Exam|4480,4483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Finding|Molecular Function|General Exam|4480,4483|false|false|false|C1418669;C2248810|PMCH gene;mesaconyl-CoA hydratase activity|MCH
Procedure|Laboratory Procedure|General Exam|4480,4483|false|false|false|C0369183|Mean corpuscular hemoglobin determination|MCH
Procedure|Laboratory Procedure|General Exam|4490,4494|false|false|false|C0474535|Mean corpuscular hemoglobin concentration determination|MCHC
Event|Event|General Exam|4500,4503|false|false|false|||RDW
Procedure|Laboratory Procedure|General Exam|4510,4513|false|false|false|C0201617|Primed lymphocyte test|Plt
Disorder|Disease or Syndrome|General Exam|4533,4538|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4533,4538|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4533,4538|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4543,4546|false|false|false|C2959585|Proliferating trichilemmal tumor|PTT
Event|Event|General Exam|4543,4546|false|false|false|||PTT
Procedure|Laboratory Procedure|General Exam|4543,4546|false|false|false|C0030605;C5552692|Partial Thromboplastin Time;Partial thromboplastin time, activated (procedure)|PTT
Disorder|Disease or Syndrome|General Exam|4569,4574|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4569,4574|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4569,4574|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Drug|Organic Chemical|General Exam|4569,4582|false|false|false|C0005802|Blood Glucose|BLOOD Glucose
Lab|Laboratory or Test Result|General Exam|4569,4582|false|false|false|C0428554|Finding of blood glucose level|BLOOD Glucose
Procedure|Laboratory Procedure|General Exam|4569,4582|false|false|false|C0392201|Blood glucose measurement|BLOOD Glucose
Drug|Biologically Active Substance|General Exam|4575,4582|false|false|false|C0017725|glucose|Glucose
Drug|Organic Chemical|General Exam|4575,4582|false|false|false|C0017725|glucose|Glucose
Drug|Pharmacologic Substance|General Exam|4575,4582|false|false|false|C0017725|glucose|Glucose
Event|Event|General Exam|4575,4582|false|false|false|||Glucose
Lab|Laboratory or Test Result|General Exam|4575,4582|false|false|false|C5781949|Glucose^1.5H post dose glucagon|Glucose
Procedure|Laboratory Procedure|General Exam|4575,4582|false|false|false|C0337438|Glucose measurement|Glucose
Event|Event|General Exam|4619,4620|false|false|false|||5
Drug|Inorganic Chemical|General Exam|4630,4634|false|false|false|C0005367|Bicarbonates|HCO3
Drug|Pharmacologic Substance|General Exam|4630,4634|false|false|false|C0005367|Bicarbonates|HCO3
Procedure|Laboratory Procedure|General Exam|4630,4634|false|false|false|C0202059|Bicarbonate measurement|HCO3
Disorder|Disease or Syndrome|General Exam|4659,4664|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4659,4664|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4659,4664|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Disorder|Neoplastic Process|General Exam|4665,4668|false|false|false|C1266129;C1370889|Atypical Lipoma;Liposarcoma, well differentiated|ALT
Drug|Amino Acid, Peptide, or Protein|General Exam|4665,4668|false|false|false|C0001899|Alanine Transaminase|ALT
Drug|Enzyme|General Exam|4665,4668|false|false|false|C0001899|Alanine Transaminase|ALT
Event|Event|General Exam|4665,4668|false|false|false|||ALT
Finding|Gene or Genome|General Exam|4665,4668|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Intellectual Product|General Exam|4665,4668|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Finding|Molecular Function|General Exam|4665,4668|false|false|false|C1140170;C1415274;C2257651|Alternative Billing Concepts;GPT gene|ALT
Procedure|Therapeutic or Preventive Procedure|General Exam|4665,4668|false|false|false|C4553172|Antibiotic Lock Therapy|ALT
Anatomy|Body Space or Junction|General Exam|4673,4676|false|false|false|C1185650|Asterion|AST
Disorder|Neoplastic Process|General Exam|4673,4676|false|false|false|C4522245|Atypical Spitz Nevus|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4673,4676|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Biologically Active Substance|General Exam|4673,4676|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Drug|Enzyme|General Exam|4673,4676|false|false|false|C0004002;C0242192;C1121182|Aspartate Transaminase;SGOT - Glutamate oxaloacetate transaminase;SLC17A5 protein, human|AST
Event|Event|General Exam|4673,4676|false|false|false|||AST
Finding|Gene or Genome|General Exam|4673,4676|false|false|false|C1415181;C1420113;C5960784|GOT1 gene;SLC17A5 gene;SLC17A5 wt Allele|AST
Drug|Amino Acid, Peptide, or Protein|General Exam|4682,4689|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Drug|Enzyme|General Exam|4682,4689|false|false|false|C0002059|Alkaline Phosphatase|AlkPhos
Disorder|Disease or Syndrome|General Exam|4718,4723|false|false|false|C0851353|Blood and lymphatic system disorders|BLOOD
Event|Event|General Exam|4718,4723|false|false|false|||BLOOD
Finding|Body Substance|General Exam|4718,4723|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|BLOOD
Procedure|Laboratory Procedure|General Exam|4718,4731|false|false|false|C0729820|Blood calcium measurement|BLOOD Calcium
Drug|Biologically Active Substance|General Exam|4724,4731|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|4724,4731|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|4724,4731|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|4724,4731|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|4724,4731|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|4724,4731|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|4724,4731|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|4724,4731|false|false|false|C0201925|Calcium measurement|Calcium
Disorder|Disease or Syndrome|General Exam|4758,4761|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|4758,4761|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|4758,4761|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|4758,4761|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|4758,4761|false|false|false|||HIV
Event|Event|General Exam|4765,4770|false|false|false|||HAART
Procedure|Therapeutic or Preventive Procedure|General Exam|4765,4770|false|false|false|C0887947|Antiretroviral Therapy, Highly Active|HAART
Disorder|Disease or Syndrome|General Exam|4772,4776|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|4772,4776|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|4772,4776|false|false|false|||COPD
Finding|Gene or Genome|General Exam|4772,4776|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|General Exam|4783,4787|false|false|false|||home
Finding|Idea or Concept|General Exam|4783,4787|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|4783,4787|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|4783,4787|false|false|false|C1553498|home health encounter|home
Disorder|Disease or Syndrome|General Exam|4792,4795|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|General Exam|4792,4795|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Disease or Syndrome|General Exam|4796,4805|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|General Exam|4796,4805|false|false|false|||cirrhosis
Disorder|Disease or Syndrome|General Exam|4822,4829|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|4822,4829|false|false|false|||ascites
Finding|Pathologic Function|General Exam|4822,4829|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|General Exam|4830,4839|false|false|false|||requiring
Drug|Organic Chemical|General Exam|4849,4860|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|General Exam|4849,4860|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|General Exam|4849,4860|false|false|false|||therapeutic
Finding|Functional Concept|General Exam|4849,4860|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|General Exam|4849,4860|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|General Exam|4849,4860|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|General Exam|4862,4874|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|4862,4874|false|false|false|C0034115|Paracentesis|paracenteses
Anatomy|Body Location or Region|General Exam|4876,4883|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|General Exam|4876,4898|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|General Exam|4884,4898|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|General Exam|4884,4898|false|false|false|||encephalopathy
Anatomy|Tissue|General Exam|4907,4917|true|false|false|C0332835|Transplanted tissue|transplant
Finding|Finding|General Exam|4907,4917|true|false|false|C0478647;C3841811|Transplant;Transplanted organ and tissue status|transplant
Procedure|Therapeutic or Preventive Procedure|General Exam|4907,4917|true|false|false|C0040732|Transplantation|transplant
Event|Event|General Exam|4918,4922|true|false|false|||list
Finding|Intellectual Product|General Exam|4918,4922|true|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|General Exam|4928,4941|false|false|false|||comorbidities
Finding|Finding|General Exam|4928,4941|false|false|false|C0009488|Comorbidity|comorbidities
Disorder|Disease or Syndrome|General Exam|4946,4949|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Event|Event|General Exam|4946,4949|false|false|false|||AMS
Finding|Gene or Genome|General Exam|4946,4949|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|General Exam|4946,4949|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Event|Event|General Exam|4951,4962|false|false|false|||hypotension
Finding|Finding|General Exam|4951,4962|false|false|false|C0020649|Hypotension|hypotension
Event|Event|General Exam|4973,4985|false|false|false|||hyperkalemia
Finding|Finding|General Exam|4973,4985|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Finding|Mental Process|General Exam|4996,5002|false|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|General Exam|4996,5009|false|false|false|C0488568;C0488569||mental status
Finding|Finding|General Exam|4996,5009|false|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|General Exam|5003,5009|false|false|false|C5889824||status
Event|Event|General Exam|5003,5009|false|false|false|||status
Finding|Idea or Concept|General Exam|5003,5009|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|5010,5018|false|false|false|||improved
Drug|Organic Chemical|General Exam|5024,5033|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|General Exam|5024,5033|false|false|false|C0022957|lactulose|lactulose
Event|Event|General Exam|5024,5033|false|false|false|||lactulose
Event|Event|General Exam|5035,5046|false|false|false|||Hypotension
Finding|Finding|General Exam|5035,5046|false|false|false|C0020649|Hypotension|Hypotension
Event|Event|General Exam|5052,5056|false|false|false|||felt
Drug|Substance|General Exam|5070,5075|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Event|Event|General Exam|5070,5075|false|false|false|||fluid
Finding|Intellectual Product|General Exam|5070,5075|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Physiologic Function|General Exam|5070,5082|false|false|false|C0242705|Fluid Shifts|fluid shifts
Event|Event|General Exam|5076,5082|false|false|false|||shifts
Finding|Functional Concept|General Exam|5076,5082|false|false|false|C0333051|shift displacement|shifts
Event|Event|General Exam|5088,5100|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|General Exam|5088,5100|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Idea or Concept|General Exam|5108,5111|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|General Exam|5108,5111|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|General Exam|5122,5131|false|false|false|||admission
Procedure|Health Care Activity|General Exam|5122,5131|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|General Exam|5135,5139|false|false|false|C5575035|Well (answer to question)|well
Finding|Finding|General Exam|5143,5146|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|5143,5146|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Event|Event|General Exam|5150,5156|false|false|false|||intake
Finding|Functional Concept|General Exam|5150,5156|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|General Exam|5150,5156|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Finding|Mental Process|General Exam|5164,5171|false|false|false|C0542559|contextual factors|setting
Disorder|Disease or Syndrome|General Exam|5176,5179|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Event|Event|General Exam|5176,5179|false|false|false|||AMS
Finding|Gene or Genome|General Exam|5176,5179|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|General Exam|5176,5179|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Event|Event|General Exam|5181,5192|false|false|false|||Hypotension
Finding|Finding|General Exam|5181,5192|false|false|false|C0020649|Hypotension|Hypotension
Event|Event|General Exam|5201,5209|false|false|false|||resolved
Drug|Amino Acid, Peptide, or Protein|General Exam|5218,5225|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|General Exam|5218,5225|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|General Exam|5218,5225|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|General Exam|5218,5225|false|false|false|||albumin
Finding|Gene or Genome|General Exam|5218,5225|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|General Exam|5218,5225|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|General Exam|5218,5225|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|General Exam|5227,5239|false|false|false|||Hyperkalemia
Finding|Finding|General Exam|5227,5239|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Event|Event|General Exam|5241,5249|false|false|false|||resolved
Drug|Amino Acid, Peptide, or Protein|General Exam|5255,5262|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|General Exam|5255,5262|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|General Exam|5255,5262|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|General Exam|5255,5262|false|false|false|||insulin
Finding|Gene or Genome|General Exam|5255,5262|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|General Exam|5255,5262|false|false|false|C0202098|Insulin measurement|insulin
Drug|Organic Chemical|General Exam|5267,5277|false|false|false|C0124498|Kayexalate|kayexalate
Drug|Pharmacologic Substance|General Exam|5267,5277|false|false|false|C0124498|Kayexalate|kayexalate
Event|Event|General Exam|5267,5277|false|false|false|||kayexalate
Event|Event|General Exam|5282,5293|false|false|false|||Hypotension
Finding|Finding|General Exam|5282,5293|false|false|false|C0020649|Hypotension|Hypotension
Finding|Body Substance|General Exam|5295,5302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|5295,5302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|5295,5302|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|5303,5312|false|false|false|||presented
Attribute|Clinical Attribute|General Exam|5318,5321|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|General Exam|5318,5321|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|General Exam|5318,5321|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|General Exam|5318,5321|false|false|false|||SBP
Finding|Gene or Genome|General Exam|5318,5321|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|General Exam|5318,5321|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|General Exam|5333,5341|false|false|false|||improved
Finding|Finding|General Exam|5333,5341|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Finding|Intellectual Product|General Exam|5333,5341|false|false|false|C0184511;C1561611;C4084203|Admission Level of Care Code - Improved;Improved;Improved - answer to question|improved
Drug|Amino Acid, Peptide, or Protein|General Exam|5348,5355|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|General Exam|5348,5355|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|General Exam|5348,5355|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|General Exam|5348,5355|false|false|false|||albumin
Finding|Gene or Genome|General Exam|5348,5355|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|General Exam|5348,5355|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|General Exam|5348,5355|false|false|false|C0201838|Albumin measurement|albumin
Event|Event|General Exam|5381,5385|false|false|false|||felt
Drug|Substance|General Exam|5400,5405|false|false|false|C0302908;C1704353|Liquid substance;fluid - substance|fluid
Finding|Intellectual Product|General Exam|5400,5405|false|false|false|C1546638|Fluid Specimen Code|fluid
Finding|Physiologic Function|General Exam|5400,5412|false|false|false|C0242705|Fluid Shifts|fluid shifts
Event|Event|General Exam|5406,5412|false|false|false|||shifts
Finding|Functional Concept|General Exam|5406,5412|false|false|false|C0333051|shift displacement|shifts
Event|Event|General Exam|5418,5430|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|General Exam|5418,5430|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Finding|General Exam|5442,5446|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|5450,5456|false|false|false|||likely
Finding|Finding|General Exam|5450,5456|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5450,5456|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|General Exam|5458,5469|false|false|false|C0546884|Hypovolemia|hypovolemia
Disorder|Disease or Syndrome|General Exam|5476,5479|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Event|Event|General Exam|5476,5479|false|false|false|||AMS
Finding|Gene or Genome|General Exam|5476,5479|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|General Exam|5476,5479|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Event|Event|General Exam|5484,5493|false|false|false|||decreased
Finding|Finding|General Exam|5484,5503|false|false|false|C1504561|Hypophagia|decreased PO intake
Event|Event|General Exam|5497,5503|false|false|false|||intake
Finding|Functional Concept|General Exam|5497,5503|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|General Exam|5497,5503|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Event|Event|General Exam|5508,5515|true|false|false|||concern
Finding|Idea or Concept|General Exam|5508,5515|true|false|false|C2699424|Concern|concern
Event|Event|General Exam|5521,5529|true|false|false|||bleeding
Finding|Pathologic Function|General Exam|5521,5529|true|false|false|C0019080|Hemorrhage|bleeding
Disorder|Disease or Syndrome|General Exam|5533,5539|true|false|false|C0036690;C0243026|Sepsis;Septicemia|sepsis
Event|Event|General Exam|5533,5539|true|false|false|||sepsis
Drug|Biomedical or Dental Material|General Exam|5545,5553|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|5545,5553|false|false|false|||baseline
Finding|Idea or Concept|General Exam|5545,5553|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Anatomy|Cell Component|General Exam|5554,5557|false|false|false|C2263086|Nuclear cap binding complex location|CBC
Event|Event|General Exam|5554,5557|false|false|false|||CBC
Procedure|Laboratory Procedure|General Exam|5554,5557|false|false|false|C0009555|Complete Blood Count|CBC
Event|Event|General Exam|5570,5575|false|false|false|||fever
Finding|Finding|General Exam|5570,5575|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Finding|Sign or Symptom|General Exam|5570,5575|false|false|false|C0015967;C0424755|Fever;Fever symptoms (finding)|fever
Event|Event|General Exam|5582,5591|false|false|false|||continued
Event|Event|General Exam|5595,5603|false|false|false|||received
Drug|Amino Acid, Peptide, or Protein|General Exam|5607,5614|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|General Exam|5607,5614|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|General Exam|5607,5614|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|General Exam|5607,5614|false|false|false|||albumin
Finding|Gene or Genome|General Exam|5607,5614|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|General Exam|5607,5614|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|General Exam|5607,5614|false|false|false|C0201838|Albumin measurement|albumin
Finding|Idea or Concept|General Exam|5626,5634|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|General Exam|5626,5641|false|false|false|C0488549||hospital course
Finding|Finding|General Exam|5626,5641|false|false|false|C0489547|Hospital course|hospital course
Event|Event|General Exam|5635,5641|false|false|false|||course
Attribute|Clinical Attribute|General Exam|5659,5662|false|false|false|C0871470|Systolic Pressure|SBP
Drug|Amino Acid, Peptide, or Protein|General Exam|5659,5662|false|false|false|C0085805|Androgen Binding Protein|SBP
Drug|Biologically Active Substance|General Exam|5659,5662|false|false|false|C0085805|Androgen Binding Protein|SBP
Event|Event|General Exam|5659,5662|false|false|false|||SBP
Finding|Gene or Genome|General Exam|5659,5662|false|false|false|C1705296;C3274833|CCHCR1 wt Allele;SHBG wt Allele|SBP
Procedure|Diagnostic Procedure|General Exam|5659,5662|false|false|false|C1306620|Systolic blood pressure measurement|SBP
Event|Event|General Exam|5663,5671|false|false|false|||improved
Finding|Body Substance|General Exam|5683,5690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|5683,5690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|5683,5690|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|5691,5699|false|false|false|||remained
Event|Event|General Exam|5701,5713|false|false|false|||asymptomatic
Finding|Finding|General Exam|5701,5713|false|false|false|C0231221;C0332151|Asymptomatic (finding);Asymptomatic diagnosis of|asymptomatic
Event|Event|General Exam|5720,5732|false|false|false|||Hyperkalemia
Finding|Finding|General Exam|5720,5732|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Finding|Body Substance|General Exam|5734,5741|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|5734,5741|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|5734,5741|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|5742,5751|false|false|false|||presented
Event|Event|General Exam|5768,5771|false|false|false|||EKG
Finding|Intellectual Product|General Exam|5768,5771|false|false|false|C0013798;C5945056|Electrocardiogram;Electrocardiogram image|EKG
Procedure|Diagnostic Procedure|General Exam|5768,5771|false|false|false|C1623258|Electrocardiography|EKG
Event|Event|General Exam|5772,5779|false|false|false|||changes
Finding|Functional Concept|General Exam|5772,5779|false|false|false|C0392747|Changing|changes
Finding|Finding|General Exam|5788,5791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|5788,5791|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|General Exam|5796,5802|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5796,5802|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Finding|General Exam|5807,5813|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Functional Concept|General Exam|5807,5813|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Idea or Concept|General Exam|5807,5813|false|false|false|C1274040;C1546471;C2825142|Experimental Result;Result;What subject filter - Result|result
Finding|Finding|General Exam|5817,5820|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|5817,5820|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Part, Organ, or Organ Component|General Exam|5831,5839|false|false|false|C0003842|Arteries|arterial
Event|Event|General Exam|5840,5846|false|false|false|||volume
Finding|Intellectual Product|General Exam|5840,5846|false|false|false|C1705102|Volume (publication)|volume
Event|Event|General Exam|5848,5855|false|false|false|||leading
Finding|Intellectual Product|General Exam|5859,5863|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|General Exam|5866,5875|false|false|false|||excretion
Finding|Body Substance|General Exam|5866,5875|false|false|false|C0221102;C0504085|Body Excretions;Excretory function|excretion
Finding|Physiologic Function|General Exam|5866,5875|false|false|false|C0221102;C0504085|Body Excretions;Excretory function|excretion
Finding|Finding|General Exam|5882,5888|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|5882,5888|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|5889,5901|false|false|false|||exacerbation
Finding|Finding|General Exam|5889,5901|false|true|false|C4086268|Exacerbation|exacerbation
Drug|Hormone|General Exam|5916,5924|false|false|false|C0020268|hydrocortisone|cortisol
Drug|Organic Chemical|General Exam|5916,5924|false|false|false|C0020268|hydrocortisone|cortisol
Drug|Pharmacologic Substance|General Exam|5916,5924|false|false|false|C0020268|hydrocortisone|cortisol
Event|Event|General Exam|5916,5924|false|false|false|||cortisol
Procedure|Laboratory Procedure|General Exam|5916,5924|false|false|false|C0201968|Cortisol Measurement|cortisol
Event|Event|General Exam|5929,5935|false|false|false|||normal
Event|Event|General Exam|5939,5947|false|false|false|||improved
Drug|Amino Acid, Peptide, or Protein|General Exam|5953,5960|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Hormone|General Exam|5953,5960|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Drug|Pharmacologic Substance|General Exam|5953,5960|false|false|false|C0021641;C0795635;C1533581;C1579433;C3714501;C4721402|INS protein, human;Insulin;Insulin Drug Class;Insulin [EPC];Therapeutic Insulin;insulin, regular, human|insulin
Event|Event|General Exam|5953,5960|false|false|false|||insulin
Finding|Gene or Genome|General Exam|5953,5960|false|false|false|C1337112|INS gene|insulin
Procedure|Laboratory Procedure|General Exam|5953,5960|false|false|false|C0202098|Insulin measurement|insulin
Drug|Organic Chemical|General Exam|5965,5975|false|false|false|C0124498|Kayexalate|kayexalate
Drug|Pharmacologic Substance|General Exam|5965,5975|false|false|false|C0124498|Kayexalate|kayexalate
Event|Event|General Exam|5965,5975|false|false|false|||kayexalate
Finding|Idea or Concept|General Exam|5994,5997|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|General Exam|5994,5997|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|General Exam|6001,6010|false|false|false|||discharge
Finding|Body Substance|General Exam|6001,6010|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|6001,6010|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|6001,6010|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|6001,6010|false|false|false|C0030685|Patient Discharge|discharge
Drug|Organic Chemical|General Exam|6012,6019|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|General Exam|6012,6019|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|General Exam|6024,6028|false|false|false|||held
Finding|Idea or Concept|General Exam|6037,6045|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|General Exam|6037,6052|false|false|false|C0488549||hospital course
Finding|Finding|General Exam|6037,6052|false|false|false|C0489547|Hospital course|hospital course
Event|Event|General Exam|6046,6052|false|false|false|||course
Finding|Body Substance|General Exam|6063,6070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|6063,6070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|6063,6070|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|6071,6080|false|false|false|||presented
Drug|Biomedical or Dental Material|General Exam|6098,6106|false|false|false|C0168634|BaseLine dental cement|baseline
Event|Event|General Exam|6098,6106|false|false|false|||baseline
Finding|Idea or Concept|General Exam|6098,6106|false|false|false|C1552824|baseline - TableCellVerticalAlign|baseline
Event|Event|General Exam|6130,6134|false|false|false|||felt
Event|Event|General Exam|6141,6147|false|false|false|||likely
Finding|Finding|General Exam|6141,6147|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|6141,6147|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Event|Event|General Exam|6155,6161|false|false|false|||volume
Finding|Intellectual Product|General Exam|6155,6161|false|true|false|C1705102|Volume (publication)|volume
Event|Event|General Exam|6162,6167|false|false|false|||shift
Finding|Functional Concept|General Exam|6162,6167|false|true|false|C0333051|shift displacement|shift
Phenomenon|Phenomenon or Process|General Exam|6162,6167|false|true|false|C2347509|Physical Shift|shift
Event|Event|General Exam|6178,6190|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|General Exam|6178,6190|false|false|false|C0034115|Paracentesis|paracentesis
Finding|Idea or Concept|General Exam|6198,6201|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Finding|Intellectual Product|General Exam|6198,6201|false|false|false|C1561538;C1561539|Precision - day;Transaction counts and value totals - day|day
Event|Event|General Exam|6211,6220|false|false|false|||admission
Procedure|Health Care Activity|General Exam|6211,6220|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Finding|Finding|General Exam|6224,6228|false|false|false|C5575035|Well (answer to question)|well
Event|Event|General Exam|6236,6239|false|false|false|||low
Finding|Finding|General Exam|6236,6239|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|6236,6239|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Anatomy|Body Part, Organ, or Organ Component|General Exam|6251,6259|false|false|false|C0003842|Arteries|arterial
Event|Event|General Exam|6260,6266|false|false|false|||volume
Finding|Intellectual Product|General Exam|6260,6266|false|false|false|C1705102|Volume (publication)|volume
Finding|Finding|General Exam|6268,6274|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|6268,6274|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Intellectual Product|General Exam|6279,6283|false|false|false|C1547310;C4723750|International Metastatic Renal Cell Carcinoma Database Consortium (IMDC) Criteria - Poor-Risk Group;Patient Condition Code - Poor|poor
Event|Event|General Exam|6287,6293|false|false|false|||intake
Finding|Functional Concept|General Exam|6287,6293|false|false|false|C1512806|Intake|intake
Procedure|Health Care Activity|General Exam|6287,6293|false|false|false|C3251814;C4521161|Intake (treatment);Measurement of fluid intake|intake
Disorder|Disease or Syndrome|General Exam|6298,6301|false|false|false|C1860224|ABLEPHARON-MACROSTOMIA SYNDROME|AMS
Event|Event|General Exam|6298,6301|false|false|false|||AMS
Finding|Gene or Genome|General Exam|6298,6301|false|false|false|C4284022|TWIST2 wt Allele|AMS
Procedure|Laboratory Procedure|General Exam|6298,6301|false|false|false|C4521393|Accelerator Mass Spectrometry|AMS
Event|Event|General Exam|6307,6315|false|false|false|||improved
Drug|Amino Acid, Peptide, or Protein|General Exam|6328,6335|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Biologically Active Substance|General Exam|6328,6335|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Drug|Pharmacologic Substance|General Exam|6328,6335|false|false|false|C0001924;C5966160|Albumin;Albumins|albumin
Event|Event|General Exam|6328,6335|false|false|false|||albumin
Finding|Gene or Genome|General Exam|6328,6335|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Finding|Physiologic Function|General Exam|6328,6335|false|false|false|C1412332;C4553023|ALB gene;Albumin metabolic function|albumin
Procedure|Laboratory Procedure|General Exam|6328,6335|false|false|false|C0201838|Albumin measurement|albumin
Procedure|Therapeutic or Preventive Procedure|General Exam|6328,6350|false|false|false|C1293861|Administration of albumin|albumin administration
Event|Event|General Exam|6336,6350|false|false|false|||administration
Event|Occupational Activity|General Exam|6336,6350|false|false|false|C0001554|Administration occupational activities|administration
Procedure|Therapeutic or Preventive Procedure|General Exam|6336,6350|false|false|false|C1533734|Administration (procedure)|administration
Drug|Organic Chemical|General Exam|6352,6362|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|General Exam|6352,6362|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|General Exam|6368,6375|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|General Exam|6368,6375|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|General Exam|6381,6385|false|false|false|||held
Finding|Idea or Concept|General Exam|6393,6401|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|General Exam|6393,6408|false|false|false|C0488549||hospital course
Finding|Finding|General Exam|6393,6408|false|false|false|C0489547|Hospital course|hospital course
Event|Event|General Exam|6402,6408|false|false|false|||course
Disorder|Anatomical Abnormality|General Exam|6415,6418|false|false|false|C0399558|Glandular odontogenic cyst|GOC
Event|Event|General Exam|6415,6418|false|false|false|||GOC
Finding|Gene or Genome|General Exam|6428,6431|false|false|false|C1420310|SON gene|son
Disorder|Disease or Syndrome|General Exam|6433,6436|false|false|false|C0162531|Hereditary Coproporphyria|HCP
Event|Event|General Exam|6433,6436|false|false|false|||HCP
Finding|Gene or Genome|General Exam|6433,6436|false|false|false|C1335283;C1412376;C1413681;C1705637;C5780748|AMBP gene;AMBP wt Allele;CPOX gene;PTPN6 gene;PTPN6 wt Allele|HCP
Event|Event|General Exam|6438,6441|false|false|false|||met
Finding|Classification|General Exam|6456,6466|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|6456,6466|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|General Exam|6467,6479|false|false|false|||hepatologist
Finding|Idea or Concept|General Exam|6492,6500|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|General Exam|6492,6507|false|false|false|C0488549||hospital course
Finding|Finding|General Exam|6492,6507|false|false|false|C0489547|Hospital course|hospital course
Event|Event|General Exam|6501,6507|false|false|false|||course
Event|Event|General Exam|6515,6524|true|false|false|||discussed
Finding|Body Substance|General Exam|6534,6541|true|false|true|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6534,6541|true|false|true|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6534,6541|true|false|true|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Anatomy|Tissue|General Exam|6551,6561|true|false|false|C0332835|Transplanted tissue|transplant
Finding|Finding|General Exam|6551,6561|true|false|false|C0478647;C3841811|Transplant;Transplanted organ and tissue status|transplant
Procedure|Therapeutic or Preventive Procedure|General Exam|6551,6561|true|false|false|C0040732|Transplantation|transplant
Event|Event|General Exam|6562,6571|true|false|false|||candidate
Finding|Conceptual Entity|General Exam|6562,6571|true|false|true|C4527371|Candidate|candidate
Finding|Finding|General Exam|6584,6594|true|false|false|C4722602|Underlying|underlying
Anatomy|Body Location or Region|General Exam|6595,6599|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Anatomy|Body Part, Organ, or Organ Component|General Exam|6595,6599|true|false|false|C0024109;C4037972|Chest>Lung;Lung|lung
Disorder|Disease or Syndrome|General Exam|6595,6599|true|false|false|C0024115|Lung diseases|lung
Finding|Finding|General Exam|6595,6599|true|false|false|C0740941|Lung Problem|lung
Disorder|Disease or Syndrome|General Exam|6595,6607|true|false|false|C0024115|Lung diseases|lung disease
Disorder|Disease or Syndrome|General Exam|6600,6607|false|false|false|C0012634|Disease|disease
Event|Event|General Exam|6600,6607|false|false|false|||disease
Attribute|Clinical Attribute|General Exam|6609,6613|false|false|false|C0802965||FEV1
Procedure|Diagnostic Procedure|General Exam|6609,6613|false|false|false|C0849974|Pulmonary Function Test/Forced Expiratory Volume 1|FEV1
Event|Event|General Exam|6621,6628|false|false|false|||hypoxia
Finding|Finding|General Exam|6621,6628|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Finding|Pathologic Function|General Exam|6621,6628|false|false|false|C0242184;C1963140|Hypoxia;Hypoxia, CTCAE|hypoxia
Event|Event|General Exam|6634,6642|false|false|false|||dilation
Finding|Finding|General Exam|6634,6642|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Finding|Pathologic Function|General Exam|6634,6642|false|false|false|C0012359;C0700124|Dilated;Pathological Dilatation|dilation
Procedure|Therapeutic or Preventive Procedure|General Exam|6634,6642|false|false|false|C1322279|Dilate procedure|dilation
Finding|Finding|General Exam|6647,6655|false|false|false|C0442811;C5202917|IPSS-R Risk Category Very Low;Very low (qualifier value)|very low
Finding|Finding|General Exam|6652,6655|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|General Exam|6652,6655|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Finding|General Exam|6652,6659|false|false|false|C5233331|Low BMI|low BMI
Attribute|Clinical Attribute|General Exam|6656,6659|false|false|false|C1305855;C1542867|Body mass index|BMI
Event|Event|General Exam|6656,6659|false|false|false|||BMI
Finding|Finding|General Exam|6656,6659|false|false|false|C0578022|Finding of body mass index|BMI
Finding|Functional Concept|General Exam|6681,6689|false|false|false|C5445118|Approach (contact)|approach
Event|Event|General Exam|6695,6706|false|false|false|||recommended
Finding|Body Substance|General Exam|6715,6722|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6715,6722|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6715,6722|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|6727,6739|false|false|false|||transitioned
Attribute|Clinical Attribute|General Exam|6743,6746|false|false|false|C4285234||DNR
Drug|Antibiotic|General Exam|6743,6746|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|General Exam|6743,6746|false|false|false|C0011015|daunorubicin|DNR
Event|Event|General Exam|6743,6746|false|false|false|||DNR
Finding|Finding|General Exam|6743,6746|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|General Exam|6743,6746|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Body Substance|General Exam|6757,6764|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6757,6764|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6757,6764|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|6765,6771|false|false|false|||agreed
Disorder|Disease or Syndrome|General Exam|6782,6786|false|false|false|C0270724|Infantile Neuroaxonal Dystrophy|plan
Event|Event|General Exam|6782,6786|false|false|false|||plan
Finding|Functional Concept|General Exam|6782,6786|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Intellectual Product|General Exam|6782,6786|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Finding|Mental Process|General Exam|6782,6786|false|false|false|C0032074;C0599880;C1301732|Planned;Treatment Plan|plan
Event|Event|General Exam|6796,6803|true|false|false|||treated
Event|Event|General Exam|6813,6817|true|false|false|||goal
Finding|Idea or Concept|General Exam|6813,6817|true|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Finding|Intellectual Product|General Exam|6813,6817|true|false|false|C0018017;C1571704|Act Mood - Goal;objective (goal)|goal
Event|Event|General Exam|6822,6830|true|false|false|||treating
Event|Event|General Exam|6851,6857|true|false|false|||issues
Finding|Functional Concept|General Exam|6859,6865|false|false|false|C0728831|Social|Social
Event|Occupational Activity|General Exam|6866,6870|false|false|false|C0043227|Work|work
Event|Event|General Exam|6871,6874|false|false|false|||met
Finding|Body Substance|General Exam|6885,6892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6885,6892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6885,6892|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|6902,6911|false|false|false|||discharge
Finding|Body Substance|General Exam|6902,6911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Intellectual Product|General Exam|6902,6911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Finding|Sign or Symptom|General Exam|6902,6911|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|discharge
Procedure|Health Care Activity|General Exam|6902,6911|false|false|false|C0030685|Patient Discharge|discharge
Finding|Body Substance|General Exam|6917,6924|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|6917,6924|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|6917,6924|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|6929,6939|false|false|false|||interested
Finding|Mental Process|General Exam|6929,6939|false|false|false|C0543488|Interested|interested
Event|Event|General Exam|6944,6953|false|false|false|||following
Finding|Finding|General Exam|6962,6977|false|false|false|C0700049|Encounter due to palliative care|palliative care
Procedure|Health Care Activity|General Exam|6962,6977|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|palliative care
Procedure|Therapeutic or Preventive Procedure|General Exam|6962,6977|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|palliative care
Event|Activity|General Exam|6973,6977|false|false|false|C1947933|care activity|care
Event|Event|General Exam|6973,6977|false|false|false|||care
Finding|Finding|General Exam|6973,6977|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|General Exam|6973,6977|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|General Exam|6992,7002|false|false|false|||outpatient
Finding|Classification|General Exam|6992,7002|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|6992,7002|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|General Exam|7004,7012|false|false|false|||referral
Procedure|Health Care Activity|General Exam|7004,7012|false|false|false|C0034927|Patient referral|referral
Event|Event|General Exam|7017,7021|false|false|false|||made
Finding|Mental Process|General Exam|7036,7042|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|7036,7049|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|General Exam|7036,7049|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|General Exam|7043,7049|false|false|false|C5889824||Status
Finding|Idea or Concept|General Exam|7043,7049|false|false|false|C1546481|What subject filter - Status|Status
Finding|Body Substance|General Exam|7051,7058|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|7051,7058|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|7051,7058|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|7059,7068|false|false|false|||presented
Disorder|Mental or Behavioral Dysfunction|General Exam|7074,7083|false|false|false|C0009676|Confusion|confusion
Event|Event|General Exam|7074,7083|false|false|false|||confusion
Finding|Finding|General Exam|7074,7083|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Idea or Concept|General Exam|7094,7105|false|false|false|C0750501|most likely|most likely
Finding|Finding|General Exam|7099,7105|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Finding|Idea or Concept|General Exam|7099,7105|false|false|false|C0332148;C0750492|Probable diagnosis;Probably|likely
Disorder|Neoplastic Process|General Exam|7106,7115|false|false|false|C0027627|Neoplasm Metastasis|secondary
Event|Event|General Exam|7106,7115|false|false|false|||secondary
Finding|Functional Concept|General Exam|7106,7115|false|false|false|C1522484|metastatic qualifier|secondary
Anatomy|Body Location or Region|General Exam|7119,7126|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|General Exam|7119,7141|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|General Exam|7127,7141|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|General Exam|7127,7141|false|false|false|||encephalopathy
Finding|Classification|General Exam|7153,7163|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|7153,7163|true|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|General Exam|7164,7171|true|false|false|||records
Finding|Idea or Concept|General Exam|7164,7171|true|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Intellectual Product|General Exam|7164,7171|true|false|false|C0034869;C1548330|Quantity limited request - Records;Records|records
Finding|Body Substance|General Exam|7173,7180|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|7173,7180|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|7173,7180|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Functional Concept|General Exam|7173,7184|false|false|false|C0332310|Has patient|patient has
Disorder|Disease or Syndrome|General Exam|7208,7231|true|false|false|C1619727|Decompensated cirrhosis of liver|decompensated cirrhosis
Disorder|Disease or Syndrome|General Exam|7222,7231|true|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|cirrhosis
Event|Event|General Exam|7222,7231|true|false|false|||cirrhosis
Finding|Mental Process|General Exam|7236,7242|true|false|false|C0229992|Psyche structure|mental
Attribute|Clinical Attribute|General Exam|7236,7249|true|false|false|C0488568;C0488569||mental status
Finding|Finding|General Exam|7236,7249|true|false|false|C0278060|Mental state|mental status
Attribute|Clinical Attribute|General Exam|7243,7249|true|false|false|C5889824||status
Event|Event|General Exam|7243,7249|true|false|false|||status
Finding|Idea or Concept|General Exam|7243,7249|true|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|7254,7259|true|false|false|||signs
Finding|Finding|General Exam|7254,7259|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Finding|Functional Concept|General Exam|7254,7259|true|false|false|C0220912;C0311392|Aspects of signs;Physical findings|signs
Disorder|Disease or Syndrome|General Exam|7263,7272|true|false|false|C0009450|Communicable Diseases|infection
Event|Event|General Exam|7263,7272|true|false|false|||infection
Finding|Pathologic Function|General Exam|7263,7272|true|false|false|C3714514|Infection|infection
Anatomy|Body Location or Region|General Exam|7278,7282|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Anatomy|Body Part, Organ, or Organ Component|General Exam|7278,7282|true|false|false|C0018670;C0152336|Head;Structure of head of caudate nucleus|head
Disorder|Disease or Syndrome|General Exam|7278,7282|true|false|false|C0362076|Problems with head|head
Procedure|Therapeutic or Preventive Procedure|General Exam|7278,7282|true|false|false|C0876917|Procedure on head|head
Procedure|Diagnostic Procedure|General Exam|7278,7285|true|false|false|C0202691|CAT scan of head|head CT
Event|Event|General Exam|7283,7285|true|false|false|||CT
Event|Event|General Exam|7290,7298|false|false|false|||negative
Finding|Classification|General Exam|7290,7298|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Finding|Finding|General Exam|7290,7298|false|false|false|C0205160;C1513916;C2699077|Negative;Negative Finding;Rh Negative Blood Group|negative
Lab|Laboratory or Test Result|General Exam|7290,7298|false|false|false|C5237010|Expression Negative|negative
Event|Event|General Exam|7302,7306|false|false|false|||well
Finding|Finding|General Exam|7302,7306|false|false|false|C5575035|Well (answer to question)|well
Finding|Mental Process|General Exam|7308,7314|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|General Exam|7308,7321|false|false|false|C0488568;C0488569||Mental status
Finding|Finding|General Exam|7308,7321|false|false|false|C0278060|Mental state|Mental status
Attribute|Clinical Attribute|General Exam|7315,7321|false|false|false|C5889824||status
Event|Event|General Exam|7315,7321|false|false|false|||status
Finding|Idea or Concept|General Exam|7315,7321|false|false|false|C1546481|What subject filter - Status|status
Event|Event|General Exam|7322,7330|false|false|false|||improved
Drug|Organic Chemical|General Exam|7337,7346|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|General Exam|7337,7346|false|false|false|C0022957|lactulose|lactulose
Event|Event|General Exam|7337,7346|false|false|false|||lactulose
Finding|Body Substance|General Exam|7361,7368|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|7361,7368|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|7361,7368|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|7369,7376|false|false|false|||reports
Drug|Organic Chemical|General Exam|7407,7416|true|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|General Exam|7407,7416|true|false|false|C0022957|lactulose|lactulose
Finding|Finding|General Exam|7427,7434|true|false|false|C4534363|At home|at home
Event|Event|General Exam|7430,7434|true|false|false|||home
Finding|Idea or Concept|General Exam|7430,7434|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|7430,7434|true|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|7430,7434|true|false|false|C1553498|home health encounter|home
Finding|Body Substance|General Exam|7436,7443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|7436,7443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|7436,7443|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|7453,7462|false|false|false|||continued
Drug|Organic Chemical|General Exam|7467,7476|false|false|false|C0073374|rifaximin|rifaximin
Drug|Pharmacologic Substance|General Exam|7467,7476|false|false|false|C0073374|rifaximin|rifaximin
Event|Event|General Exam|7467,7476|false|false|false|||rifaximin
Disorder|Disease or Syndrome|General Exam|7484,7487|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Disorder|Virus|General Exam|7484,7487|false|false|false|C0019196;C0220847|Hepatitis C;hepatitis C virus|HCV
Event|Event|General Exam|7484,7487|false|false|false|||HCV
Disorder|Disease or Syndrome|General Exam|7488,7497|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|General Exam|7488,7497|false|false|false|||Cirrhosis
Procedure|Laboratory Procedure|General Exam|7499,7507|false|false|false|C1285573|Genotype determination|Genotype
Event|Event|General Exam|7508,7510|false|false|false|||3a
Finding|Body Substance|General Exam|7512,7519|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|7512,7519|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|7512,7519|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Event|Event|General Exam|7523,7536|false|false|false|||decompensated
Disorder|Disease or Syndrome|General Exam|7554,7561|false|false|false|C0003962|Ascites|ascites
Event|Event|General Exam|7554,7561|false|false|false|||ascites
Finding|Pathologic Function|General Exam|7554,7561|false|false|false|C5441966|Peritoneal Effusion|ascites
Event|Event|General Exam|7566,7575|false|false|false|||worsening
Anatomy|Body Location or Region|General Exam|7576,7583|false|false|false|C0205054|Hepatic|hepatic
Disorder|Disease or Syndrome|General Exam|7576,7598|false|false|false|C0019151|Hepatic Encephalopathy|hepatic encephalopathy
Disorder|Disease or Syndrome|General Exam|7584,7598|false|false|false|C0085584|Encephalopathies|encephalopathy
Event|Event|General Exam|7584,7598|false|false|false|||encephalopathy
Event|Event|General Exam|7608,7617|false|false|false|||dependent
Finding|Functional Concept|General Exam|7608,7617|false|false|false|C3244310|dependent|dependent
Event|Event|General Exam|7634,7646|false|false|false|||paracentesis
Procedure|Therapeutic or Preventive Procedure|General Exam|7634,7646|false|false|false|C0034115|Paracentesis|paracentesis
Drug|Organic Chemical|General Exam|7648,7662|false|false|false|C0037982|spironolactone|Spironolactone
Drug|Pharmacologic Substance|General Exam|7648,7662|false|false|false|C0037982|spironolactone|Spironolactone
Event|Event|General Exam|7648,7662|false|false|false|||Spironolactone
Event|Event|General Exam|7677,7684|false|false|false|||stopped
Event|Event|General Exam|7692,7704|false|false|false|||hyperkalemia
Finding|Finding|General Exam|7692,7704|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Finding|Body Substance|General Exam|7706,7713|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|7706,7713|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|7706,7713|true|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Anatomy|Tissue|General Exam|7724,7734|true|false|false|C0332835|Transplanted tissue|transplant
Finding|Finding|General Exam|7724,7734|true|false|false|C0478647;C3841811|Transplant;Transplanted organ and tissue status|transplant
Procedure|Therapeutic or Preventive Procedure|General Exam|7724,7734|true|false|false|C0040732|Transplantation|transplant
Event|Event|General Exam|7735,7744|true|false|false|||candidate
Finding|Conceptual Entity|General Exam|7735,7744|true|false|false|C4527371|Candidate|candidate
Finding|Finding|General Exam|7755,7768|true|false|false|C0009488|Comorbidity|comorbidities
Disorder|Disease or Syndrome|General Exam|7769,7773|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|7769,7773|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|7769,7773|false|false|false|||COPD
Finding|Gene or Genome|General Exam|7769,7773|false|false|false|C1412502|ARCN1 gene|COPD
Event|Event|General Exam|7778,7788|false|false|false|||outpatient
Finding|Classification|General Exam|7778,7788|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|7778,7788|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Event|Event|General Exam|7790,7802|false|false|false|||hepatologist
Finding|Body Substance|General Exam|7808,7815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Idea or Concept|General Exam|7808,7815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Finding|Intellectual Product|General Exam|7808,7815|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|patient
Event|Event|General Exam|7822,7826|false|false|false|||like
Event|Event|General Exam|7830,7838|false|false|false|||continue
Event|Event|General Exam|7849,7861|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|7849,7861|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|General Exam|7868,7878|false|false|false|||outpatient
Finding|Classification|General Exam|7868,7878|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|7868,7878|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Disorder|Disease or Syndrome|General Exam|7883,7886|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|7883,7886|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|7883,7886|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|7883,7886|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|7883,7886|false|false|false|||HIV
Drug|Amino Acid, Peptide, or Protein|General Exam|7900,7903|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Biologically Active Substance|General Exam|7900,7903|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Drug|Immunologic Factor|General Exam|7900,7903|false|false|false|C0003323;C4048280|CD4 Antigens;T-Cell Surface Glycoprotein CD4, human|CD4
Finding|Gene or Genome|General Exam|7900,7903|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Finding|Receptor|General Exam|7900,7903|false|false|false|C0003323;C1332714|CD4 Antigens;CD4 gene|CD4
Procedure|Laboratory Procedure|General Exam|7900,7909|false|false|false|C0243009;C3541261|CD4 Count determination procedure;CD4 Expressing Cell Count|CD4 count
Event|Event|General Exam|7904,7909|false|false|false|||count
Disorder|Disease or Syndrome|General Exam|7922,7925|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|7922,7925|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|7922,7925|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|7922,7925|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|7922,7925|false|false|false|||HIV
Procedure|Laboratory Procedure|General Exam|7922,7936|false|false|false|C1168369|HIV viral load|HIV viral load
Finding|Functional Concept|General Exam|7926,7931|false|false|false|C0521026|Viral|viral
Finding|Finding|General Exam|7926,7936|false|false|false|C0376705|Viral Load result|viral load
Procedure|Laboratory Procedure|General Exam|7926,7936|false|false|false|C1261478|Viral load (procedure)|viral load
Event|Activity|General Exam|7932,7936|false|false|false|C1708715|Loading Technique|load
Event|Event|General Exam|7932,7936|false|false|false|||load
Finding|Idea or Concept|General Exam|7932,7936|false|false|false|C1550025|Load - Remote control command|load
Attribute|Clinical Attribute|General Exam|7949,7961|false|false|false|C3827727|Undetectable|undetectable
Event|Event|General Exam|7949,7961|false|false|false|||undetectable
Event|Event|General Exam|7971,7980|false|false|false|||continued
Finding|Idea or Concept|General Exam|7988,7992|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|7988,7992|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|7988,7992|false|false|false|C1553498|home health encounter|home
Event|Event|General Exam|7993,8000|false|false|false|||regimen
Finding|Intellectual Product|General Exam|7993,8000|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|General Exam|7993,8000|false|false|false|C0040808|Treatment Protocols|regimen
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8005,8016|false|false|false|C1871526|raltegravir|raltegravir
Drug|Pharmacologic Substance|General Exam|8005,8016|false|false|false|C1871526|raltegravir|raltegravir
Event|Event|General Exam|8005,8016|false|false|false|||raltegravir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8018,8031|false|false|false|C0909839|emtricitabine|emtricitabine
Drug|Pharmacologic Substance|General Exam|8018,8031|false|false|false|C0909839|emtricitabine|emtricitabine
Event|Event|General Exam|8018,8031|false|false|false|||emtricitabine
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8037,8046|false|false|false|C0384228|tenofovir|tenofovir
Drug|Pharmacologic Substance|General Exam|8037,8046|false|false|false|C0384228|tenofovir|tenofovir
Event|Event|General Exam|8037,8046|false|false|false|||tenofovir
Drug|Organic Chemical|General Exam|8048,8055|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|General Exam|8048,8055|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|General Exam|8057,8068|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|General Exam|8057,8068|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Event|Event|General Exam|8073,8077|false|false|false|||held
Event|Event|General Exam|8085,8094|false|false|false|||admission
Procedure|Health Care Activity|General Exam|8085,8094|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|admission
Event|Event|General Exam|8106,8118|false|false|false|||hyperkalemia
Finding|Finding|General Exam|8106,8118|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|hyperkalemia
Disorder|Disease or Syndrome|General Exam|8127,8131|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|8127,8131|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|8127,8131|false|false|false|||COPD
Finding|Gene or Genome|General Exam|8127,8131|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Body Substance|General Exam|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Idea or Concept|General Exam|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Intellectual Product|General Exam|8133,8140|false|false|false|C1550655;C1578481;C1578483;C1578484;C1578485;C1578486|Disabled Person Code - Patient;Mail Claim Party - Patient;Relationship modifier - Patient;Report source - Patient;Specimen Type - Patient|Patient
Finding|Finding|General Exam|8150,8157|false|false|false|C4534363|At home|at home
Event|Event|General Exam|8153,8157|false|false|false|||home
Finding|Idea or Concept|General Exam|8153,8157|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|8153,8157|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|8153,8157|false|false|false|C1553498|home health encounter|home
Event|Event|General Exam|8167,8176|false|false|false|||continued
Event|Event|General Exam|8184,8188|false|false|false|||home
Finding|Idea or Concept|General Exam|8184,8188|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Finding|Intellectual Product|General Exam|8184,8188|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|home
Procedure|Health Care Activity|General Exam|8184,8188|false|false|false|C1553498|home health encounter|home
Event|Event|General Exam|8190,8197|false|false|false|||regimen
Finding|Intellectual Product|General Exam|8190,8197|false|false|false|C5237222|GDC Regimen Terminology|regimen
Procedure|Therapeutic or Preventive Procedure|General Exam|8190,8197|false|false|false|C0040808|Treatment Protocols|regimen
Finding|Idea or Concept|General Exam|8200,8212|false|false|false|C1548597|Marketing basis - Transitional|TRANSITIONAL
Event|Event|General Exam|8213,8219|false|false|false|||ISSUES
Finding|Functional Concept|General Exam|8222,8228|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|General Exam|8222,8228|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|General Exam|8222,8231|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|General Exam|8222,8231|false|false|false|C1522577|follow-up|Follow up
Event|Event|General Exam|8229,8231|false|false|false|||up
Finding|Finding|General Exam|8237,8252|false|false|false|C0700049|Encounter due to palliative care|Palliative Care
Procedure|Health Care Activity|General Exam|8237,8252|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Procedure|Therapeutic or Preventive Procedure|General Exam|8237,8252|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Event|Activity|General Exam|8248,8252|false|false|false|C1947933|care activity|Care
Event|Event|General Exam|8248,8252|false|false|false|||Care
Finding|Finding|General Exam|8248,8252|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|General Exam|8248,8252|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|General Exam|8256,8266|false|false|false|||outpatient
Finding|Classification|General Exam|8256,8266|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|8256,8266|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|General Exam|8268,8275|false|false|false|C0591139|Bactrim|Bactrim
Drug|Pharmacologic Substance|General Exam|8268,8275|false|false|false|C0591139|Bactrim|Bactrim
Event|Event|General Exam|8276,8287|false|false|false|||prophylaxis
Procedure|Therapeutic or Preventive Procedure|General Exam|8276,8287|false|false|false|C0199176|Prophylactic treatment|prophylaxis
Disorder|Disease or Syndrome|General Exam|8289,8292|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|8289,8292|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|8289,8292|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|8289,8292|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|8289,8292|false|false|false|||HIV
Lab|Laboratory or Test Result|General Exam|8289,8293|false|false|false|C0019699|HIV Seropositivity|HIV+
Event|Event|General Exam|8299,8303|false|false|false|||held
Finding|Idea or Concept|General Exam|8311,8319|false|false|false|C1547192|Organization unit type - Hospital|hospital
Attribute|Clinical Attribute|General Exam|8311,8326|false|false|false|C0488549||hospital course
Finding|Finding|General Exam|8311,8326|false|false|false|C0489547|Hospital course|hospital course
Event|Event|General Exam|8320,8326|false|false|false|||course
Event|Event|General Exam|8340,8348|false|false|false|||Consider
Event|Event|General Exam|8349,8359|false|false|false|||restarting
Event|Event|General Exam|8363,8373|false|false|false|||outpatient
Finding|Classification|General Exam|8363,8373|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|8363,8373|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Drug|Organic Chemical|General Exam|8376,8386|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|General Exam|8376,8386|false|false|false|C0016860|furosemide|Furosemide
Event|Event|General Exam|8376,8386|false|false|false|||Furosemide
Event|Event|General Exam|8391,8395|false|false|false|||held
Event|Event|General Exam|8408,8416|false|false|false|||consider
Event|Event|General Exam|8417,8427|false|false|false|||restarting
Event|Event|General Exam|8432,8442|false|false|false|||outpatient
Finding|Classification|General Exam|8432,8442|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Idea or Concept|General Exam|8432,8442|false|false|false|C1548439;C1549405|Patient Class - Outpatient;Referral category - Outpatient|outpatient
Finding|Functional Concept|General Exam|8444,8450|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Intellectual Product|General Exam|8444,8450|false|false|false|C1719822;C4281991|Follow;Follow - dosing instruction imperative|Follow
Finding|Finding|General Exam|8444,8453|false|false|false|C0589120|Follow-up status|Follow up
Procedure|Health Care Activity|General Exam|8444,8453|false|false|false|C1522577|follow-up|Follow up
Event|Event|General Exam|8451,8453|false|false|false|||up
Event|Event|General Exam|8459,8469|false|false|false|||hepatology
Event|Event|General Exam|8471,8479|false|false|false|||Continue
Finding|Idea or Concept|General Exam|8471,8479|false|false|false|C0549178|Continuous|Continue
Event|Event|General Exam|8502,8514|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|General Exam|8502,8514|false|false|false|C0034115|Paracentesis|paracenteses
Event|Occupational Activity|General Exam|8516,8520|false|false|false|C0009219|Coding|Code
Finding|Intellectual Product|General Exam|8516,8520|false|false|false|C0805701;C0919279;C1554100|A Codes;Code;MDF Attribute Type - Code|Code
Procedure|Health Care Activity|General Exam|8516,8527|false|false|false|C0742531|CODE STATUS|Code status
Attribute|Clinical Attribute|General Exam|8521,8527|false|false|false|C5889824||status
Event|Event|General Exam|8521,8527|false|false|false|||status
Finding|Idea or Concept|General Exam|8521,8527|false|false|false|C1546481|What subject filter - Status|status
Attribute|Clinical Attribute|General Exam|8529,8532|false|false|false|C4285234||DNR
Drug|Antibiotic|General Exam|8529,8532|false|false|false|C0011015|daunorubicin|DNR
Drug|Organic Chemical|General Exam|8529,8532|false|false|false|C0011015|daunorubicin|DNR
Event|Event|General Exam|8529,8532|false|false|false|||DNR
Finding|Finding|General Exam|8529,8532|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Finding|Intellectual Product|General Exam|8529,8532|false|false|false|C0079252;C0582114|Do not resuscitate status;Do-Not-Resuscitate Orders|DNR
Attribute|Clinical Attribute|General Exam|8539,8550|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|General Exam|8539,8550|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|General Exam|8539,8550|false|false|false|||Medications
Finding|Intellectual Product|General Exam|8539,8550|false|false|false|C4284232|Medications|Medications
Finding|Finding|General Exam|8539,8563|false|false|false|C1627937|Medications on admission|Medications on Admission
Event|Event|General Exam|8554,8563|false|false|false|||Admission
Procedure|Health Care Activity|General Exam|8554,8563|false|false|false|C0184666;C0809949|Admission activity;Hospital admission|Admission
Drug|Pharmacologic Substance|General Exam|8582,8592|false|false|false|C0013227|Pharmaceutical Preparations|Medication
Finding|Intellectual Product|General Exam|8582,8592|false|false|false|C3244316;C4284232|Medications;medication - HL7 publishing domain|Medication
Finding|Intellectual Product|General Exam|8582,8597|false|false|false|C0746470|MEDICATION LIST|Medication list
Event|Event|General Exam|8593,8597|false|false|false|||list
Finding|Intellectual Product|General Exam|8593,8597|false|false|false|C0745732;C3272378|List;Sequence Data Type|list
Event|Event|General Exam|8601,8609|false|false|false|||accurate
Drug|Organic Chemical|General Exam|8614,8622|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Pharmacologic Substance|General Exam|8614,8622|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Drug|Vitamin|General Exam|8614,8622|false|false|false|C1815293|Complete, Multiple Vitamins with Iron|complete
Event|Event|General Exam|8614,8622|false|false|false|||complete
Finding|Functional Concept|General Exam|8614,8622|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Finding|Idea or Concept|General Exam|8614,8622|false|false|false|C1548561;C1706059;C3853530|Completion Status for valid values - Complete;Data operation - complete;Finish - dosing instruction imperative|complete
Drug|Organic Chemical|General Exam|8627,8636|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|General Exam|8627,8636|false|false|false|C0022957|lactulose|Lactulose
Event|Event|General Exam|8646,8649|false|false|false|||TID
Drug|Organic Chemical|General Exam|8654,8664|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|General Exam|8654,8664|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|General Exam|8654,8664|false|false|false|||Tiotropium
Drug|Organic Chemical|General Exam|8654,8672|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|General Exam|8654,8672|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|General Exam|8665,8672|false|false|false|C0006222|Bromides|Bromide
Event|Event|General Exam|8665,8672|false|false|false|||Bromide
Procedure|Laboratory Procedure|General Exam|8665,8672|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|General Exam|8675,8678|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|General Exam|8675,8678|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|General Exam|8675,8678|false|false|false|||CAP
Finding|Gene or Genome|General Exam|8675,8678|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|General Exam|8675,8678|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8692,8703|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|General Exam|8692,8703|false|false|false|C1871526|raltegravir|Raltegravir
Disorder|Mental or Behavioral Dysfunction|General Exam|8714,8717|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8714,8717|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8714,8717|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8714,8717|false|false|false|||BID
Finding|Gene or Genome|General Exam|8714,8717|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8722,8735|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|General Exam|8722,8735|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|General Exam|8722,8745|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|General Exam|8722,8745|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8736,8745|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|General Exam|8736,8745|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|8747,8754|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|General Exam|8747,8754|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|General Exam|8758,8761|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|General Exam|8758,8761|false|false|false|||TAB
Drug|Organic Chemical|General Exam|8775,8785|false|false|false|C0016860|furosemide|Furosemide
Drug|Pharmacologic Substance|General Exam|8775,8785|false|false|false|C0016860|furosemide|Furosemide
Drug|Organic Chemical|General Exam|8805,8813|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|General Exam|8805,8813|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|General Exam|8805,8813|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|General Exam|8805,8813|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|General Exam|8815,8821|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|General Exam|8815,8821|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|General Exam|8836,8839|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|8840,8844|false|false|false|C2598155||Pain
Event|Event|General Exam|8840,8844|false|false|false|||Pain
Finding|Functional Concept|General Exam|8840,8844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Finding|Sign or Symptom|General Exam|8840,8844|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|Pain
Drug|Organic Chemical|General Exam|8849,8860|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|General Exam|8849,8860|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|General Exam|8849,8860|false|false|false|||Fluticasone
Drug|Organic Chemical|General Exam|8849,8871|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|General Exam|8849,8871|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|General Exam|8861,8871|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|General Exam|8872,8878|false|false|false|||110mcg
Event|Event|General Exam|8881,8885|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|General Exam|8889,8892|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8889,8892|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8889,8892|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8889,8892|false|false|false|||BID
Finding|Gene or Genome|General Exam|8889,8892|false|false|false|C1332410|BID gene|BID
Drug|Biologically Active Substance|General Exam|8897,8904|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|8897,8904|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|8897,8904|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|8897,8904|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|8897,8904|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|8897,8904|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|8897,8904|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|8897,8904|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|General Exam|8897,8914|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|General Exam|8897,8914|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|General Exam|8905,8914|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|General Exam|8905,8914|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|General Exam|8905,8914|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Event|Event|General Exam|8905,8914|false|false|false|||Carbonate
Disorder|Mental or Behavioral Dysfunction|General Exam|8925,8928|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8925,8928|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8925,8928|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8925,8928|false|false|false|||BID
Finding|Gene or Genome|General Exam|8925,8928|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8933,8942|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|General Exam|8933,8942|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|General Exam|8953,8956|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|8953,8956|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|8953,8956|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|8953,8956|false|false|false|||BID
Finding|Gene or Genome|General Exam|8953,8956|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|8962,8971|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|General Exam|8962,8971|false|false|false|C0001927|albuterol|albuterol
Event|Event|General Exam|8962,8971|false|false|false|||albuterol
Drug|Organic Chemical|General Exam|8962,8979|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|General Exam|8962,8979|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|General Exam|8972,8979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|General Exam|8972,8979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|General Exam|8972,8979|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|General Exam|8972,8979|false|false|false|||sulfate
Finding|Functional Concept|General Exam|8997,9007|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|General Exam|8997,9007|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|General Exam|9008,9011|false|false|false|||Q6H
Finding|Gene or Genome|General Exam|9012,9015|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|General Exam|9017,9025|false|false|false|C0043144|Wheezing|Wheezing
Drug|Antibiotic|General Exam|9041,9053|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Organic Chemical|General Exam|9041,9053|false|false|false|C0041041|trimethoprim|Trimethoprim
Drug|Biomedical or Dental Material|General Exam|9059,9062|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|General Exam|9059,9062|false|false|false|||TAB
Event|Event|General Exam|9076,9085|false|false|false|||Discharge
Finding|Body Substance|General Exam|9076,9085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|9076,9085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|9076,9085|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|9076,9085|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|9076,9097|false|false|false|C0806915|Medication.discharge|Discharge Medications
Attribute|Clinical Attribute|General Exam|9086,9097|false|false|false|C0802604;C2598133||Medications
Drug|Pharmacologic Substance|General Exam|9086,9097|false|false|false|C0013227|Pharmaceutical Preparations|Medications
Event|Event|General Exam|9086,9097|false|false|false|||Medications
Finding|Intellectual Product|General Exam|9086,9097|false|false|false|C4284232|Medications|Medications
Drug|Biologically Active Substance|General Exam|9102,9109|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Element, Ion, or Isotope|General Exam|9102,9109|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Inorganic Chemical|General Exam|9102,9109|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Pharmacologic Substance|General Exam|9102,9109|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Drug|Vitamin|General Exam|9102,9109|false|false|false|C0006675;C0006726;C2936886;C3540037;C3714611|CALCIUM SUPPLEMENTS;Calcium Drug Class;Calcium [EPC];Calcium, Dietary;calcium|Calcium
Event|Event|General Exam|9102,9109|false|false|false|||Calcium
Finding|Physiologic Function|General Exam|9102,9109|false|false|false|C4553026|Calcium metabolic function|Calcium
Procedure|Laboratory Procedure|General Exam|9102,9109|false|false|false|C0201925|Calcium measurement|Calcium
Drug|Inorganic Chemical|General Exam|9102,9119|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Pharmacologic Substance|General Exam|9102,9119|false|false|false|C0006681|calcium carbonate|Calcium Carbonate
Drug|Element, Ion, or Isotope|General Exam|9110,9119|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Organic Chemical|General Exam|9110,9119|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Drug|Pharmacologic Substance|General Exam|9110,9119|false|false|false|C0007026;C3715099|Carbonates;carbonate ion|Carbonate
Disorder|Mental or Behavioral Dysfunction|General Exam|9130,9133|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9130,9133|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9130,9133|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9130,9133|false|false|false|||BID
Finding|Gene or Genome|General Exam|9130,9133|false|false|false|C1332410|BID gene|BID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|9138,9151|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Pharmacologic Substance|General Exam|9138,9151|false|false|false|C0909839|emtricitabine|Emtricitabine
Drug|Organic Chemical|General Exam|9138,9161|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Pharmacologic Substance|General Exam|9138,9161|false|false|false|C1532298|Emtricitabine- and tenofovir-containing product|Emtricitabine-Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|9152,9161|false|false|false|C0384228|tenofovir|Tenofovir
Drug|Pharmacologic Substance|General Exam|9152,9161|false|false|false|C0384228|tenofovir|Tenofovir
Event|Event|General Exam|9152,9161|false|false|false|||Tenofovir
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|9163,9170|false|false|false|C1528494|Truvada|Truvada
Drug|Pharmacologic Substance|General Exam|9163,9170|false|false|false|C1528494|Truvada|Truvada
Drug|Biomedical or Dental Material|General Exam|9174,9177|false|false|false|C0039225|Tablet Dosage Form|TAB
Event|Event|General Exam|9174,9177|false|false|false|||TAB
Drug|Organic Chemical|General Exam|9191,9202|false|false|false|C0082607|fluticasone|Fluticasone
Drug|Pharmacologic Substance|General Exam|9191,9202|false|false|false|C0082607|fluticasone|Fluticasone
Event|Event|General Exam|9191,9202|false|false|false|||Fluticasone
Drug|Organic Chemical|General Exam|9191,9213|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Pharmacologic Substance|General Exam|9191,9213|false|false|false|C0117996|fluticasone propionate|Fluticasone Propionate
Drug|Organic Chemical|General Exam|9203,9213|false|false|false|C0033474;C0392214|Propionates;propionate|Propionate
Event|Event|General Exam|9223,9227|false|false|false|||PUFF
Disorder|Mental or Behavioral Dysfunction|General Exam|9231,9234|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9231,9234|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9231,9234|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9231,9234|false|false|false|||BID
Finding|Gene or Genome|General Exam|9231,9234|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|9239,9248|false|false|false|C0022957|lactulose|Lactulose
Drug|Pharmacologic Substance|General Exam|9239,9248|false|false|false|C0022957|lactulose|Lactulose
Event|Event|General Exam|9239,9248|false|false|false|||Lactulose
Event|Event|General Exam|9258,9261|false|false|false|||TID
Drug|Nucleic Acid, Nucleoside, or Nucleotide|General Exam|9266,9277|false|false|false|C1871526|raltegravir|Raltegravir
Drug|Pharmacologic Substance|General Exam|9266,9277|false|false|false|C1871526|raltegravir|Raltegravir
Disorder|Mental or Behavioral Dysfunction|General Exam|9288,9291|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9288,9291|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9288,9291|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9288,9291|false|false|false|||BID
Finding|Gene or Genome|General Exam|9288,9291|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|9296,9305|false|false|false|C0073374|rifaximin|Rifaximin
Drug|Pharmacologic Substance|General Exam|9296,9305|false|false|false|C0073374|rifaximin|Rifaximin
Disorder|Mental or Behavioral Dysfunction|General Exam|9316,9319|false|false|false|C4546282|Body integrity dysphoria|BID
Drug|Amino Acid, Peptide, or Protein|General Exam|9316,9319|false|false|false|C1530795|BID protein, human|BID
Drug|Biologically Active Substance|General Exam|9316,9319|false|false|false|C1530795|BID protein, human|BID
Event|Event|General Exam|9316,9319|false|false|false|||BID
Finding|Gene or Genome|General Exam|9316,9319|false|false|false|C1332410|BID gene|BID
Drug|Organic Chemical|General Exam|9324,9332|false|false|false|C0040610|tramadol|TraMADOL
Drug|Pharmacologic Substance|General Exam|9324,9332|false|false|false|C0040610|tramadol|TraMADOL
Event|Event|General Exam|9324,9332|false|false|false|||TraMADOL
Procedure|Laboratory Procedure|General Exam|9324,9332|false|false|false|C1266765|Tramadol measurement (procedure)|TraMADOL
Drug|Organic Chemical|General Exam|9334,9340|false|false|false|C0724054|Ultram|Ultram
Drug|Pharmacologic Substance|General Exam|9334,9340|false|false|false|C0724054|Ultram|Ultram
Finding|Gene or Genome|General Exam|9356,9359|false|false|false|C1422467|CIAO3 gene|PRN
Attribute|Clinical Attribute|General Exam|9360,9364|false|false|false|C2598155||pain
Event|Event|General Exam|9360,9364|false|false|false|||pain
Finding|Functional Concept|General Exam|9360,9364|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Finding|Sign or Symptom|General Exam|9360,9364|false|false|false|C0030193;C1549543|Administration Method - Pain;Pain|pain
Drug|Organic Chemical|General Exam|9369,9378|false|false|false|C0001927|albuterol|albuterol
Drug|Pharmacologic Substance|General Exam|9369,9378|false|false|false|C0001927|albuterol|albuterol
Event|Event|General Exam|9369,9378|false|false|false|||albuterol
Drug|Organic Chemical|General Exam|9369,9386|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Pharmacologic Substance|General Exam|9369,9386|false|false|false|C0543495|albuterol sulfate|albuterol sulfate
Drug|Element, Ion, or Isotope|General Exam|9379,9386|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Inorganic Chemical|General Exam|9379,9386|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Drug|Pharmacologic Substance|General Exam|9379,9386|false|false|false|C0038720;C0475337;C3536965|Sulfates, Inorganic;Sulfates, Unspecified or Sulfate Ion;sulfate ion|sulfate
Event|Event|General Exam|9379,9386|false|false|false|||sulfate
Finding|Functional Concept|General Exam|9404,9414|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Finding|Organism Function|General Exam|9404,9414|false|false|false|C0004048;C0205535|Inhalation Route of Administration;Inspiration (function)|inhalation
Event|Event|General Exam|9415,9418|false|false|false|||Q6H
Finding|Gene or Genome|General Exam|9419,9422|false|false|false|C1422467|CIAO3 gene|PRN
Finding|Sign or Symptom|General Exam|9424,9432|false|false|false|C0043144|Wheezing|Wheezing
Drug|Organic Chemical|General Exam|9437,9447|false|false|false|C0213771|tiotropium|Tiotropium
Drug|Pharmacologic Substance|General Exam|9437,9447|false|false|false|C0213771|tiotropium|Tiotropium
Event|Event|General Exam|9437,9447|false|false|false|||Tiotropium
Drug|Organic Chemical|General Exam|9437,9455|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Pharmacologic Substance|General Exam|9437,9455|false|false|false|C1306772|tiotropium bromide|Tiotropium Bromide
Drug|Inorganic Chemical|General Exam|9448,9455|false|false|false|C0006222|Bromides|Bromide
Event|Event|General Exam|9448,9455|false|false|false|||Bromide
Procedure|Laboratory Procedure|General Exam|9448,9455|false|false|false|C0202341|Bromides measurement|Bromide
Disorder|Congenital Abnormality|General Exam|9458,9461|false|false|false|C1855179|CATARACT, ANTERIOR POLAR|CAP
Drug|Biomedical or Dental Material|General Exam|9458,9461|false|false|false|C0006935|capsule (pharmacologic)|CAP
Event|Event|General Exam|9458,9461|false|false|false|||CAP
Finding|Gene or Genome|General Exam|9458,9461|false|false|false|C1416891;C1418551;C1419093;C1422073;C1422760;C2985259;C4522312|BRD4 gene;BRD4 wt Allele;CAP1 gene;HACD1 gene;LNPEP gene;SERPINB6 gene;SORBS1 gene|CAP
Procedure|Therapeutic or Preventive Procedure|General Exam|9458,9461|false|false|false|C0278651;C0280547;C1879916|CAP Regimen;cisplatin/cyclophosphamide/doxorubicin protocol;cyclophosphamide/doxorubicin/prednisone protocol|CAP
Event|Event|General Exam|9475,9484|false|false|false|||Discharge
Finding|Body Substance|General Exam|9475,9484|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|9475,9484|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|9475,9484|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|9475,9484|false|false|false|C0030685|Patient Discharge|Discharge
Attribute|Clinical Attribute|General Exam|9475,9496|false|false|false|C4019243||Discharge Disposition
Finding|Finding|General Exam|9475,9496|false|false|false|C4759848|Discharge disposition|Discharge Disposition
Attribute|Clinical Attribute|General Exam|9485,9496|false|false|false|C2926604||Disposition
Event|Event|General Exam|9485,9496|false|false|false|||Disposition
Procedure|Health Care Activity|General Exam|9485,9496|false|false|false|C0184758|Patient disposition|Disposition
Event|Event|General Exam|9498,9502|false|false|false|||Home
Finding|Idea or Concept|General Exam|9498,9502|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Finding|Intellectual Product|General Exam|9498,9502|false|false|false|C1548341;C1549632|Address type - Home;Visit User Code - Home|Home
Procedure|Health Care Activity|General Exam|9498,9502|false|false|false|C1553498|home health encounter|Home
Event|Event|General Exam|9505,9514|false|false|false|||Discharge
Finding|Body Substance|General Exam|9505,9514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Intellectual Product|General Exam|9505,9514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Finding|Sign or Symptom|General Exam|9505,9514|false|false|false|C0012621;C0600083;C1546601;C2926602|Body Fluid Discharge;Body Substance Discharge;Discharge Body Fluid|Discharge
Procedure|Health Care Activity|General Exam|9505,9514|false|false|false|C0030685|Patient Discharge|Discharge
Finding|Finding|General Exam|9505,9524|false|false|false|C1555319|discharge diagnosis|Discharge Diagnosis
Attribute|Clinical Attribute|General Exam|9515,9524|false|false|false|C0945731||Diagnosis
Event|Event|General Exam|9515,9524|false|false|false|||Diagnosis
Finding|Classification|General Exam|9515,9524|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Finding|Functional Concept|General Exam|9515,9524|false|false|false|C1546899;C1704338|Diagnosis Classification - Diagnosis;diagnosis aspects|Diagnosis
Procedure|Diagnostic Procedure|General Exam|9515,9524|false|false|false|C0011900|Diagnosis|Diagnosis
Finding|Finding|General Exam|9535,9546|false|false|false|C0020649|Hypotension|Hypotension
Event|Event|General Exam|9547,9559|false|false|false|||Hyperkalemia
Finding|Finding|General Exam|9547,9559|false|false|false|C0020461;C5700154|Hyperkalemia;Serum potassium level above reference range|Hyperkalemia
Finding|Intellectual Product|General Exam|9560,9565|false|false|false|C1547229;C1547295|Acute - Triage Code;Admission Level of Care Code - Acute|Acute
Disorder|Disease or Syndrome|General Exam|9560,9579|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute Kidney Injury
Disorder|Injury or Poisoning|General Exam|9560,9579|false|false|false|C0022660;C2609414|Acute kidney injury;Kidney Failure, Acute|Acute Kidney Injury
Anatomy|Body Part, Organ, or Organ Component|General Exam|9566,9572|false|false|false|C0022646;C0227665|Both kidneys;Kidney|Kidney
Disorder|Neoplastic Process|General Exam|9566,9572|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|Kidney
Event|Event|General Exam|9566,9572|false|false|false|||Kidney
Finding|Sign or Symptom|General Exam|9566,9572|false|false|false|C0812426|Kidney problem|Kidney
Procedure|Diagnostic Procedure|General Exam|9566,9572|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Procedure|Therapeutic or Preventive Procedure|General Exam|9566,9572|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|Kidney
Disorder|Injury or Poisoning|General Exam|9566,9579|false|false|false|C0160420|Injury of kidney|Kidney Injury
Disorder|Injury or Poisoning|General Exam|9573,9579|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|Injury
Event|Event|General Exam|9573,9579|false|false|false|||Injury
Disorder|Neoplastic Process|General Exam|9581,9590|false|false|false|C0027627|Neoplasm Metastasis|Secondary
Event|Event|General Exam|9581,9590|false|false|false|||Secondary
Finding|Functional Concept|General Exam|9581,9590|false|false|false|C1522484|metastatic qualifier|Secondary
Disorder|Disease or Syndrome|General Exam|9592,9595|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Disorder|Virus|General Exam|9592,9595|false|false|false|C0019682;C0019693|HIV;HIV Infections|HIV
Drug|Immunologic Factor|General Exam|9592,9595|false|false|false|C0086413|HIV Vaccine|HIV
Drug|Pharmacologic Substance|General Exam|9592,9595|false|false|false|C0086413|HIV Vaccine|HIV
Event|Event|General Exam|9592,9595|false|false|false|||HIV
Disorder|Disease or Syndrome|General Exam|9596,9605|false|false|false|C0023890;C1623038|Cirrhosis;Liver Cirrhosis|Cirrhosis
Event|Event|General Exam|9596,9605|false|false|false|||Cirrhosis
Disorder|Disease or Syndrome|General Exam|9606,9610|false|false|false|C0024117;C3714496|Chronic Obstructive Airway Disease;Chronic obstructive pulmonary disease of horses|COPD
Drug|Pharmacologic Substance|General Exam|9606,9610|false|false|false|C1647218|COPD pharmacologic substance|COPD
Event|Event|General Exam|9606,9610|false|false|false|||COPD
Finding|Gene or Genome|General Exam|9606,9610|false|false|false|C1412502|ARCN1 gene|COPD
Finding|Mental Process|Discharge Condition|9634,9640|false|false|false|C0229992|Psyche structure|Mental
Attribute|Clinical Attribute|Discharge Condition|9634,9647|false|false|false|C0488568;C0488569||Mental Status
Finding|Finding|Discharge Condition|9634,9647|false|false|false|C0278060|Mental state|Mental Status
Attribute|Clinical Attribute|Discharge Condition|9641,9647|false|false|false|C5889824||Status
Finding|Idea or Concept|Discharge Condition|9641,9647|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9649,9654|false|false|false|||Clear
Finding|Idea or Concept|Discharge Condition|9649,9654|false|false|false|C1550016|Remote control command - Clear|Clear
Event|Event|Discharge Condition|9659,9667|false|false|false|||coherent
Finding|Finding|Discharge Condition|9659,9667|false|false|false|C4068804|Coherent|coherent
Event|Event|Discharge Condition|9669,9674|false|false|false|||Level
Attribute|Clinical Attribute|Discharge Condition|9669,9691|false|false|false|C4050479||Level of Consciousness
Finding|Finding|Discharge Condition|9669,9691|false|false|false|C0234425|Level of consciousness|Level of Consciousness
Event|Event|Discharge Condition|9678,9691|false|false|false|||Consciousness
Finding|Finding|Discharge Condition|9678,9691|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Finding|Mental Process|Discharge Condition|9678,9691|false|false|false|C0009791;C0234421;C0517960|Conscious;Consciousness related finding|Consciousness
Attribute|Clinical Attribute|Discharge Condition|9693,9698|false|false|false|C5890168||Alert
Drug|Organic Chemical|Discharge Condition|9693,9698|false|false|false|C0718338|Alert brand of caffeine|Alert
Drug|Pharmacologic Substance|Discharge Condition|9693,9698|false|false|false|C0718338|Alert brand of caffeine|Alert
Event|Event|Discharge Condition|9693,9698|false|false|false|||Alert
Finding|Finding|Discharge Condition|9693,9698|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Functional Concept|Discharge Condition|9693,9698|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Finding|Intellectual Product|Discharge Condition|9693,9698|false|false|false|C0239110;C0424536;C2004580;C3665546|Alert;Alert note;Consciousness clear;Mentally alert|Alert
Event|Event|Discharge Condition|9703,9714|false|false|false|||interactive
Finding|Functional Concept|Discharge Condition|9703,9714|false|false|false|C1704675|Interaction|interactive
Event|Activity|Discharge Condition|9716,9724|false|false|false|C0441655|Activities|Activity
Finding|Daily or Recreational Activity|Discharge Condition|9716,9724|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Finding|Finding|Discharge Condition|9716,9724|false|false|false|C0026606;C3668946|Activity (animal life circumstance);Physical activity|Activity
Attribute|Clinical Attribute|Discharge Condition|9725,9731|false|false|false|C5889824||Status
Event|Event|Discharge Condition|9725,9731|false|false|false|||Status
Finding|Idea or Concept|Discharge Condition|9725,9731|false|false|false|C1546481|What subject filter - Status|Status
Event|Event|Discharge Condition|9733,9743|false|false|false|||Ambulatory
Finding|Functional Concept|Discharge Condition|9733,9743|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Idea or Concept|Discharge Condition|9733,9743|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Finding|Intellectual Product|Discharge Condition|9733,9743|false|false|false|C0439841;C1547135;C1561561;C5401192|Ambulatory;Ambulatory (qualifier value);Level of Care - Ambulatory;Referral category - Ambulatory|Ambulatory
Procedure|Health Care Activity|Discharge Condition|9733,9743|false|false|false|C1561560|ambulatory encounter|Ambulatory
Event|Event|Discharge Condition|9746,9757|false|false|false|||Independent
Finding|Finding|Discharge Condition|9746,9757|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Idea or Concept|Discharge Condition|9746,9757|false|false|false|C0085862;C1299583;C1549571;C1608386|Coordination of Benefits - Independent;Independence;Independently able;Religious Affiliation - Independent|Independent
Finding|Gene or Genome|Discharge Instructions|9785,9789|false|false|false|C4320303|FBXW7-AS1 gene|Dear
Event|Event|Discharge Instructions|9809,9817|false|false|false|||admitted
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|9836,9845|false|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|9836,9845|false|false|false|||confusion
Finding|Finding|Discharge Instructions|9836,9845|false|false|false|C0683369|Clouded consciousness|confusion
Finding|Finding|Discharge Instructions|9847,9850|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Finding|Intellectual Product|Discharge Instructions|9847,9850|false|false|false|C1550472;C4522223;C5203106|IPSS Risk Category Low;IPSS-R Risk Category Low;low confidentiality|low
Disorder|Disease or Syndrome|Discharge Instructions|9851,9856|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|9851,9856|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|9851,9856|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Event|Event|Discharge Instructions|9858,9866|false|false|false|||pressure
Finding|Finding|Discharge Instructions|9858,9866|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|9858,9866|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|9858,9866|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|9858,9866|false|false|false|C0033095||pressure
Finding|Finding|Discharge Instructions|9874,9878|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Idea or Concept|Discharge Instructions|9874,9878|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Intellectual Product|Discharge Instructions|9874,9878|false|false|false|C1561958;C3887512;C4522209;C5200928;C5202936|High (finding);IPSS Risk Category High;IPSS-R Risk Category High;Message Waiting Priority - High;high - ActExposureLevelCode|high
Finding|Finding|Discharge Instructions|9874,9888|false|false|false|C0856882|Potassium increased|high potassium
Drug|Biologically Active Substance|Discharge Instructions|9879,9888|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Discharge Instructions|9879,9888|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Discharge Instructions|9879,9888|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Discharge Instructions|9879,9888|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Discharge Instructions|9879,9888|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Discharge Instructions|9879,9888|false|false|false|||potassium
Finding|Physiologic Function|Discharge Instructions|9879,9888|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Discharge Instructions|9879,9888|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Discharge Instructions|9889,9894|false|false|false|||value
Finding|Intellectual Product|Discharge Instructions|9889,9894|false|false|false|C1554112|MDF Attribute Type - Value|value
Disorder|Mental or Behavioral Dysfunction|Discharge Instructions|9901,9910|false|false|false|C0009676|Confusion|confusion
Event|Event|Discharge Instructions|9901,9910|false|false|false|||confusion
Finding|Finding|Discharge Instructions|9901,9910|false|false|false|C0683369|Clouded consciousness|confusion
Event|Event|Discharge Instructions|9911,9919|false|false|false|||improved
Drug|Organic Chemical|Discharge Instructions|9926,9935|false|false|false|C0022957|lactulose|lactulose
Drug|Pharmacologic Substance|Discharge Instructions|9926,9935|false|false|false|C0022957|lactulose|lactulose
Event|Event|Discharge Instructions|9926,9935|false|false|false|||lactulose
Disorder|Disease or Syndrome|Discharge Instructions|9942,9947|false|false|false|C0851353|Blood and lymphatic system disorders|blood
Event|Event|Discharge Instructions|9942,9947|false|false|false|||blood
Finding|Body Substance|Discharge Instructions|9942,9947|false|false|false|C0005767;C0005768;C0229664|Blood;In Blood;peripheral blood|blood
Finding|Finding|Discharge Instructions|9942,9956|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Finding|Organism Function|Discharge Instructions|9942,9956|false|false|false|C0005823;C1271104;C1272641|Blood Pressure;Blood pressure finding;Systemic arterial pressure|blood pressure
Procedure|Health Care Activity|Discharge Instructions|9942,9956|false|false|false|C0005824|Blood pressure determination|blood pressure
Event|Event|Discharge Instructions|9948,9956|false|false|false|||pressure
Finding|Finding|Discharge Instructions|9948,9956|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Functional Concept|Discharge Instructions|9948,9956|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Finding|Organ or Tissue Function|Discharge Instructions|9948,9956|false|false|false|C0234222;C0460139;C1306345|Baresthesia;Pressure (finding)|pressure
Phenomenon|Phenomenon or Process|Discharge Instructions|9948,9956|false|false|false|C0033095||pressure
Event|Event|Discharge Instructions|9957,9965|false|false|false|||improved
Drug|Substance|Discharge Instructions|9977,9983|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|9977,9983|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|9977,9983|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|9977,9983|false|false|false|C0016286|Fluid Therapy|fluids
Drug|Biologically Active Substance|Discharge Instructions|9994,10003|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Element, Ion, or Isotope|Discharge Instructions|9994,10003|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Food|Discharge Instructions|9994,10003|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Inorganic Chemical|Discharge Instructions|9994,10003|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Drug|Pharmacologic Substance|Discharge Instructions|9994,10003|false|false|false|C0032821;C0162800;C0304475;C3714637|Dietary Potassium;Potassium Drug Class;Potassium supplement;potassium|potassium
Event|Event|Discharge Instructions|9994,10003|false|false|false|||potassium
Finding|Physiologic Function|Discharge Instructions|9994,10003|false|false|false|C4553027|Potassium metabolic function|potassium
Procedure|Laboratory Procedure|Discharge Instructions|9994,10003|false|false|false|C0202194|Potassium measurement|potassium
Event|Event|Discharge Instructions|10004,10012|false|false|false|||improved
Finding|Finding|Discharge Instructions|10016,10020|false|false|false|C5575035|Well (answer to question)|well
Event|Event|Discharge Instructions|10041,10047|false|false|false|||degree
Finding|Intellectual Product|Discharge Instructions|10041,10047|false|false|false|C0542560|Academic degree|degree
Anatomy|Body Part, Organ, or Organ Component|Discharge Instructions|10052,10058|false|false|false|C0022646;C0227665|Both kidneys;Kidney|kidney
Disorder|Neoplastic Process|Discharge Instructions|10052,10058|false|false|false|C0496892;C0496927|Benign neoplasm of kidney;Neoplasm of uncertain or unknown behavior of kidney|kidney
Event|Event|Discharge Instructions|10052,10058|false|false|false|||kidney
Finding|Sign or Symptom|Discharge Instructions|10052,10058|false|false|false|C0812426|Kidney problem|kidney
Procedure|Diagnostic Procedure|Discharge Instructions|10052,10058|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10052,10058|false|false|false|C0869841;C4554465|Procedures on Kidney;examination of kidney|kidney
Disorder|Injury or Poisoning|Discharge Instructions|10052,10065|false|false|false|C0160420|Injury of kidney|kidney injury
Disorder|Injury or Poisoning|Discharge Instructions|10059,10065|false|false|false|C3263722;C3263723|Traumatic AND/OR non-traumatic injury;Traumatic injury|injury
Event|Event|Discharge Instructions|10059,10065|false|false|false|||injury
Event|Event|Discharge Instructions|10075,10079|false|false|false|||came
Finding|Idea or Concept|Discharge Instructions|10087,10095|false|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10112,10120|false|false|false|||improved
Drug|Substance|Discharge Instructions|10126,10132|false|false|false|C0302908|Liquid substance|fluids
Event|Event|Discharge Instructions|10126,10132|false|false|false|||fluids
Finding|Body Substance|Discharge Instructions|10126,10132|false|false|false|C1521806|Mouse Body Fluid or Substance|fluids
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10126,10132|false|false|false|C0016286|Fluid Therapy|fluids
Event|Event|Discharge Instructions|10159,10168|false|false|false|||discussed
Event|Event|Discharge Instructions|10170,10178|false|false|false|||changing
Attribute|Clinical Attribute|Discharge Instructions|10184,10189|false|false|false|C2979882||goals
Event|Event|Discharge Instructions|10184,10189|false|false|false|||goals
Finding|Idea or Concept|Discharge Instructions|10184,10189|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Finding|Intellectual Product|Discharge Instructions|10184,10189|false|false|false|C0018017;C0679840;C1546459|What subject filter - Goals;objective (goal);treatment goals|goals
Procedure|Health Care Activity|Discharge Instructions|10184,10197|false|false|false|C2930505|Goals of Care|goals of care
Event|Activity|Discharge Instructions|10193,10197|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|10193,10197|false|false|false|||care
Finding|Finding|Discharge Instructions|10193,10197|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10193,10197|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Event|Event|Discharge Instructions|10201,10209|false|false|false|||focusing
Attribute|Clinical Attribute|Discharge Instructions|10213,10220|false|false|false|C3854129||symptom
Finding|Sign or Symptom|Discharge Instructions|10213,10220|false|false|false|C1457887|Symptoms|symptom
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10213,10231|false|false|false|C0030231;C1536570|Palliative Care;Symptom Management|symptom management
Event|Event|Discharge Instructions|10221,10231|false|false|false|||management
Event|Occupational Activity|Discharge Instructions|10221,10231|false|false|false|C0001554;C1273870|Administration occupational activities;Management procedure|management
Procedure|Health Care Activity|Discharge Instructions|10221,10231|false|false|false|C0376636|Disease Management|management
Event|Event|Discharge Instructions|10237,10246|false|false|false|||treatment
Finding|Conceptual Entity|Discharge Instructions|10237,10246|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Finding|Functional Concept|Discharge Instructions|10237,10246|false|false|false|C0039798;C1522326;C1705169|Biomaterial Treatment;Treating;therapeutic aspects|treatment
Procedure|Health Care Activity|Discharge Instructions|10237,10246|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10237,10246|false|false|false|C0087111;C1533734;C3887704|Administration (procedure);Therapeutic procedure;treatment - ActInformationManagementReason|treatment
Finding|Functional Concept|Discharge Instructions|10250,10260|false|false|false|C0205343|Reversible|reversible
Event|Event|Discharge Instructions|10261,10270|false|false|false|||processes
Disorder|Disease or Syndrome|Discharge Instructions|10283,10292|false|false|false|C0009450|Communicable Diseases|infection
Event|Event|Discharge Instructions|10283,10292|false|false|false|||infection
Finding|Pathologic Function|Discharge Instructions|10283,10292|false|false|false|C3714514|Infection|infection
Finding|Idea or Concept|Discharge Instructions|10317,10325|true|false|false|C1547192|Organization unit type - Hospital|hospital
Event|Event|Discharge Instructions|10336,10340|false|false|false|||seen
Finding|Functional Concept|Discharge Instructions|10356,10362|false|false|false|C0728831|Social|social
Event|Event|Discharge Instructions|10363,10370|false|false|false|||workers
Event|Event|Discharge Instructions|10386,10392|false|false|false|||follow
Finding|Finding|Discharge Instructions|10401,10416|false|false|false|C0700049|Encounter due to palliative care|Palliative Care
Procedure|Health Care Activity|Discharge Instructions|10401,10416|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10401,10416|false|false|false|C0030231;C3816218|Palliative Care;Palliative Nursing|Palliative Care
Event|Activity|Discharge Instructions|10412,10416|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|10412,10416|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|10412,10416|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Event|Event|Discharge Instructions|10443,10451|false|false|false|||continue
Drug|Organic Chemical|Discharge Instructions|10460,10471|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Drug|Pharmacologic Substance|Discharge Instructions|10460,10471|false|false|false|C0723712|Therapeutic brand of coal tar|therapeutic
Event|Event|Discharge Instructions|10460,10471|false|false|false|||therapeutic
Finding|Functional Concept|Discharge Instructions|10460,10471|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Finding|Intellectual Product|Discharge Instructions|10460,10471|false|false|false|C0302350;C1547427|Therapeutic;Therapeutic - Location Service Code|therapeutic
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10460,10471|false|false|false|C0087111|Therapeutic procedure|therapeutic
Event|Event|Discharge Instructions|10472,10484|false|false|false|||paracenteses
Procedure|Therapeutic or Preventive Procedure|Discharge Instructions|10472,10484|false|false|false|C0034115|Paracentesis|paracenteses
Event|Event|Discharge Instructions|10501,10509|false|false|false|||pleasure
Finding|Intellectual Product|Discharge Instructions|10501,10509|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Finding|Mental Process|Discharge Instructions|10501,10509|false|false|false|C0679105;C1610547|Production Class Code - Pleasure;pleasurable emotion|pleasure
Event|Activity|Discharge Instructions|10517,10521|false|false|false|C1947933|care activity|care
Event|Event|Discharge Instructions|10517,10521|false|false|false|||care
Finding|Finding|Discharge Instructions|10517,10521|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10517,10521|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|care
Finding|Intellectual Product|Discharge Instructions|10517,10524|false|false|false|C1555558|care of - AddressPartType|care of
Disorder|Disease or Syndrome|Discharge Instructions|10554,10558|false|false|false|C0339510|Vitelliform Macular Dystrophy|best
Event|Event|Discharge Instructions|10554,10558|false|false|false|||best
Finding|Gene or Genome|Discharge Instructions|10554,10558|false|false|false|C1826421;C5781213|BEST1 gene;BEST1 wt Allele|best
Event|Activity|Discharge Instructions|10569,10573|false|false|false|C1947933|care activity|Care
Finding|Finding|Discharge Instructions|10569,10573|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Finding|Intellectual Product|Discharge Instructions|10569,10573|false|false|false|C0580931;C2362566|Continuity Assessment Record and Evaluation;In care (finding)|Care
Attribute|Clinical Attribute|Discharge Instructions|10569,10578|false|false|false|C4321316||Care team
Finding|Finding|Discharge Instructions|10569,10578|false|false|false|C4321315|Care team|Care team
Procedure|Health Care Activity|Discharge Instructions|10581,10589|false|false|false|C1522577|follow-up|Followup
Attribute|Clinical Attribute|Discharge Instructions|10590,10602|false|false|false|C3263700||Instructions
Event|Event|Discharge Instructions|10590,10602|false|false|false|||Instructions
Finding|Intellectual Product|Discharge Instructions|10590,10602|false|false|false|C0302828;C1442085|Instruction [Publication Type];Instructions|Instructions

