 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
MEDICINE|156,164
<EOL>|164,165
<EOL>|166,167
Allergies|167,176
:|176,177
<EOL>|178,179
lisinopril|179,189
<EOL>|189,190
<EOL>|191,192
Attending|192,201
:|201,202
_|203,204
_|204,205
_|205,206
<EOL>|206,207
<EOL>|208,209
Chief|209,214
Complaint|215,224
:|224,225
<EOL>|225,226
Chest|226,231
pain|232,236
<EOL>|236,237
<EOL>|238,239
Major|239,244
Surgical|245,253
or|254,256
Invasive|257,265
Procedure|266,275
:|275,276
<EOL>|276,277
Cardiac|277,284
cath|285,289
(|290,291
_|291,292
_|292,293
_|293,294
)|294,295
<EOL>|295,296
<EOL>|296,297
<EOL>|298,299
Past|299,303
Medical|304,311
History|312,319
:|319,320
<EOL>|320,321
-|321,322
COPD|322,326
<EOL>|326,327
-|327,328
CAD|328,331
s|332,333
/|333,334
p|334,335
BMS|336,339
proximal|340,348
-|348,349
LAD|349,352
_|353,354
_|354,355
_|355,356
,|356,357
DES|358,361
to|362,364
mid|365,368
LAD|369,372
_|373,374
_|374,375
_|375,376
,|376,377
DES|378,381
to|382,384
edge|385,389
<EOL>|390,391
ISR|391,394
of|395,397
mid|398,401
LAD|402,405
DES|406,409
and|410,413
stenosis|414,422
distal|423,429
to|430,432
stent|433,438
_|439,440
_|440,441
_|441,442
,|442,443
DES|444,447
to|448,450
OM1|451,454
<EOL>|455,456
_|456,457
_|457,458
_|458,459
,|459,460
s|461,462
/|462,463
p|463,464
3|465,466
v|467,468
CABG|469,473
LIMA|474,478
-|478,479
LAD|479,482
,|482,483
SVG|484,487
-|487,488
OM1|488,491
,|491,492
<EOL>|493,494
_|494,495
_|495,496
_|496,497
<EOL>|498,499
-|499,500
HFpEF|500,505
<EOL>|505,506
-|506,507
Depression|507,517
<EOL>|519,520
-|520,521
DM|521,523
<EOL>|525,526
-|526,527
GERD|527,531
<EOL>|533,534
-|534,535
Hypertension|535,547
<EOL>|547,548
-|548,549
Migraines|549,558
<EOL>|558,559
-|559,560
Chronic|560,567
shoulder|568,576
pain|577,581
on|582,584
narcotics|585,594
<EOL>|594,595
-|595,596
OSA|596,599
<EOL>|599,600
-|600,601
Peripheral|601,611
neuropathy|612,622
<EOL>|622,623
-|623,624
Restless|624,632
leg|633,636
<EOL>|636,637
<EOL>|638,639
Social|639,645
History|646,653
:|653,654
<EOL>|654,655
_|655,656
_|656,657
_|657,658
<EOL>|658,659
Family|659,665
History|666,673
:|673,674
<EOL>|674,675
Patient|675,682
was|683,686
ward|687,691
of|692,694
the|695,698
state|699,704
,|704,705
does|706,710
n't|710,713
know|714,718
full|719,723
details|724,731
of|732,734
<EOL>|735,736
family|736,742
history|743,750
.|750,751
Mother|752,758
with|759,763
possible|764,772
alcohol|773,780
abuse|781,786
.|786,787
Father|788,794
<EOL>|795,796
deceased|796,804
at|805,807
_|808,809
_|809,810
_|810,811
from|812,816
Hodgkin|817,824
's|824,826
Disease|827,834
per|835,838
old|839,842
records|843,850
.|850,851
<EOL>|851,852
<EOL>|853,854
Physical|854,862
Exam|863,867
:|867,868
<EOL>|868,869
ADMISSION|869,878
EXAM|879,883
<EOL>|883,884
=|884,885
=|885,886
=|886,887
=|887,888
=|888,889
=|889,890
=|890,891
=|891,892
=|892,893
=|893,894
=|894,895
=|895,896
=|896,897
=|897,898
<EOL>|898,899
GENERAL|899,906
:|906,907
NAD|907,910
AOx3|911,915
Pleasant|916,924
woman|925,930
.|930,931
<EOL>|932,933
HEENT|933,938
:|938,939
NCAT|940,944
.|944,945
Sclera|946,952
anicteric|953,962
.|962,963
PERRL|964,969
,|969,970
EOMI|971,975
.|975,976
Conjunctiva|977,988
pink|989,993
,|993,994
no|995,997
<EOL>|998,999
pallor|999,1005
or|1006,1008
cyanosis|1009,1017
of|1018,1020
the|1021,1024
oral|1025,1029
mucosa|1030,1036
<EOL>|1036,1037
NECK|1037,1041
:|1041,1042
Supple|1043,1049
with|1050,1054
no|1055,1057
JVD|1058,1061
<EOL>|1061,1062
CARDIAC|1062,1069
:|1069,1070
RRR|1071,1074
normal|1075,1081
S1|1082,1084
/|1084,1085
S2|1085,1087
.|1087,1088
No|1089,1091
thrills|1092,1099
,|1099,1100
lifts|1101,1106
.|1106,1107
<EOL>|1109,1110
LUNGS|1110,1115
:|1115,1116
CTAB|1117,1121
.|1121,1122
No|1123,1125
crackles|1126,1134
,|1134,1135
wheezes|1136,1143
or|1144,1146
rhonchi|1147,1154
.|1154,1155
<EOL>|1157,1158
ABDOMEN|1158,1165
:|1165,1166
Soft|1167,1171
,|1171,1172
NTND|1173,1177
.|1177,1178
No|1179,1181
HSM|1182,1185
or|1186,1188
tenderness|1189,1199
.|1199,1200
<EOL>|1202,1203
EXTREMITIES|1203,1214
:|1214,1215
No|1216,1218
_|1219,1220
_|1220,1221
_|1221,1222
edema|1223,1228
<EOL>|1228,1229
PULSES|1229,1235
:|1235,1236
_|1237,1238
_|1238,1239
_|1239,1240
and|1241,1244
DP|1245,1247
palpable|1248,1256
on|1257,1259
the|1260,1263
right|1264,1269
side|1270,1274
.|1274,1275
Did|1276,1279
not|1280,1283
take|1284,1288
<EOL>|1289,1290
bandage|1290,1297
down|1298,1302
for|1303,1306
exam|1307,1311
as|1312,1314
podiatry|1315,1323
had|1324,1327
just|1328,1332
dressed|1333,1340
.|1340,1341
<EOL>|1342,1343
<EOL>|1344,1345
<EOL>|1345,1346
DISCHARGE|1346,1355
EXAM|1356,1360
<EOL>|1360,1361
=|1361,1362
=|1362,1363
=|1363,1364
=|1364,1365
=|1365,1366
=|1366,1367
=|1367,1368
=|1368,1369
=|1369,1370
=|1370,1371
=|1371,1372
=|1372,1373
=|1373,1374
=|1374,1375
<EOL>|1375,1376
VITALS|1376,1382
:|1382,1383
_|1385,1386
_|1386,1387
_|1387,1388
0412|1389,1393
Temp|1394,1398
:|1398,1399
97.8|1400,1404
PO|1405,1407
BP|1408,1410
:|1410,1411
105|1412,1415
/|1415,1416
67|1416,1418
R|1419,1420
Lying|1421,1426
HR|1427,1429
:|1429,1430
71|1431,1433
<EOL>|1433,1434
RR|1434,1436
:|1436,1437
18|1438,1440
O2|1441,1443
sat|1444,1447
:|1447,1448
97|1449,1451
%|1451,1452
O2|1453,1455
delivery|1456,1464
:|1464,1465
Ra|1466,1468
<EOL>|1469,1470
GENERAL|1470,1477
:|1477,1478
NAD|1478,1481
AOx3|1482,1486
Pleasant|1487,1495
woman|1496,1501
.|1501,1502
<EOL>|1503,1504
HEENT|1504,1509
:|1509,1510
NCAT|1511,1515
.|1515,1516
Sclera|1517,1523
anicteric|1524,1533
.|1533,1534
PERRL|1535,1540
,|1540,1541
EOMI|1542,1546
.|1546,1547
Conjunctiva|1548,1559
pink|1560,1564
,|1564,1565
no|1566,1568
<EOL>|1568,1569
pallor|1569,1575
or|1576,1578
cyanosis|1579,1587
of|1588,1590
the|1591,1594
oral|1595,1599
mucosa|1600,1606
<EOL>|1606,1607
NECK|1607,1611
:|1611,1612
Supple|1613,1619
with|1620,1624
no|1625,1627
JVD|1628,1631
<EOL>|1631,1632
CARDIAC|1632,1639
:|1639,1640
RRR|1641,1644
normal|1645,1651
S1|1652,1654
/|1654,1655
S2|1655,1657
.|1657,1658
No|1659,1661
thrills|1662,1669
,|1669,1670
lifts|1671,1676
.|1676,1677
<EOL>|1679,1680
LUNGS|1680,1685
:|1685,1686
CTAB|1687,1691
.|1691,1692
No|1693,1695
crackles|1696,1704
,|1704,1705
wheezes|1706,1713
or|1714,1716
rhonchi|1717,1724
.|1724,1725
<EOL>|1727,1728
ABDOMEN|1728,1735
:|1735,1736
Soft|1737,1741
,|1741,1742
NTND|1743,1747
.|1747,1748
<EOL>|1749,1750
EXTREMITIES|1750,1761
:|1761,1762
No|1763,1765
_|1766,1767
_|1767,1768
_|1768,1769
edema|1770,1775
<EOL>|1775,1776
PULSES|1776,1782
:|1782,1783
_|1784,1785
_|1785,1786
_|1786,1787
and|1788,1791
DP|1792,1794
palpable|1795,1803
on|1804,1806
the|1807,1810
right|1811,1816
side|1817,1821
.|1821,1822
Did|1823,1826
not|1827,1830
take|1831,1835
<EOL>|1835,1836
bandage|1836,1843
down|1844,1848
for|1849,1852
exam|1853,1857
as|1858,1860
podiatry|1861,1869
had|1870,1873
just|1874,1878
dressed|1879,1886
.|1886,1887
<EOL>|1887,1888
<EOL>|1888,1889
Per|1889,1892
podiatry|1893,1901
exam|1902,1906
(|1907,1908
_|1908,1909
_|1909,1910
_|1910,1911
)|1911,1912
[|1913,1914
See|1914,1917
attached|1918,1926
picture|1927,1934
on|1935,1937
OMR|1938,1941
]|1941,1942
<EOL>|1942,1943
_|1943,1944
_|1944,1945
_|1945,1946
pulses|1947,1953
palpable|1954,1962
b|1963,1964
/|1964,1965
l|1965,1966
.|1966,1967
CFT|1968,1971
<|1972,1973
3|1973,1974
sec|1975,1978
to|1979,1981
digits|1982,1988
<EOL>|1988,1989
bilaterally|1989,2000
.|2000,2001
There|2002,2007
is|2008,2010
a|2011,2012
L|2013,2014
hallux|2015,2021
wound|2022,2027
present|2028,2035
at|2036,2038
the|2039,2042
medial|2043,2049
<EOL>|2049,2050
aspect|2050,2056
of|2057,2059
the|2060,2063
toe|2064,2067
at|2068,2070
the|2071,2074
level|2075,2080
of|2081,2083
the|2084,2087
IPJ|2088,2091
.|2091,2092
Wound|2093,2098
has|2099,2102
eschar|2103,2109
over|2110,2114
<EOL>|2114,2115
top|2115,2118
of|2119,2121
the|2122,2125
base|2126,2130
w|2131,2132
/|2132,2133
surrounding|2134,2145
hyperkeratotic|2146,2160
skin|2161,2165
and|2166,2169
<EOL>|2169,2170
surrounding|2170,2181
erythema|2182,2190
.|2190,2191
There|2192,2197
is|2198,2200
no|2201,2203
malodor|2204,2211
or|2212,2214
proximal|2215,2223
streaking|2224,2233
<EOL>|2233,2234
present|2234,2241
.|2241,2242
Once|2243,2247
the|2248,2251
wound|2252,2257
was|2258,2261
debrided|2262,2270
and|2271,2274
the|2275,2278
eschar|2279,2285
was|2286,2289
<EOL>|2290,2291
deroofed|2291,2299
,|2299,2300
<EOL>|2300,2301
there|2301,2306
is|2307,2309
fibrotic|2310,2318
skin|2319,2323
at|2324,2326
the|2327,2330
base|2331,2335
of|2336,2338
the|2339,2342
wound|2343,2348
.|2348,2349
It|2350,2352
does|2353,2357
not|2358,2361
<EOL>|2361,2362
probe|2362,2367
deep|2368,2372
to|2373,2375
bone|2376,2380
.|2380,2381
2cc|2382,2385
of|2386,2388
purulent|2389,2397
drainage|2398,2406
was|2407,2410
expressed|2411,2420
from|2421,2425
<EOL>|2425,2426
wound.|2426,2432
Wound|2433,2438
is|2439,2441
extremely|2442,2451
TTP|2452,2455
.|2455,2456
Gross|2457,2462
sensation|2463,2472
is|2473,2475
intact|2476,2482
to|2483,2485
b|2486,2487
/|2487,2488
l|2488,2489
<EOL>|2489,2490
lower|2490,2495
extremities|2496,2507
.|2507,2508
MMT|2509,2512
_|2513,2514
_|2514,2515
_|2515,2516
to|2517,2519
all|2520,2523
_|2524,2525
_|2525,2526
_|2526,2527
muscle|2528,2534
groups|2535,2541
crossing|2542,2550
the|2551,2554
<EOL>|2554,2555
ankle|2555,2560
jt|2561,2563
.|2563,2564
No|2565,2567
gross|2568,2573
deformities|2574,2585
noted|2586,2591
.|2591,2592
<EOL>|2593,2594
<EOL>|2595,2596
Pertinent|2596,2605
Results|2606,2613
:|2613,2614
<EOL>|2614,2615
ADMISSION|2615,2624
LABS|2625,2629
<EOL>|2629,2630
=|2630,2631
=|2631,2632
=|2632,2633
=|2633,2634
=|2634,2635
=|2635,2636
=|2636,2637
=|2637,2638
=|2638,2639
=|2639,2640
=|2640,2641
=|2641,2642
=|2642,2643
=|2643,2644
<EOL>|2644,2645
_|2645,2646
_|2646,2647
_|2647,2648
12|2649,2651
:|2651,2652
50AM|2652,2656
BLOOD|2657,2662
WBC|2663,2666
-|2666,2667
12|2667,2669
.|2669,2670
7|2670,2671
*|2671,2672
RBC|2673,2676
-|2676,2677
4|2677,2678
.|2678,2679
34|2679,2681
Hgb|2682,2685
-|2685,2686
14.4|2686,2690
Hct|2691,2694
-|2694,2695
41.7|2695,2699
<EOL>|2700,2701
MCV|2701,2704
-|2704,2705
96|2705,2707
MCH|2708,2711
-|2711,2712
33|2712,2714
.|2714,2715
2|2715,2716
*|2716,2717
MCHC|2718,2722
-|2722,2723
34.5|2723,2727
RDW|2728,2731
-|2731,2732
11.8|2732,2736
RDWSD|2737,2742
-|2742,2743
41.3|2743,2747
Plt|2748,2751
_|2752,2753
_|2753,2754
_|2754,2755
<EOL>|2755,2756
_|2756,2757
_|2757,2758
_|2758,2759
12|2760,2762
:|2762,2763
50AM|2763,2767
BLOOD|2768,2773
Glucose|2774,2781
-|2781,2782
318|2782,2785
*|2785,2786
UreaN|2787,2792
-|2792,2793
21|2793,2795
*|2795,2796
Creat|2797,2802
-|2802,2803
1.1|2803,2806
Na|2807,2809
-|2809,2810
134|2810,2813
*|2813,2814
<EOL>|2815,2816
K|2816,2817
-|2817,2818
4.2|2818,2821
Cl|2822,2824
-|2824,2825
92|2825,2827
*|2827,2828
HCO3|2829,2833
-|2833,2834
19|2834,2836
*|2836,2837
AnGap|2838,2843
-|2843,2844
23|2844,2846
*|2846,2847
<EOL>|2847,2848
_|2848,2849
_|2849,2850
_|2850,2851
12|2852,2854
:|2854,2855
50AM|2855,2859
BLOOD|2860,2865
cTropnT|2866,2873
-|2873,2874
<|2874,2875
0|2875,2876
.|2876,2877
01|2877,2879
<EOL>|2879,2880
_|2880,2881
_|2881,2882
_|2882,2883
06|2884,2886
:|2886,2887
00AM|2887,2891
BLOOD|2892,2897
cTropnT|2898,2905
-|2905,2906
<|2906,2907
0|2907,2908
.|2908,2909
01|2909,2911
<EOL>|2911,2912
_|2912,2913
_|2913,2914
_|2914,2915
11|2916,2918
:|2918,2919
40AM|2919,2923
BLOOD|2924,2929
cTropnT|2930,2937
-|2937,2938
<|2938,2939
0|2939,2940
.|2940,2941
01|2941,2943
<EOL>|2943,2944
_|2944,2945
_|2945,2946
_|2946,2947
05|2948,2950
:|2950,2951
20PM|2951,2955
BLOOD|2956,2961
CK|2962,2964
-|2964,2965
MB|2965,2967
-|2967,2968
1|2968,2969
cTropnT|2970,2977
-|2977,2978
<|2978,2979
0|2979,2980
.|2980,2981
01|2981,2983
<EOL>|2983,2984
_|2984,2985
_|2985,2986
_|2986,2987
05|2988,2990
:|2990,2991
20PM|2991,2995
BLOOD|2996,3001
Albumin|3002,3009
-|3009,3010
3.5|3010,3013
Calcium|3014,3021
-|3021,3022
8.6|3022,3025
Phos|3026,3030
-|3030,3031
3.6|3031,3034
Mg|3035,3037
-|3037,3038
1.8|3038,3041
<EOL>|3041,3042
_|3042,3043
_|3043,3044
_|3044,3045
05|3046,3048
:|3048,3049
20PM|3049,3053
BLOOD|3054,3059
%|3060,3061
HbA1c|3061,3066
-|3066,3067
12|3067,3069
.|3069,3070
0|3070,3071
*|3071,3072
eAG|3073,3076
-|3076,3077
298|3077,3080
*|3080,3081
<EOL>|3081,3082
_|3082,3083
_|3083,3084
_|3084,3085
12|3086,3088
:|3088,3089
50AM|3089,3093
BLOOD|3094,3099
CRP|3100,3103
-|3103,3104
36|3104,3106
.|3106,3107
4|3107,3108
*|3108,3109
<EOL>|3109,3110
_|3110,3111
_|3111,3112
_|3112,3113
12|3114,3116
:|3116,3117
50AM|3117,3121
BLOOD|3122,3127
ASA|3128,3131
-|3131,3132
NEG|3132,3135
Acetmnp|3136,3143
-|3143,3144
NEG|3144,3147
Tricycl|3148,3155
-|3155,3156
NEG|3156,3159
<EOL>|3159,3160
<EOL>|3160,3161
STUDIES|3161,3168
<EOL>|3168,3169
=|3169,3170
=|3170,3171
=|3171,3172
=|3172,3173
=|3173,3174
=|3174,3175
=|3175,3176
<EOL>|3176,3177
_|3177,3178
_|3178,3179
_|3179,3180
Coronary|3181,3189
Angiogram|3190,3199
<EOL>|3199,3200
Coronary|3200,3208
Anatomy|3209,3216
<EOL>|3216,3217
Dominance|3217,3226
:|3226,3227
Right|3228,3233
<EOL>|3233,3234
*|3234,3235
Left|3236,3240
Main|3241,3245
Coronary|3246,3254
Artery|3255,3261
<EOL>|3261,3262
The|3262,3265
LMCA|3266,3270
is|3271,3273
.|3273,3274
<EOL>|3274,3275
*|3275,3276
Left|3277,3281
Anterior|3282,3290
Descending|3291,3301
<EOL>|3301,3302
The|3302,3305
LAD|3306,3309
has|3310,3313
diffuse|3314,3321
60|3322,3324
%|3324,3325
in|3326,3328
-|3328,3329
stent|3329,3334
restenosis|3335,3345
with|3346,3350
patent|3351,3357
LIMA|3358,3362
to|3363,3365
<EOL>|3366,3367
distal|3367,3373
vessel|3374,3380
.|3380,3381
<EOL>|3381,3382
The|3382,3385
_|3386,3387
_|3387,3388
_|3388,3389
Diagonal|3390,3398
is|3399,3401
small|3402,3407
and|3408,3411
diffusely|3412,3421
diseased|3422,3430
.|3430,3431
<EOL>|3431,3432
*|3432,3433
Circumflex|3434,3444
<EOL>|3444,3445
The|3445,3448
Circumflex|3449,3459
is|3460,3462
occluded|3463,3471
after|3472,3477
a|3478,3479
small|3480,3485
OM1|3486,3489
.|3489,3490
There|3491,3496
is|3497,3499
a|3500,3501
patent|3502,3508
<EOL>|3509,3510
SVG|3510,3513
to|3514,3516
OM2|3517,3520
.|3520,3521
<EOL>|3521,3522
*|3522,3523
Right|3524,3529
Coronary|3530,3538
Artery|3539,3545
<EOL>|3545,3546
The|3546,3549
RCA|3550,3553
has|3554,3557
focal|3558,3563
mid|3564,3567
50|3568,3570
%|3570,3571
stenosis|3572,3580
.|3580,3581
<EOL>|3581,3582
SVG|3582,3585
to|3586,3588
OM|3589,3591
patent|3592,3598
.|3598,3599
<EOL>|3599,3600
LIMA|3600,3604
to|3605,3607
LAD|3608,3611
patent|3612,3618
.|3618,3619
<EOL>|3619,3620
Intra-procedural|3620,3636
Complications|3637,3650
:|3650,3651
None|3652,3656
<EOL>|3656,3657
Impressions|3657,3668
:|3668,3669
<EOL>|3669,3670
1.|3670,3672
three|3673,3678
vessel|3679,3685
CAD|3686,3689
.|3689,3690
<EOL>|3690,3691
2.|3691,3693
Patent|3694,3700
SVG|3701,3704
to|3705,3707
OM|3708,3710
and|3711,3714
LIMA|3715,3719
to|3720,3722
LAD|3723,3726
.|3726,3727
<EOL>|3727,3728
Recommendations|3728,3743
<EOL>|3743,3744
1.|3744,3746
Medical|3747,3754
therapy|3755,3762
.|3762,3763
<EOL>|3763,3764
<EOL>|3764,3765
Pharmacological|3765,3780
MIBI|3781,3785
_|3786,3787
_|3787,3788
_|3788,3789
<EOL>|3789,3790
IMPRESSION|3790,3800
:|3800,3801
<EOL>|3802,3803
<EOL>|3805,3806
1.|3806,3808
Reversible|3809,3819
,|3819,3820
medium|3821,3827
sized|3828,3833
,|3833,3834
moderate|3835,3843
severity|3844,3852
perfusion|3853,3862
defect|3863,3869
<EOL>|3870,3871
involving|3871,3880
the|3881,3884
<EOL>|3885,3886
LAD|3886,3889
territory|3890,3899
.|3899,3900
<EOL>|3901,3902
<EOL>|3904,3905
2.|3905,3907
Normal|3908,3914
left|3915,3919
ventricular|3920,3931
cavity|3932,3938
size|3939,3943
and|3944,3947
systolic|3948,3956
function|3957,3965
.|3965,3966
<EOL>|3969,3970
<EOL>|3972,3973
Compared|3973,3981
to|3982,3984
the|3985,3988
prior|3989,3994
study|3995,4000
of|4001,4003
_|4004,4005
_|4005,4006
_|4006,4007
,|4007,4008
the|4009,4012
perfusion|4013,4022
defect|4023,4029
<EOL>|4030,4031
is|4031,4033
new|4034,4037
.|4037,4038
<EOL>|4039,4040
<EOL>|4042,4043
<EOL>|4043,4044
ECHO|4044,4048
_|4049,4050
_|4050,4051
_|4051,4052
<EOL>|4052,4053
LEFT|4053,4057
ATRIUM|4058,4064
:|4064,4065
Normal|4066,4072
LA|4073,4075
volume|4076,4082
index|4083,4088
.|4088,4089
<EOL>|4090,4091
<EOL>|4091,4092
LEFT|4092,4096
VENTRICLE|4097,4106
:|4106,4107
Normal|4108,4114
LV|4115,4117
wall|4118,4122
thickness|4123,4132
,|4132,4133
cavity|4134,4140
size|4141,4145
,|4145,4146
and|4147,4150
<EOL>|4151,4152
regional|4152,4160
/|4160,4161
global|4161,4167
systolic|4168,4176
function|4177,4185
(|4186,4187
biplane|4187,4194
LVEF|4195,4199
>|4199,4200
55|4200,4202
%|4202,4203
)|4203,4204
.|4204,4205
Doppler|4206,4213
<EOL>|4214,4215
parameters|4215,4225
are|4226,4229
most|4230,4234
consistent|4235,4245
with|4246,4250
normal|4251,4257
LV|4258,4260
diastolic|4261,4270
<EOL>|4271,4272
function|4272,4280
.|4280,4281
<EOL>|4282,4283
<EOL>|4283,4284
RIGHT|4284,4289
VENTRICLE|4290,4299
:|4299,4300
Normal|4301,4307
RV|4308,4310
chamber|4311,4318
size|4319,4323
and|4324,4327
free|4328,4332
wall|4333,4337
motion|4338,4344
.|4344,4345
<EOL>|4346,4347
Paradoxic|4347,4356
septal|4357,4363
motion|4364,4370
consistent|4371,4381
with|4382,4386
prior|4387,4392
cardiac|4393,4400
surgery|4401,4408
.|4408,4409
<EOL>|4410,4411
<EOL>|4411,4412
AORTA|4412,4417
:|4417,4418
Normal|4419,4425
diameter|4426,4434
of|4435,4437
aorta|4438,4443
at|4444,4446
the|4447,4450
sinus|4451,4456
,|4456,4457
ascending|4458,4467
and|4468,4471
arch|4472,4476
<EOL>|4477,4478
levels|4478,4484
.|4484,4485
<EOL>|4486,4487
<EOL>|4487,4488
AORTIC|4488,4494
VALVE|4495,4500
:|4500,4501
Normal|4502,4508
aortic|4509,4515
valve|4516,4521
leaflets|4522,4530
(|4531,4532
3|4532,4533
)|4533,4534
.|4534,4535
No|4536,4538
AS|4539,4541
.|4541,4542
No|4543,4545
AR|4546,4548
.|4548,4549
<EOL>|4550,4551
<EOL>|4551,4552
MITRAL|4552,4558
VALVE|4559,4564
:|4564,4565
Normal|4566,4572
mitral|4573,4579
valve|4580,4585
leaflets|4586,4594
with|4595,4599
trivial|4600,4607
MR|4608,4610
.|4610,4611
<EOL>|4612,4613
_|4613,4614
_|4614,4615
_|4615,4616
mitral|4617,4623
valve|4624,4629
supporting|4630,4640
structures|4641,4651
.|4651,4652
No|4653,4655
MS|4656,4658
.|4658,4659
<EOL>|4660,4661
<EOL>|4661,4662
_|4662,4663
_|4663,4664
_|4664,4665
VALVE|4666,4671
:|4671,4672
Normal|4673,4679
tricuspid|4680,4689
valve|4690,4695
leaflets|4696,4704
with|4705,4709
trivial|4710,4717
<EOL>|4718,4719
TR|4719,4721
.|4721,4722
Normal|4723,4729
PA|4730,4732
systolic|4733,4741
pressure|4742,4750
.|4750,4751
<EOL>|4752,4753
<EOL>|4753,4754
PULMONIC|4754,4762
VALVE|4763,4768
/|4768,4769
PULMONARY|4769,4778
ARTERY|4779,4785
:|4785,4786
Pulmonic|4787,4795
valve|4796,4801
not|4802,4805
visualized|4806,4816
.|4816,4817
<EOL>|4818,4819
No|4819,4821
PS|4822,4824
.|4824,4825
Physiologic|4826,4837
PR|4838,4840
.|4840,4841
<EOL>|4842,4843
<EOL>|4843,4844
PERICARDIUM|4844,4855
:|4855,4856
No|4857,4859
pericardial|4860,4871
effusion|4872,4880
.|4880,4881
<EOL>|4884,4885
Conclusions|4885,4896
<EOL>|4899,4900
The|4901,4904
left|4905,4909
atrial|4910,4916
volume|4917,4923
index|4924,4929
is|4930,4932
normal|4933,4939
.|4939,4940
Normal|4941,4947
left|4948,4952
ventricular|4953,4964
<EOL>|4965,4966
wall|4966,4970
thickness|4971,4980
,|4980,4981
cavity|4982,4988
size|4989,4993
,|4993,4994
and|4995,4998
regional|4999,5007
/|5007,5008
global|5008,5014
systolic|5015,5023
<EOL>|5024,5025
function|5025,5033
(|5034,5035
biplane|5035,5042
LVEF|5043,5047
=|5048,5049
63|5050,5052
%|5053,5054
)|5054,5055
.|5055,5056
Doppler|5057,5064
parameters|5065,5075
are|5076,5079
most|5080,5084
<EOL>|5085,5086
consistent|5086,5096
with|5097,5101
normal|5102,5108
left|5109,5113
ventricular|5114,5125
diastolic|5126,5135
function|5136,5144
.|5144,5145
<EOL>|5146,5147
Right|5147,5152
ventricular|5153,5164
chamber|5165,5172
size|5173,5177
and|5178,5181
free|5182,5186
wall|5187,5191
motion|5192,5198
are|5199,5202
normal|5203,5209
.|5209,5210
<EOL>|5211,5212
The|5212,5215
diameters|5216,5225
of|5226,5228
aorta|5229,5234
at|5235,5237
the|5238,5241
sinus|5242,5247
,|5247,5248
ascending|5249,5258
and|5259,5262
arch|5263,5267
levels|5268,5274
<EOL>|5275,5276
are|5276,5279
normal|5280,5286
.|5286,5287
The|5288,5291
aortic|5292,5298
valve|5299,5304
leaflets|5305,5313
(|5314,5315
3|5315,5316
)|5316,5317
appear|5318,5324
structurally|5325,5337
<EOL>|5338,5339
normal|5339,5345
with|5346,5350
good|5351,5355
leaflet|5356,5363
excursion|5364,5373
and|5374,5377
no|5378,5380
aortic|5381,5387
stenosis|5388,5396
or|5397,5399
<EOL>|5400,5401
aortic|5401,5407
regurgitation|5408,5421
.|5421,5422
The|5423,5426
mitral|5427,5433
valve|5434,5439
appears|5440,5447
structurally|5448,5460
<EOL>|5461,5462
normal|5462,5468
with|5469,5473
trivial|5474,5481
mitral|5482,5488
regurgitation|5489,5502
.|5502,5503
The|5504,5507
estimated|5508,5517
<EOL>|5518,5519
pulmonary|5519,5528
artery|5529,5535
systolic|5536,5544
pressure|5545,5553
is|5554,5556
normal|5557,5563
.|5563,5564
There|5565,5570
is|5571,5573
no|5574,5576
<EOL>|5577,5578
pericardial|5578,5589
effusion|5590,5598
.|5598,5599
<EOL>|5600,5601
<EOL>|5601,5602
IMPRESSION|5603,5613
:|5613,5614
<EOL>|5615,5616
1|5617,5618
)|5618,5619
Normal|5620,5626
biventricular|5627,5640
regional|5641,5649
/|5649,5650
global|5650,5656
systolic|5657,5665
function|5666,5674
.|5674,5675
<EOL>|5676,5677
<EOL>|5677,5678
Compared|5679,5687
with|5688,5692
the|5693,5696
prior|5697,5702
study|5703,5708
(|5709,5710
images|5710,5716
reviewed|5717,5725
)|5725,5726
of|5727,5729
_|5730,5731
_|5731,5732
_|5732,5733
,|5733,5734
<EOL>|5735,5736
no|5736,5738
clinically|5739,5749
significant|5750,5761
change|5762,5768
noted|5769,5774
<EOL>|5775,5776
<EOL>|5776,5777
DISCHARGE|5777,5786
LABS|5787,5791
<EOL>|5791,5792
=|5792,5793
=|5793,5794
=|5794,5795
=|5795,5796
=|5796,5797
=|5797,5798
=|5798,5799
=|5799,5800
=|5800,5801
=|5801,5802
=|5802,5803
=|5803,5804
=|5804,5805
=|5805,5806
<EOL>|5806,5807
_|5807,5808
_|5808,5809
_|5809,5810
06|5811,5813
:|5813,5814
10AM|5814,5818
BLOOD|5819,5824
WBC|5825,5828
-|5828,5829
7.7|5829,5832
RBC|5833,5836
-|5836,5837
3|5837,5838
.|5838,5839
53|5839,5841
*|5841,5842
Hgb|5843,5846
-|5846,5847
11.6|5847,5851
Hct|5852,5855
-|5855,5856
33|5856,5858
.|5858,5859
8|5859,5860
*|5860,5861
<EOL>|5862,5863
MCV|5863,5866
-|5866,5867
96|5867,5869
MCH|5870,5873
-|5873,5874
32|5874,5876
.|5876,5877
9|5877,5878
*|5878,5879
MCHC|5880,5884
-|5884,5885
34.3|5885,5889
RDW|5890,5893
-|5893,5894
11.7|5894,5898
RDWSD|5899,5904
-|5904,5905
40.6|5905,5909
Plt|5910,5913
_|5914,5915
_|5915,5916
_|5916,5917
<EOL>|5917,5918
_|5918,5919
_|5919,5920
_|5920,5921
06|5922,5924
:|5924,5925
10AM|5925,5929
BLOOD|5930,5935
Glucose|5936,5943
-|5943,5944
245|5944,5947
*|5947,5948
UreaN|5949,5954
-|5954,5955
12|5955,5957
Creat|5958,5963
-|5963,5964
1.0|5964,5967
Na|5968,5970
-|5970,5971
140|5971,5974
<EOL>|5975,5976
K|5976,5977
-|5977,5978
4.3|5978,5981
Cl|5982,5984
-|5984,5985
101|5985,5988
HCO3|5989,5993
-|5993,5994
25|5994,5996
AnGap|5997,6002
-|6002,6003
14|6003,6005
<EOL>|6005,6006
_|6006,6007
_|6007,6008
_|6008,6009
02|6010,6012
:|6012,6013
45AM|6013,6017
BLOOD|6018,6023
ALT|6024,6027
-|6027,6028
14|6028,6030
AST|6031,6034
-|6034,6035
17|6035,6037
AlkPhos|6038,6045
-|6045,6046
50|6046,6048
TotBili|6049,6056
-|6056,6057
0.4|6057,6060
<EOL>|6060,6061
_|6061,6062
_|6062,6063
_|6063,6064
06|6065,6067
:|6067,6068
10AM|6068,6072
BLOOD|6073,6078
Calcium|6079,6086
-|6086,6087
8|6087,6088
.|6088,6089
0|6089,6090
*|6090,6091
Phos|6092,6096
-|6096,6097
2|6097,6098
.|6098,6099
6|6099,6100
*|6100,6101
Mg|6102,6104
-|6104,6105
1.|6105,6107
_|6107,6108
_|6108,6109
_|6109,6110
year|6111,6115
old|6116,6119
female|6120,6126
with|6127,6131
CAD|6132,6135
(|6135,6136
s|6136,6137
/|6137,6138
p|6138,6139
BMS|6140,6143
proximal|6144,6152
-|6152,6153
LAD|6153,6156
_|6157,6158
_|6158,6159
_|6159,6160
,|6160,6161
DES|6162,6165
to|6166,6168
<EOL>|6169,6170
mid|6170,6173
LAD|6174,6177
_|6178,6179
_|6179,6180
_|6180,6181
,|6181,6182
DES|6183,6186
to|6187,6189
edge|6190,6194
ISR|6195,6198
of|6199,6201
mid|6202,6205
LAD|6206,6209
DES|6210,6213
and|6214,6217
stenosis|6218,6226
distal|6227,6233
<EOL>|6234,6235
to|6235,6237
stent|6238,6243
_|6244,6245
_|6245,6246
_|6246,6247
,|6247,6248
DES|6249,6252
to|6253,6255
_|6256,6257
_|6257,6258
_|6258,6259
,|6259,6260
s|6261,6262
/|6262,6263
p|6263,6264
3|6265,6266
v|6267,6268
CABG|6269,6273
LIMA|6274,6278
-|6278,6279
LAD|6279,6282
,|6282,6283
<EOL>|6284,6285
SVG|6285,6288
-|6288,6289
OM1|6289,6292
,|6292,6293
SVG|6294,6297
-|6297,6298
D1|6298,6300
(|6300,6301
occluded|6301,6309
)|6309,6310
_|6311,6312
_|6312,6313
_|6313,6314
,|6314,6315
HFpEF|6316,6321
,|6321,6322
IDDM|6323,6327
,|6327,6328
HTN|6329,6332
who|6333,6336
<EOL>|6337,6338
presented|6338,6347
with|6348,6352
several|6353,6360
days|6361,6365
atypical|6366,6374
chest|6375,6380
pain|6381,6385
both|6386,6390
with|6391,6395
<EOL>|6396,6397
exertion|6397,6405
and|6406,6409
at|6410,6412
rest|6413,6417
,|6417,6418
with|6419,6423
mild|6424,6428
T|6429,6430
wave|6431,6435
deepening|6436,6445
but|6446,6449
no|6450,6452
other|6453,6458
<EOL>|6459,6460
EKG|6460,6463
changes|6464,6471
or|6472,6474
troponin|6475,6483
.|6483,6484
She|6485,6488
also|6489,6493
presented|6494,6503
with|6504,6508
mild|6509,6513
DKA|6514,6517
and|6518,6521
<EOL>|6522,6523
diabetic|6523,6531
foot|6532,6536
ulcer|6537,6542
.|6542,6543
She|6544,6547
had|6548,6551
a|6552,6553
stress|6554,6560
test|6561,6565
with|6566,6570
reversible|6571,6581
<EOL>|6582,6583
ischemia|6583,6591
in|6592,6594
the|6595,6598
LAD|6599,6602
territory|6603,6612
(|6613,6614
_|6614,6615
_|6615,6616
_|6616,6617
)|6617,6618
and|6619,6622
went|6623,6627
to|6628,6630
cardiac|6631,6638
<EOL>|6639,6640
catheterization|6640,6655
_|6656,6657
_|6657,6658
_|6658,6659
which|6660,6665
showed|6666,6672
stable|6673,6679
disease|6680,6687
and|6688,6691
no|6692,6694
new|6695,6698
<EOL>|6699,6700
obstructive|6700,6711
lesions|6712,6719
.|6719,6720
Overall|6721,6728
her|6729,6732
chest|6733,6738
pain|6739,6743
was|6744,6747
felt|6748,6752
to|6753,6755
have|6756,6760
<EOL>|6761,6762
been|6762,6766
either|6767,6773
musculoskeletal|6774,6789
or|6790,6792
demand|6793,6799
in|6800,6802
the|6803,6806
setting|6807,6814
of|6815,6817
DKA|6818,6821
and|6822,6825
<EOL>|6826,6827
diabetic|6827,6835
foot|6836,6840
ulcer|6841,6846
.|6846,6847
She|6848,6851
was|6852,6855
discharged|6856,6866
on|6867,6869
ASA|6870,6873
81|6874,6876
,|6876,6877
atorvastatin|6878,6890
<EOL>|6891,6892
80|6892,6894
,|6894,6895
Metoprolol|6896,6906
XL|6907,6909
100mg|6910,6915
daily|6916,6921
.|6921,6922
<EOL>|6923,6924
<EOL>|6924,6925
#|6925,6926
DKA|6926,6929
/|6929,6930
IDDM|6930,6934
:|6934,6935
Patient|6936,6943
presented|6944,6953
with|6954,6958
anion|6959,6964
gap|6965,6968
metabolic|6969,6978
acidosis|6979,6987
<EOL>|6988,6989
and|6989,6992
felt|6993,6997
to|6998,7000
be|7001,7003
in|7004,7006
mild|7007,7011
DKA|7012,7015
.|7015,7016
She|7017,7020
had|7021,7024
insulin|7025,7032
gtt|7033,7036
in|7037,7039
the|7040,7043
ED|7044,7046
but|7047,7050
<EOL>|7051,7052
was|7052,7055
rapidly|7056,7063
switched|7064,7072
to|7073,7075
subcutaneous|7076,7088
insulin|7089,7096
.|7096,7097
Her|7098,7101
A1c|7102,7105
returned|7106,7114
<EOL>|7115,7116
at|7116,7118
12|7119,7121
%|7121,7122
,|7122,7123
which|7124,7129
is|7130,7132
the|7133,7136
highest|7137,7144
it|7145,7147
has|7148,7151
been|7152,7156
recorded|7157,7165
for|7166,7169
her|7170,7173
in|7174,7176
our|7177,7180
<EOL>|7181,7182
records|7182,7189
.|7189,7190
She|7191,7194
had|7195,7198
followed|7199,7207
with|7208,7212
_|7213,7214
_|7214,7215
_|7215,7216
previously|7217,7227
and|7228,7231
was|7232,7235
<EOL>|7236,7237
on|7237,7239
canagliflozin|7240,7253
and|7254,7257
glipizide|7258,7267
as|7268,7270
well|7271,7275
as|7276,7278
SC|7279,7281
insulin|7282,7289
prior|7290,7295
to|7296,7298
<EOL>|7299,7300
admission|7300,7309
.|7309,7310
However|7311,7318
,|7318,7319
she|7320,7323
reported|7324,7332
intermittent|7333,7345
adherence|7346,7355
to|7356,7358
her|7359,7362
<EOL>|7363,7364
medications|7364,7375
and|7376,7379
this|7380,7384
was|7385,7388
the|7389,7392
likely|7393,7399
reason|7400,7406
for|7407,7410
her|7411,7414
DKA|7415,7418
.|7418,7419
While|7420,7425
<EOL>|7426,7427
she|7427,7430
was|7431,7434
in|7435,7437
house|7438,7443
the|7444,7447
_|7448,7449
_|7449,7450
_|7450,7451
followed|7452,7460
along|7461,7466
and|7467,7470
she|7471,7474
met|7475,7478
<EOL>|7479,7480
with|7480,7484
a|7485,7486
diabetes|7487,7495
educator|7496,7504
.|7504,7505
Her|7506,7509
canagliflozin|7510,7523
was|7524,7527
stopped|7528,7535
at|7536,7538
<EOL>|7539,7540
discharge|7540,7549
due|7550,7553
to|7554,7556
increased|7557,7566
risk|7567,7571
of|7572,7574
amputation|7575,7585
.|7585,7586
<EOL>|7587,7588
<EOL>|7588,7589
#|7589,7590
Diabetic|7590,7598
foot|7599,7603
ulcer|7604,7609
:|7609,7610
Present|7611,7618
for|7619,7622
at|7623,7625
least|7626,7631
3|7632,7633
weeks|7634,7639
prior|7640,7645
to|7646,7648
<EOL>|7649,7650
admission|7650,7659
.|7659,7660
She|7661,7664
underwent|7665,7674
bedside|7675,7682
debridement|7683,7694
by|7695,7697
Podiatry|7698,7706
in|7707,7709
ED|7710,7712
.|7712,7713
<EOL>|7714,7715
XR|7715,7717
suggested|7718,7727
presence|7728,7736
of|7737,7739
osteomyelitis|7740,7753
.|7754,7755
She|7756,7759
was|7760,7763
maintained|7764,7774
on|7775,7777
<EOL>|7778,7779
vanc|7779,7783
/|7783,7784
cefepime|7784,7792
/|7792,7793
flagyl|7793,7799
in|7800,7802
house|7803,7808
,|7808,7809
and|7810,7813
was|7814,7817
switched|7818,7826
to|7827,7829
cipro|7830,7835
/|7835,7836
clinda|7836,7842
<EOL>|7843,7844
at|7844,7846
discharge|7847,7856
per|7857,7860
podiatry|7861,7869
recs|7870,7874
with|7875,7879
plans|7880,7885
for|7886,7889
close|7890,7895
follow|7896,7902
up|7903,7905
.|7905,7906
<EOL>|7907,7908
Her|7908,7911
wound|7912,7917
swab|7918,7922
at|7923,7925
time|7926,7930
of|7931,7933
discharge|7934,7943
was|7944,7947
polymicrobial|7948,7961
but|7962,7965
was|7966,7969
<EOL>|7970,7971
growing|7971,7978
Group|7979,7984
B|7985,7986
strep|7987,7992
(|7993,7994
sensitivities|7994,8007
pending|8008,8015
)|8015,8016
and|8017,8020
klebsiella|8021,8031
<EOL>|8032,8033
(|8033,8034
pan|8034,8037
sensitive|8038,8047
)|8047,8048
.|8048,8049
<EOL>|8050,8051
<EOL>|8051,8052
#|8052,8053
Med|8053,8056
noncompliance|8057,8070
:|8070,8071
She|8072,8075
reported|8076,8084
intermittent|8085,8097
medication|8098,8108
<EOL>|8109,8110
compliance|8110,8120
related|8121,8128
to|8129,8131
difficulty|8132,8142
remembering|8143,8154
to|8155,8157
take|8158,8162
her|8163,8166
<EOL>|8167,8168
medications|8168,8179
as|8180,8182
well|8183,8187
as|8188,8190
periods|8191,8198
of|8199,8201
depression|8202,8212
and|8213,8216
stress|8217,8223
where|8224,8229
<EOL>|8230,8231
taking|8231,8237
her|8238,8241
medication|8242,8252
was|8253,8256
not|8257,8260
a|8261,8262
priority|8263,8271
.|8271,8272
She|8273,8276
has|8277,8280
recently|8281,8289
<EOL>|8290,8291
obtained|8291,8299
a|8300,8301
pillbox|8302,8309
and|8310,8313
her|8314,8317
granddaughter|8318,8331
is|8332,8334
helping|8335,8342
her|8343,8346
with|8347,8351
<EOL>|8352,8353
remembering|8353,8364
to|8365,8367
take|8368,8372
her|8373,8376
medications|8377,8388
.|8388,8389
<EOL>|8390,8391
<EOL>|8391,8392
#|8392,8393
HFpEF|8393,8398
:|8398,8399
Metoprolol|8400,8410
as|8411,8413
above|8414,8419
,|8419,8420
continued|8421,8430
torsemide|8431,8440
20mg|8441,8445
and|8446,8449
she|8450,8453
<EOL>|8454,8455
appeared|8455,8463
euvolemic|8464,8473
throughout|8474,8484
admission|8485,8494
.|8494,8495
<EOL>|8496,8497
#|8497,8498
HL|8498,8500
:|8500,8501
Continued|8502,8511
atorvastatin|8512,8524
<EOL>|8524,8525
#|8525,8526
HTN|8526,8529
:|8529,8530
Metoprolol|8531,8541
lowered|8542,8549
to|8550,8552
XL|8553,8555
100mg|8556,8561
daily|8562,8567
,|8567,8568
losartan|8569,8577
kept|8578,8582
at|8583,8585
<EOL>|8586,8587
25mg|8587,8591
daily|8592,8597
.|8597,8598
Imdur|8599,8604
stopped|8605,8612
.|8612,8613
<EOL>|8613,8614
#|8614,8615
COPD|8615,8619
:|8619,8620
Duonebs|8621,8628
q6h|8629,8632
in|8633,8635
house|8636,8641
,|8641,8642
continued|8643,8652
home|8653,8657
inhalers|8658,8666
on|8667,8669
<EOL>|8670,8671
discharge|8671,8680
.|8680,8681
<EOL>|8682,8683
#|8683,8684
Restless|8684,8692
legs|8693,8697
:|8697,8698
continued|8699,8708
ropinerole|8709,8719
<EOL>|8720,8721
<EOL>|8721,8722
Transitional|8722,8734
issues|8735,8741
:|8741,8742
<EOL>|8743,8744
-|8744,8745
Please|8746,8752
follow|8753,8759
up|8760,8762
her|8763,8766
diabetic|8767,8775
foot|8776,8780
ulcer|8781,8786
in|8787,8789
_|8790,8791
_|8791,8792
_|8792,8793
clinic|8794,8800
.|8800,8801
<EOL>|8802,8803
Plan|8803,8807
at|8808,8810
time|8811,8815
of|8816,8818
discharge|8819,8828
was|8829,8832
to|8833,8835
take|8836,8840
to|8841,8843
OR|8844,8846
for|8847,8850
further|8851,8858
surgical|8859,8867
<EOL>|8868,8869
debridement|8869,8880
,|8880,8881
patient|8882,8889
was|8890,8893
discharged|8894,8904
with|8905,8909
cipro|8910,8915
/|8915,8916
clinda|8916,8922
until|8923,8928
<EOL>|8929,8930
Podiatry|8930,8938
follow|8939,8945
up|8946,8948
<EOL>|8949,8950
-|8950,8951
Please|8952,8958
review|8959,8965
her|8966,8969
blood|8970,8975
sugars|8976,8982
at|8983,8985
home|8986,8990
and|8991,8994
continue|8995,9003
to|9004,9006
<EOL>|9007,9008
reinforce|9008,9017
compliance|9018,9028
with|9029,9033
diabetes|9034,9042
medications|9043,9054
.|9054,9055
Her|9056,9059
<EOL>|9060,9061
Canagliflozin|9061,9074
was|9075,9078
stopped|9079,9086
due|9087,9090
to|9091,9093
increased|9094,9103
risk|9104,9108
of|9109,9111
amputation|9112,9122
.|9122,9123
<EOL>|9124,9125
Consider|9125,9133
reintroducing|9134,9147
metformin|9148,9157
as|9158,9160
this|9161,9165
was|9166,9169
stopped|9170,9177
_|9178,9179
_|9179,9180
_|9180,9181
years|9182,9187
ago|9188,9191
<EOL>|9192,9193
for|9193,9196
diarrhea|9197,9205
but|9206,9209
may|9210,9213
be|9214,9216
a|9217,9218
better|9219,9225
option|9226,9232
for|9233,9236
her|9237,9240
.|9240,9241
<EOL>|9242,9243
-|9243,9244
Follow|9245,9251
up|9252,9254
blood|9255,9260
pressures|9261,9270
and|9271,9274
heart|9275,9280
rate|9281,9285
on|9286,9288
the|9289,9292
current|9293,9300
<EOL>|9301,9302
regimen|9302,9309
.|9309,9310
Suspect|9311,9318
that|9319,9323
due|9324,9327
to|9328,9330
noncompliance|9331,9344
her|9345,9348
medications|9349,9360
were|9361,9365
<EOL>|9366,9367
uptitrated|9367,9377
to|9378,9380
higher|9381,9387
doses|9388,9393
than|9394,9398
she|9399,9402
actually|9403,9411
needs|9412,9417
.|9417,9418
We|9419,9421
cut|9422,9425
back|9426,9430
<EOL>|9431,9432
her|9432,9435
Metoprolol|9436,9446
and|9447,9450
stoped|9451,9457
her|9458,9461
imdur|9462,9467
<EOL>|9467,9468
-|9468,9469
Can|9470,9473
restart|9474,9481
imdur|9482,9487
if|9488,9490
requiring|9491,9500
for|9501,9504
chest|9505,9510
pain|9511,9515
on|9516,9518
outpatient|9519,9529
<EOL>|9530,9531
basis|9531,9536
<EOL>|9536,9537
-|9537,9538
Please|9539,9545
continue|9546,9554
to|9555,9557
work|9558,9562
with|9563,9567
patient|9568,9575
on|9576,9578
med|9579,9582
compliance|9583,9593
and|9594,9597
<EOL>|9598,9599
possible|9599,9607
barriers|9608,9616
.|9616,9617
She|9618,9621
denied|9622,9628
depression|9629,9639
with|9640,9644
our|9645,9648
social|9649,9655
worker|9656,9662
<EOL>|9663,9664
but|9664,9667
does|9668,9672
endorse|9673,9680
that|9681,9685
stress|9686,9692
makes|9693,9698
it|9699,9701
hard|9702,9706
to|9707,9709
take|9710,9714
her|9715,9718
<EOL>|9719,9720
medications|9720,9731
.|9731,9732
<EOL>|9733,9734
-|9734,9735
f|9736,9737
/|9737,9738
u|9738,9739
final|9740,9745
wound|9746,9751
swab|9752,9756
cultures|9757,9765
<EOL>|9766,9767
<EOL>|9767,9768
<EOL>|9769,9770
Medications|9770,9781
on|9782,9784
Admission|9785,9794
:|9794,9795
<EOL>|9795,9796
The|9796,9799
Preadmission|9800,9812
Medication|9813,9823
list|9824,9828
is|9829,9831
accurate|9832,9840
and|9841,9844
complete|9845,9853
.|9853,9854
<EOL>|9854,9855
1.|9855,9857
Losartan|9858,9866
Potassium|9867,9876
25|9877,9879
mg|9880,9882
PO|9883,9885
DAILY|9886,9891
<EOL>|9892,9893
2.|9893,9895
MetronidAZOLE|9896,9909
Topical|9910,9917
1|9918,9919
%|9920,9921
Gel|9922,9925
1|9926,9927
Appl|9928,9932
TP|9933,9935
BID|9936,9939
:|9939,9940
PRN|9940,9943
Rosacea|9944,9951
<EOL>|9952,9953
3.|9953,9955
Gabapentin|9956,9966
300|9967,9970
mg|9971,9973
PO|9974,9976
QHS|9977,9980
:|9980,9981
PRN|9981,9984
Headache|9985,9993
<EOL>|9994,9995
4.|9995,9997
Metoprolol|9998,10008
Succinate|10009,10018
XL|10019,10021
250|10022,10025
mg|10026,10028
PO|10029,10031
DAILY|10032,10037
<EOL>|10038,10039
5.|10039,10041
linaGLIPtin|10042,10053
5|10054,10055
mg|10056,10058
oral|10059,10063
DAILY|10064,10069
<EOL>|10070,10071
6.|10071,10073
Atorvastatin|10074,10086
80|10087,10089
mg|10090,10092
PO|10093,10095
QPM|10096,10099
<EOL>|10100,10101
7.|10101,10103
Furosemide|10104,10114
20|10115,10117
mg|10118,10120
PO|10121,10123
DAILY|10124,10129
<EOL>|10130,10131
8.|10131,10133
Isosorbide|10134,10144
Mononitrate|10145,10156
120|10157,10160
mg|10161,10163
PO|10164,10166
DAILY|10167,10172
<EOL>|10173,10174
9.|10174,10176
Nitroglycerin|10177,10190
SL|10191,10193
0.4|10194,10197
mg|10198,10200
SL|10201,10203
Q5MIN|10204,10209
:|10209,10210
PRN|10210,10213
angina|10214,10220
<EOL>|10221,10222
10.|10222,10225
rOPINIRole|10226,10236
0.5|10237,10240
mg|10241,10243
PO|10244,10246
QHS|10247,10250
restless|10251,10259
leg|10260,10263
syndrome|10264,10272
<EOL>|10273,10274
11|10274,10276
.|10276,10277
OxyCODONE|10278,10287
-|10287,10288
-|10288,10289
Acetaminophen|10289,10302
(|10303,10304
5mg|10304,10307
-|10307,10308
325mg|10308,10313
)|10313,10314
1|10315,10316
TAB|10317,10320
PO|10321,10323
Q6H|10324,10327
:|10327,10328
PRN|10328,10331
Pain|10332,10336
-|10337,10338
<EOL>|10339,10340
Severe|10340,10346
<EOL>|10347,10348
12.|10348,10351
Fluticasone|10352,10363
Propionate|10364,10374
110mcg|10375,10381
2|10382,10383
PUFF|10384,10388
IH|10389,10391
BID|10392,10395
<EOL>|10396,10397
13.|10397,10400
Pantoprazole|10401,10413
40|10414,10416
mg|10417,10419
PO|10420,10422
BID|10423,10426
<EOL>|10427,10428
14.|10428,10431
Aspirin|10432,10439
325|10440,10443
mg|10444,10446
PO|10447,10449
DAILY|10450,10455
<EOL>|10456,10457
15.|10457,10460
TraZODone|10461,10470
50|10471,10473
mg|10474,10476
PO|10477,10479
QHS|10480,10483
:|10483,10484
PRN|10484,10487
insomnia|10488,10496
<EOL>|10497,10498
16.|10498,10501
canagliflozin|10502,10515
100|10516,10519
mg|10520,10522
oral|10523,10527
DAILY|10528,10533
<EOL>|10534,10535
17.|10535,10538
albuterol|10539,10548
sulfate|10549,10556
90|10557,10559
mcg|10560,10563
/|10563,10564
actuation|10564,10573
inhalation|10574,10584
Q8H|10585,10588
:|10588,10589
PRN|10589,10592
<EOL>|10593,10594
18.|10594,10597
Lidocaine|10598,10607
5|10608,10609
%|10609,10610
Patch|10611,10616
1|10617,10618
PTCH|10619,10623
TD|10624,10626
QPM|10627,10630
<EOL>|10631,10632
<EOL>|10632,10633
<EOL>|10634,10635
Discharge|10635,10644
Medications|10645,10656
:|10656,10657
<EOL>|10657,10658
1.|10658,10660
Ciprofloxacin|10662,10675
HCl|10676,10679
500|10680,10683
mg|10684,10686
PO|10687,10689
Q12H|10690,10694
<EOL>|10695,10696
RX|10696,10698
*|10699,10700
ciprofloxacin|10700,10713
HCl|10714,10717
500|10718,10721
mg|10722,10724
1|10725,10726
tablet|10727,10733
(|10733,10734
s|10734,10735
)|10735,10736
by|10737,10739
mouth|10740,10745
twice|10746,10751
a|10752,10753
day|10754,10757
<EOL>|10758,10759
Disp|10759,10763
#|10764,10765
*|10765,10766
14|10766,10768
Tablet|10769,10775
Refills|10776,10783
:|10783,10784
*|10784,10785
0|10785,10786
<EOL>|10787,10788
2.|10788,10790
Clindamycin|10792,10803
300|10804,10807
mg|10808,10810
PO|10811,10813
Q6H|10814,10817
<EOL>|10818,10819
RX|10819,10821
*|10822,10823
clindamycin|10823,10834
HCl|10835,10838
300|10839,10842
mg|10843,10845
1|10846,10847
capsule|10848,10855
(|10855,10856
s|10856,10857
)|10857,10858
by|10859,10861
mouth|10862,10867
four|10868,10872
times|10873,10878
per|10879,10882
<EOL>|10883,10884
day|10884,10887
Disp|10888,10892
#|10893,10894
*|10894,10895
28|10895,10897
Capsule|10898,10905
Refills|10906,10913
:|10913,10914
*|10914,10915
0|10915,10916
<EOL>|10917,10918
3.|10918,10920
Glargine|10922,10930
50|10931,10933
Units|10934,10939
Bedtime|10940,10947
<EOL>|10947,10948
Humalog|10948,10955
18|10956,10958
Units|10959,10964
Breakfast|10965,10974
<EOL>|10974,10975
Humalog|10975,10982
18|10983,10985
Units|10986,10991
Lunch|10992,10997
<EOL>|10997,10998
Humalog|10998,11005
18|11006,11008
Units|11009,11014
Dinner|11015,11021
<EOL>|11021,11022
Insulin|11022,11029
SC|11030,11032
Sliding|11033,11040
Scale|11041,11046
using|11047,11052
HUM|11053,11056
Insulin|11057,11064
<EOL>|11065,11066
4.|11066,11068
Metoprolol|11070,11080
Succinate|11081,11090
XL|11091,11093
100|11094,11097
mg|11098,11100
PO|11101,11103
DAILY|11104,11109
<EOL>|11110,11111
RX|11111,11113
*|11114,11115
metoprolol|11115,11125
succinate|11126,11135
100|11136,11139
mg|11140,11142
1|11143,11144
tablet|11145,11151
(|11151,11152
s|11152,11153
)|11153,11154
by|11155,11157
mouth|11158,11163
daily|11164,11169
Disp|11170,11174
<EOL>|11175,11176
#|11176,11177
*|11177,11178
30|11178,11180
Tablet|11181,11187
Refills|11188,11195
:|11195,11196
*|11196,11197
0|11197,11198
<EOL>|11199,11200
5.|11200,11202
albuterol|11204,11213
sulfate|11214,11221
90|11222,11224
mcg|11225,11228
/|11228,11229
actuation|11229,11238
inhalation|11239,11249
Q8H|11250,11253
:|11253,11254
PRN|11254,11257
<EOL>|11259,11260
6.|11260,11262
Aspirin|11264,11271
325|11272,11275
mg|11276,11278
PO|11279,11281
DAILY|11282,11287
<EOL>|11289,11290
7.|11290,11292
Atorvastatin|11294,11306
80|11307,11309
mg|11310,11312
PO|11313,11315
QPM|11316,11319
<EOL>|11321,11322
8.|11322,11324
Fluticasone|11326,11337
Propionate|11338,11348
110mcg|11349,11355
2|11356,11357
PUFF|11358,11362
IH|11363,11365
BID|11366,11369
<EOL>|11371,11372
9.|11372,11374
Furosemide|11376,11386
20|11387,11389
mg|11390,11392
PO|11393,11395
DAILY|11396,11401
<EOL>|11403,11404
10.|11404,11407
Gabapentin|11409,11419
300|11420,11423
mg|11424,11426
PO|11427,11429
QHS|11430,11433
:|11433,11434
PRN|11434,11437
Headache|11438,11446
<EOL>|11448,11449
11.|11449,11452
linaGLIPtin|11454,11465
5|11466,11467
mg|11468,11470
oral|11471,11475
DAILY|11476,11481
<EOL>|11483,11484
12.|11484,11487
Losartan|11489,11497
Potassium|11498,11507
25|11508,11510
mg|11511,11513
PO|11514,11516
DAILY|11517,11522
<EOL>|11524,11525
13.|11525,11528
MetronidAZOLE|11530,11543
Topical|11544,11551
1|11552,11553
%|11554,11555
Gel|11556,11559
1|11560,11561
Appl|11562,11566
TP|11567,11569
BID|11570,11573
:|11573,11574
PRN|11574,11577
Rosacea|11578,11585
<EOL>|11587,11588
14.|11588,11591
Nitroglycerin|11593,11606
SL|11607,11609
0.4|11610,11613
mg|11614,11616
SL|11617,11619
Q5MIN|11620,11625
:|11625,11626
PRN|11626,11629
angina|11630,11636
<EOL>|11638,11639
15.|11639,11642
OxyCODONE|11644,11653
-|11653,11654
-|11654,11655
Acetaminophen|11655,11668
(|11669,11670
5mg|11670,11673
-|11673,11674
325mg|11674,11679
)|11679,11680
1|11681,11682
TAB|11683,11686
PO|11687,11689
Q6H|11690,11693
:|11693,11694
PRN|11694,11697
Pain|11698,11702
<EOL>|11703,11704
-|11704,11705
Severe|11706,11712
<EOL>|11713,11714
RX|11714,11716
*|11717,11718
oxycodone|11718,11727
-|11727,11728
acetaminophen|11728,11741
5|11742,11743
mg|11744,11746
-|11746,11747
325|11747,11750
mg|11751,11753
1|11754,11755
tablet|11756,11762
(|11762,11763
s|11763,11764
)|11764,11765
by|11766,11768
mouth|11769,11774
<EOL>|11775,11776
three|11776,11781
times|11782,11787
daily|11788,11793
Disp|11794,11798
#|11799,11800
*|11800,11801
15|11801,11803
Tablet|11804,11810
Refills|11811,11818
:|11818,11819
*|11819,11820
0|11820,11821
<EOL>|11822,11823
16|11823,11825
.|11825,11826
Pantoprazole|11828,11840
40|11841,11843
mg|11844,11846
PO|11847,11849
BID|11850,11853
<EOL>|11855,11856
17.|11856,11859
rOPINIRole|11861,11871
0.5|11872,11875
mg|11876,11878
PO|11879,11881
QHS|11882,11885
restless|11886,11894
leg|11895,11898
syndrome|11899,11907
<EOL>|11909,11910
18.|11910,11913
TraZODone|11915,11924
50|11925,11927
mg|11928,11930
PO|11931,11933
QHS|11934,11937
:|11937,11938
PRN|11938,11941
insomnia|11942,11950
<EOL>|11952,11953
19|11953,11955
.|11955,11956
HELD|11957,11961
-|11961,11962
canagliflozin|11963,11976
100|11977,11980
mg|11981,11983
oral|11984,11988
DAILY|11989,11994
This|11996,12000
medication|12001,12011
was|12012,12015
<EOL>|12016,12017
held|12017,12021
.|12021,12022
Do|12023,12025
not|12026,12029
restart|12030,12037
canagliflozin|12038,12051
until|12052,12057
you|12058,12061
speak|12062,12067
with|12068,12072
your|12073,12077
<EOL>|12078,12079
endocrinologist|12079,12094
<EOL>|12094,12095
20|12095,12097
.|12097,12098
HELD|12099,12103
-|12103,12104
Lidocaine|12105,12114
5|12115,12116
%|12116,12117
Patch|12118,12123
1|12124,12125
PTCH|12126,12130
TD|12131,12133
QPM|12134,12137
This|12139,12143
medication|12144,12154
was|12155,12158
<EOL>|12159,12160
held|12160,12164
.|12164,12165
Do|12166,12168
not|12169,12172
restart|12173,12180
Lidocaine|12181,12190
5|12191,12192
%|12192,12193
Patch|12194,12199
until|12200,12205
you|12206,12209
speak|12210,12215
with|12216,12220
<EOL>|12221,12222
your|12222,12226
PCP|12227,12230
<EOL>|12230,12231
<EOL>|12231,12232
<EOL>|12233,12234
_|12234,12235
_|12235,12236
_|12236,12237
:|12237,12238
<EOL>|12238,12239
Home|12239,12243
With|12244,12248
Service|12249,12256
<EOL>|12256,12257
<EOL>|12258,12259
Facility|12259,12267
:|12267,12268
<EOL>|12268,12269
_|12269,12270
_|12270,12271
_|12271,12272
<EOL>|12272,12273
<EOL>|12274,12275
Discharge|12275,12284
Diagnosis|12285,12294
:|12294,12295
<EOL>|12295,12296
PRIMARY|12296,12303
<EOL>|12303,12304
=|12304,12305
=|12305,12306
=|12306,12307
=|12307,12308
=|12308,12309
=|12309,12310
=|12310,12311
<EOL>|12311,12312
Diabetic|12312,12320
foot|12321,12325
ulcer|12326,12331
<EOL>|12331,12332
Diabetic|12332,12340
ketoacidosis|12341,12353
<EOL>|12354,12355
Chest|12355,12360
pain|12361,12365
<EOL>|12366,12367
<EOL>|12367,12368
SECONDARY|12368,12377
<EOL>|12377,12378
=|12378,12379
=|12379,12380
=|12380,12381
=|12381,12382
=|12382,12383
=|12383,12384
=|12384,12385
=|12385,12386
=|12386,12387
<EOL>|12387,12388
DIABETES|12388,12396
MELLITUS|12397,12405
(|12406,12407
INSULIN|12407,12414
DEPENDENT|12415,12424
)|12424,12425
<EOL>|12425,12426
COPD|12426,12430
<EOL>|12430,12431
<EOL>|12431,12432
<EOL>|12433,12434
Discharge|12434,12443
Condition|12444,12453
:|12453,12454
<EOL>|12454,12455
Mental|12455,12461
Status|12462,12468
:|12468,12469
Clear|12470,12475
and|12476,12479
coherent|12480,12488
.|12488,12489
<EOL>|12489,12490
Level|12490,12495
of|12496,12498
Consciousness|12499,12512
:|12512,12513
Alert|12514,12519
and|12520,12523
interactive|12524,12535
.|12535,12536
<EOL>|12536,12537
Activity|12537,12545
Status|12546,12552
:|12552,12553
Ambulatory|12554,12564
-|12565,12566
Independent|12567,12578
.|12578,12579
<EOL>|12579,12580
<EOL>|12580,12581
<EOL>|12582,12583
Discharge|12583,12592
Instructions|12593,12605
:|12605,12606
<EOL>|12606,12607
Dear|12607,12611
Ms.|12612,12615
_|12616,12617
_|12617,12618
_|12618,12619
,|12619,12620
<EOL>|12621,12622
<EOL>|12622,12623
It|12623,12625
was|12626,12629
a|12630,12631
pleasure|12632,12640
taking|12641,12647
care|12648,12652
of|12653,12655
you|12656,12659
at|12660,12662
the|12663,12666
_|12667,12668
_|12668,12669
_|12669,12670
<EOL>|12671,12672
_|12672,12673
_|12673,12674
_|12674,12675
!|12675,12676
<EOL>|12678,12679
<EOL>|12679,12680
WHY|12680,12683
WAS|12684,12687
I|12688,12689
IN|12690,12692
THE|12693,12696
HOSPITAL|12697,12705
?|12705,12706
<EOL>|12708,12709
=|12709,12710
=|12710,12711
=|12711,12712
=|12712,12713
=|12713,12714
=|12714,12715
=|12715,12716
=|12716,12717
=|12717,12718
=|12718,12719
=|12719,12720
=|12720,12721
=|12721,12722
=|12722,12723
=|12723,12724
=|12724,12725
=|12725,12726
=|12726,12727
=|12727,12728
=|12728,12729
=|12729,12730
=|12730,12731
=|12731,12732
=|12732,12733
=|12733,12734
=|12734,12735
<EOL>|12737,12738
-|12739,12740
You|12741,12744
were|12745,12749
admitted|12750,12758
because|12759,12766
you|12767,12770
had|12771,12774
chest|12775,12780
pain|12781,12785
.|12785,12786
<EOL>|12787,12788
-|12789,12790
You|12791,12794
also|12795,12799
had|12800,12803
a|12804,12805
process|12806,12813
called|12814,12820
DKA|12821,12824
from|12825,12829
not|12830,12833
taking|12834,12840
enough|12841,12847
<EOL>|12848,12849
insulin|12849,12856
<EOL>|12857,12858
-|12859,12860
You|12861,12864
also|12865,12869
had|12870,12873
a|12874,12875
bad|12876,12879
infection|12880,12889
in|12890,12892
your|12893,12897
foot|12898,12902
.|12902,12903
<EOL>|12904,12905
<EOL>|12905,12906
WHAT|12906,12910
HAPPENED|12911,12919
IN|12920,12922
THE|12923,12926
HOSPITAL|12927,12935
?|12935,12936
<EOL>|12938,12939
=|12939,12940
=|12940,12941
=|12941,12942
=|12942,12943
=|12943,12944
=|12944,12945
=|12945,12946
=|12946,12947
=|12947,12948
=|12948,12949
=|12949,12950
=|12950,12951
=|12951,12952
=|12952,12953
=|12953,12954
=|12954,12955
=|12955,12956
=|12956,12957
=|12957,12958
=|12958,12959
=|12959,12960
=|12960,12961
=|12961,12962
=|12962,12963
=|12963,12964
=|12964,12965
=|12965,12966
=|12966,12967
=|12967,12968
=|12968,12969
<EOL>|12971,12972
-|12973,12974
We|12976,12978
did|12979,12982
several|12983,12990
tests|12991,12996
to|12997,12999
figure|13000,13006
our|13007,13010
if|13011,13013
your|13014,13018
chest|13019,13024
pain|13025,13029
was|13030,13033
<EOL>|13034,13035
caused|13035,13041
by|13042,13044
a|13045,13046
heart|13047,13052
attack|13053,13059
.|13059,13060
The|13061,13064
first|13065,13070
was|13071,13074
a|13075,13076
stress|13077,13083
test|13084,13088
,|13088,13089
which|13090,13095
had|13096,13099
<EOL>|13100,13101
a|13101,13102
positive|13103,13111
results|13112,13119
.|13119,13120
We|13121,13123
then|13124,13128
did|13129,13132
a|13133,13134
procedure|13135,13144
called|13145,13151
a|13152,13153
cardiac|13154,13161
<EOL>|13162,13163
cath|13163,13167
,|13167,13168
which|13169,13174
showed|13175,13181
that|13182,13186
you|13187,13190
did|13191,13194
NOT|13195,13198
have|13199,13203
a|13204,13205
heart|13206,13211
attack|13212,13218
.|13218,13219
<EOL>|13220,13221
-|13222,13223
Our|13224,13227
podiatrists|13228,13239
did|13240,13243
a|13244,13245
debridement|13246,13257
of|13258,13260
your|13261,13265
foot|13266,13270
.|13270,13271
<EOL>|13272,13273
-|13274,13275
We|13276,13278
gave|13279,13283
you|13284,13287
antibiotics|13288,13299
for|13300,13303
your|13304,13308
foot|13309,13313
.|13313,13314
<EOL>|13315,13316
-|13317,13318
We|13319,13321
adjusted|13322,13330
your|13331,13335
insulin|13336,13343
levels|13344,13350
.|13350,13351
<EOL>|13352,13353
<EOL>|13353,13354
WHAT|13354,13358
SHOULD|13359,13365
I|13366,13367
DO|13368,13370
WHEN|13371,13375
I|13376,13377
GO|13378,13380
HOME|13381,13385
?|13385,13386
<EOL>|13388,13389
=|13389,13390
=|13390,13391
=|13391,13392
=|13392,13393
=|13393,13394
=|13394,13395
=|13395,13396
=|13396,13397
=|13397,13398
=|13398,13399
=|13399,13400
=|13400,13401
=|13401,13402
=|13402,13403
=|13403,13404
=|13404,13405
=|13405,13406
=|13406,13407
=|13407,13408
=|13408,13409
=|13409,13410
=|13410,13411
=|13411,13412
=|13412,13413
=|13413,13414
=|13414,13415
=|13415,13416
=|13416,13417
=|13417,13418
=|13418,13419
=|13419,13420
=|13420,13421
<EOL>|13423,13424
-|13424,13425
Take|13426,13430
all|13431,13434
of|13435,13437
your|13438,13442
medications|13443,13454
:|13454,13455
<EOL>|13456,13457
-|13459,13460
Ciproflocaxin|13461,13474
and|13475,13478
Clindamycin|13479,13490
are|13491,13494
antibiotics|13495,13506
you|13507,13510
need|13511,13515
to|13516,13518
<EOL>|13519,13520
take|13520,13524
until|13525,13530
the|13531,13534
podiatrists|13535,13546
tell|13547,13551
you|13552,13555
to|13556,13558
stop|13559,13563
.|13563,13564
You|13566,13569
are|13570,13573
scheduled|13574,13583
<EOL>|13584,13585
to|13585,13587
see|13588,13591
them|13592,13596
_|13597,13598
_|13598,13599
_|13599,13600
<EOL>|13600,13601
-|13603,13604
Your|13605,13609
insulin|13610,13617
regimen|13618,13625
will|13626,13630
be|13631,13633
slightly|13634,13642
different|13643,13652
from|13653,13657
your|13658,13662
<EOL>|13663,13664
old|13664,13667
regimen|13668,13675
.|13675,13676
<EOL>|13677,13678
-|13680,13681
You|13682,13685
need|13686,13690
to|13691,13693
take|13694,13698
aspirin|13699,13706
and|13707,13710
Atorvastatin|13711,13723
every|13724,13729
day|13730,13733
to|13734,13736
<EOL>|13737,13738
prevent|13738,13745
blockages|13746,13755
in|13756,13758
your|13759,13763
heart|13764,13769
from|13770,13774
forming|13775,13782
.|13782,13783
<EOL>|13784,13785
-|13786,13787
You|13788,13791
will|13792,13796
have|13797,13801
many|13802,13806
appointments|13807,13819
in|13820,13822
the|13823,13826
next|13827,13831
week|13832,13836
.|13836,13837
It|13838,13840
is|13841,13843
very|13844,13848
<EOL>|13849,13850
important|13850,13859
that|13860,13864
you|13865,13868
go|13869,13871
to|13872,13874
all|13875,13878
of|13879,13881
these|13882,13887
,|13887,13888
to|13889,13891
help|13892,13896
get|13897,13900
your|13901,13905
health|13906,13912
<EOL>|13913,13914
on|13914,13916
track|13917,13922
!|13922,13923
<EOL>|13924,13925
-|13926,13927
Your|13928,13932
weight|13933,13939
at|13940,13942
discharge|13943,13952
is|13953,13955
79.1|13956,13960
kg|13961,13963
(|13966,13967
174.38|13967,13973
lb|13974,13976
)|13976,13977
.|13978,13979
Please|13980,13986
<EOL>|13987,13988
weigh|13988,13993
yourself|13994,14002
today|14003,14008
at|14009,14011
home|14012,14016
and|14017,14020
use|14021,14024
this|14025,14029
as|14030,14032
your|14033,14037
new|14038,14041
baseline|14042,14050
<EOL>|14052,14053
-|14054,14055
Please|14055,14061
weigh|14062,14067
yourself|14068,14076
every|14077,14082
day|14083,14086
in|14087,14089
the|14090,14093
morning|14094,14101
.|14101,14102
Call|14103,14107
your|14108,14112
<EOL>|14113,14114
doctor|14114,14120
if|14121,14123
your|14124,14128
weight|14129,14135
goes|14136,14140
up|14141,14143
by|14144,14146
more|14147,14151
than|14152,14156
3|14157,14158
lbs|14159,14162
.|14162,14163
<EOL>|14165,14166
-|14167,14168
Seek|14169,14173
medical|14174,14181
attention|14182,14191
if|14192,14194
you|14195,14198
have|14199,14203
new|14204,14207
or|14208,14210
concerning|14211,14221
symptoms|14222,14230
<EOL>|14231,14232
or|14232,14234
you|14235,14238
develop|14239,14246
swelling|14247,14255
in|14256,14258
your|14259,14263
legs|14264,14268
,|14268,14269
abdominal|14270,14279
distention|14280,14290
,|14290,14291
or|14292,14294
<EOL>|14295,14296
shortness|14296,14305
of|14306,14308
breath|14309,14315
.|14315,14316
If|14317,14319
you|14320,14323
have|14324,14328
worsening|14329,14338
pain|14339,14343
or|14344,14346
redness|14347,14354
in|14355,14357
<EOL>|14358,14359
your|14359,14363
foot|14364,14368
,|14368,14369
urinating|14370,14379
frequently|14380,14390
or|14391,14393
very|14394,14398
thirsty|14399,14406
,|14406,14407
or|14408,14410
if|14411,14413
your|14414,14418
<EOL>|14419,14420
blood|14420,14425
sugar|14426,14431
is|14432,14434
consistently|14435,14447
above|14448,14453
300|14454,14457
or|14458,14460
below|14461,14466
70|14467,14469
please|14470,14476
cal|14477,14480
<EOL>|14481,14482
your|14482,14486
doctor|14487,14493
.|14493,14494
<EOL>|14495,14496
<EOL>|14497,14498
It|14498,14500
was|14501,14504
a|14505,14506
pleasure|14507,14515
participating|14516,14529
in|14530,14532
your|14533,14537
care|14538,14542
.|14542,14543
We|14544,14546
wish|14547,14551
you|14552,14555
the|14556,14559
<EOL>|14560,14561
_|14561,14562
_|14562,14563
_|14563,14564
!|14564,14565
<EOL>|14567,14568
-|14569,14570
Your|14570,14574
_|14575,14576
_|14576,14577
_|14577,14578
Care|14579,14583
Team|14584,14588
<EOL>|14590,14591
<EOL>|14592,14593
<EOL>|14594,14595
Followup|14595,14603
Instructions|14604,14616
:|14616,14617
<EOL>|14617,14618
_|14618,14619
_|14619,14620
_|14620,14621
<EOL>|14621,14622

