 Token Text | Text Span 
<EOL>|1,2
Name|2,6
:|6,7
_|9,10
_|10,11
_|11,12
Unit|29,33
No|34,36
:|36,37
_|40,41
_|41,42
_|42,43
<EOL>|43,44
<EOL>|45,46
Admission|46,55
Date|56,60
:|60,61
_|63,64
_|64,65
_|65,66
Discharge|80,89
Date|90,94
:|94,95
_|98,99
_|99,100
_|100,101
<EOL>|101,102
<EOL>|103,104
Date|104,108
of|109,111
Birth|112,117
:|117,118
_|120,121
_|121,122
_|122,123
Sex|136,139
:|139,140
F|143,144
<EOL>|144,145
<EOL>|146,147
Service|147,154
:|154,155
SURGERY|156,163
<EOL>|163,164
<EOL>|165,166
_|178,179
_|179,180
_|180,181
<EOL>|181,182
<EOL>|183,184
Attending|184,193
:|193,194
_|195,196
_|196,197
_|197,198
.|198,199
<EOL>|199,200
<EOL>|201,202
Nausea|219,225
/|225,226
Vomiting|226,234
<EOL>|234,235
<EOL>|236,237
Major|237,242
Surgical|243,251
or|252,254
Invasive|255,263
Procedure|264,273
:|273,274
<EOL>|274,275
Band|275,279
adjustment|280,290
<EOL>|290,291
<EOL>|291,292
<EOL>|293,294
Ms.|322,325
_|326,327
_|327,328
_|328,329
is|330,332
a|333,334
_|335,336
_|336,337
_|337,338
s|339,340
/|340,341
p|341,342
lap|343,346
band|347,351
in|352,354
_|355,356
_|356,357
_|357,358
who|359,362
prsents|363,370
with|371,375
a|376,377
1|378,379
<EOL>|379,380
week|380,384
history|385,392
of|393,395
nausea|396,402
,|402,403
non-bilious|404,415
non-bloody|416,426
emesis|427,433
of|434,436
<EOL>|436,437
undigested|437,447
food|448,452
after|453,458
eating|459,465
,|465,466
intolerance|467,478
to|479,481
solids|482,488
/|488,489
softs|489,494
,|494,495
<EOL>|495,496
hypersalivation|496,511
,|511,512
and|513,516
moderate|517,525
post-prandial|526,539
epigastric|540,550
<EOL>|550,551
discomfort|551,561
.|561,562
She|563,566
denies|567,573
fever|574,579
,|579,580
chills|581,587
,|587,588
hematemesis|589,600
,|600,601
BRBPR|602,607
,|607,608
<EOL>|609,610
melena|610,616
,|616,617
<EOL>|617,618
diarrhea|618,626
,|626,627
or|628,630
sympotoms|631,640
of|641,643
dehydration|644,655
,|655,656
but|657,660
was|661,664
recently|665,673
<EOL>|674,675
evaluated|675,684
<EOL>|684,685
for|685,688
dizziness|689,698
in|699,701
an|702,704
ED|705,707
with|708,712
a|713,714
diagnosis|715,724
given|725,730
of|731,733
BPPV|734,738
.|738,739
Of|740,742
note|743,747
,|747,748
<EOL>|748,749
the|749,752
patient|753,760
underwent|761,770
an|771,773
unfill|774,780
of|781,783
her|784,787
band|788,792
from|793,797
5.8|798,801
to|802,804
3.8|805,808
ml|808,810
on|811,813
<EOL>|813,814
_|814,815
_|815,816
_|816,817
for|818,821
similar|822,829
symptoms|830,838
,|838,839
the|840,843
band|844,848
was|849,852
subseqently|853,864
been|865,869
filled|870,876
<EOL>|876,877
to|877,879
4.8|880,883
on|884,886
_|887,888
_|888,889
_|889,890
,|890,891
5.2|892,895
on|896,898
_|899,900
_|900,901
_|901,902
,|902,903
and|904,907
most|908,912
recently|913,921
to|922,924
5.6|925,928
ml|928,930
on|931,933
<EOL>|934,935
_|935,936
_|936,937
_|937,938
.|938,939
<EOL>|939,940
<EOL>|940,941
<EOL>|942,943
PMHx|965,969
:|969,970
Hyperlipidemia|971,985
and|986,989
with|990,994
elevated|995,1003
triglyceride|1004,1016
,|1016,1017
iron|1018,1022
<EOL>|1022,1023
deficiency|1023,1033
anemia|1034,1040
,|1040,1041
irritable|1042,1051
bowel|1052,1057
syndrome|1058,1066
,|1066,1067
allergic|1068,1076
rhinitis|1077,1085
,|1085,1086
<EOL>|1086,1087
dysmenorrhea|1087,1099
,|1099,1100
vitamin|1101,1108
D|1109,1110
deficiency|1111,1121
,|1121,1122
question|1123,1131
of|1132,1134
hypothyroidism|1135,1149
<EOL>|1149,1150
with|1150,1154
elevated|1155,1163
TSH|1164,1167
level|1168,1173
,|1173,1174
thalassemia|1175,1186
trait|1187,1192
,|1192,1193
fatty|1194,1199
liver|1200,1205
and|1206,1209
<EOL>|1209,1210
cholelithiasis|1210,1224
by|1225,1227
ultrasound|1228,1238
study|1239,1244
.|1244,1245
A|1246,1247
history|1248,1255
of|1256,1258
kissing|1259,1266
tonsils|1267,1274
<EOL>|1274,1275
that|1275,1279
was|1280,1283
associated|1284,1294
with|1295,1299
obstructive|1300,1311
sleep|1312,1317
apnea|1318,1323
and|1324,1327
<EOL>|1327,1328
gastroesophageal|1328,1344
reflux|1345,1351
,|1351,1352
these|1353,1358
have|1359,1363
resolved|1364,1372
completely|1373,1383
after|1384,1389
<EOL>|1390,1391
the|1391,1394
<EOL>|1394,1395
tonsillectomy|1395,1408
in|1409,1411
_|1412,1413
_|1413,1414
_|1414,1415
.|1415,1416
History|1417,1424
of|1425,1427
polycystic|1428,1438
ovary|1439,1444
<EOL>|1444,1445
syndrome|1445,1453
<EOL>|1453,1454
<EOL>|1455,1456
:|1470,1471
<EOL>|1471,1472
_|1472,1473
_|1473,1474
_|1474,1475
<EOL>|1475,1476
:|1490,1491
<EOL>|1491,1492
bladder|1492,1499
CA|1500,1502
;|1502,1503
with|1504,1508
diabetes|1509,1517
,|1517,1518
breast|1519,1525
neoplasia|1526,1535
,|1535,1536
colon|1537,1542
CA|1543,1545
,|1545,1546
ovarian|1547,1554
<EOL>|1555,1556
CA|1556,1558
and|1559,1562
sarcoma|1563,1570
<EOL>|1570,1571
<EOL>|1572,1573
VS|1588,1590
:|1590,1591
Temp|1592,1596
:|1596,1597
97.9|1598,1602
,|1602,1603
HR|1604,1606
:|1606,1607
72|1608,1610
,|1610,1611
BP|1612,1614
:|1614,1615
113|1616,1619
/|1619,1620
64|1620,1622
,|1622,1623
RR|1624,1626
:|1626,1627
16|1628,1630
,|1630,1631
O2sat|1632,1637
:|1637,1638
100|1639,1642
%|1642,1643
RA|1644,1646
<EOL>|1647,1648
GEN|1648,1651
:|1651,1652
A|1653,1654
&|1654,1655
O|1655,1656
,|1656,1657
NAD|1658,1661
<EOL>|1661,1662
HEENT|1662,1667
:|1667,1668
No|1669,1671
scleral|1672,1679
icterus|1680,1687
,|1687,1688
MMM|1689,1692
<EOL>|1692,1693
CV|1693,1695
:|1695,1696
RRR|1697,1700
<EOL>|1700,1701
PULM|1701,1705
:|1705,1706
No|1707,1709
W|1710,1711
/|1711,1712
R|1712,1713
/|1713,1714
C|1714,1715
,|1715,1716
no|1717,1719
increased|1720,1729
work|1730,1734
of|1735,1737
breathing|1738,1747
<EOL>|1747,1748
ABD|1748,1751
:|1751,1752
Soft|1753,1757
,|1757,1758
nondistended|1759,1771
,|1771,1772
non-tender|1773,1783
to|1784,1786
palpation|1787,1796
in|1797,1799
epigastric|1800,1810
<EOL>|1811,1812
region|1812,1818
,|1818,1819
no|1820,1822
rebound|1823,1830
or|1831,1833
guarding|1834,1842
,|1842,1843
palpable|1844,1852
port|1853,1857
<EOL>|1857,1858
Ext|1858,1861
:|1861,1862
No|1863,1865
_|1866,1867
_|1867,1868
_|1868,1869
edema|1870,1875
,|1875,1876
warm|1877,1881
and|1882,1885
well|1886,1890
perfused|1891,1899
<EOL>|1899,1900
<EOL>|1900,1901
<EOL>|1902,1903
Pertinent|1903,1912
Results|1913,1920
:|1920,1921
<EOL>|1921,1922
_|1922,1923
_|1923,1924
_|1924,1925
12|1926,1928
:|1928,1929
16AM|1929,1933
PLT|1936,1939
COUNT|1940,1945
-|1945,1946
243|1946,1949
<EOL>|1949,1950
_|1950,1951
_|1951,1952
_|1952,1953
12|1954,1956
:|1956,1957
16AM|1957,1961
NEUTS|1964,1969
-|1969,1970
46.0|1970,1974
_|1975,1976
_|1976,1977
_|1977,1978
MONOS|1979,1984
-|1984,1985
6.9|1985,1988
EOS|1989,1992
-|1992,1993
1.8|1993,1996
<EOL>|1997,1998
BASOS|1998,2003
-|2003,2004
0.5|2004,2007
IM|2008,2010
_|2011,2012
_|2012,2013
_|2013,2014
AbsNeut|2015,2022
-|2022,2023
4|2023,2024
.|2024,2025
88|2025,2027
AbsLymp|2028,2035
-|2035,2036
4|2036,2037
.|2037,2038
72|2038,2040
*|2040,2041
AbsMono|2042,2049
-|2049,2050
0|2050,2051
.|2051,2052
73|2052,2054
<EOL>|2055,2056
AbsEos|2056,2062
-|2062,2063
0|2063,2064
.|2064,2065
19|2065,2067
AbsBaso|2068,2075
-|2075,2076
0|2076,2077
.|2077,2078
05|2078,2080
<EOL>|2080,2081
_|2081,2082
_|2082,2083
_|2083,2084
12|2085,2087
:|2087,2088
16AM|2088,2092
estGFR|2095,2101
-|2101,2102
Using|2102,2107
this|2108,2112
<EOL>|2112,2113
_|2113,2114
_|2114,2115
_|2115,2116
01|2117,2119
:|2119,2120
02AM|2120,2124
URINE|2125,2130
MUCOUS|2132,2138
-|2138,2139
RARE|2139,2143
<EOL>|2143,2144
_|2144,2145
_|2145,2146
_|2146,2147
01|2148,2150
:|2150,2151
02AM|2151,2155
URINE|2156,2161
HYALINE|2163,2170
-|2170,2171
1|2171,2172
*|2172,2173
<EOL>|2173,2174
_|2174,2175
_|2175,2176
_|2176,2177
01|2178,2180
:|2180,2181
02AM|2181,2185
URINE|2186,2191
RBC|2193,2196
-|2196,2197
4|2197,2198
*|2198,2199
WBC|2200,2203
-|2203,2204
4|2204,2205
BACTERIA|2206,2214
-|2214,2215
MOD|2215,2218
YEAST|2219,2224
-|2224,2225
NONE|2225,2229
<EOL>|2230,2231
EPI|2231,2234
-|2234,2235
11|2235,2237
<EOL>|2237,2238
_|2238,2239
_|2239,2240
_|2240,2241
01|2242,2244
:|2244,2245
02AM|2245,2249
URINE|2250,2255
BLOOD|2257,2262
-|2262,2263
NEG|2263,2266
NITRITE|2267,2274
-|2274,2275
NEG|2275,2278
PROTEIN|2279,2286
-|2286,2287
30|2287,2289
<EOL>|2290,2291
GLUCOSE|2291,2298
-|2298,2299
NEG|2299,2302
KETONE|2303,2309
-|2309,2310
NEG|2310,2313
BILIRUBIN|2314,2323
-|2323,2324
NEG|2324,2327
UROBILNGN|2328,2337
-|2337,2338
NEG|2338,2341
PH|2342,2344
-|2344,2345
6.5|2345,2348
<EOL>|2349,2350
LEUK|2350,2354
-|2354,2355
TR|2355,2357
<EOL>|2357,2358
_|2358,2359
_|2359,2360
_|2360,2361
01|2362,2364
:|2364,2365
02AM|2365,2369
URINE|2370,2375
COLOR|2377,2382
-|2382,2383
Yellow|2383,2389
APPEAR|2390,2396
-|2396,2397
Hazy|2397,2401
SP|2402,2404
_|2405,2406
_|2406,2407
_|2407,2408
<EOL>|2408,2409
_|2409,2410
_|2410,2411
_|2411,2412
01|2413,2415
:|2415,2416
02AM|2416,2420
URINE|2421,2426
UCG|2428,2431
-|2431,2432
NEGATIVE|2432,2440
<EOL>|2440,2441
_|2441,2442
_|2442,2443
_|2443,2444
01|2445,2447
:|2447,2448
02AM|2448,2452
URINE|2453,2458
HOURS|2460,2465
-|2465,2466
RANDOM|2466,2472
<EOL>|2472,2473
_|2473,2474
_|2474,2475
_|2475,2476
01|2477,2479
:|2479,2480
02AM|2480,2484
URINE|2485,2490
HOURS|2492,2497
-|2497,2498
RANDOM|2498,2504
<EOL>|2504,2505
<EOL>|2506,2507
_|2530,2531
_|2531,2532
_|2532,2533
was|2534,2537
admitted|2538,2546
from|2547,2551
ED|2552,2554
on|2555,2557
_|2558,2559
_|2559,2560
_|2560,2561
for|2562,2565
nausea|2566,2572
and|2573,2576
<EOL>|2577,2578
vomiting|2578,2586
after|2587,2592
any|2593,2596
po|2597,2599
intake|2600,2606
.|2606,2607
Of|2608,2610
note|2611,2615
,|2615,2616
she|2617,2620
has|2621,2624
had|2625,2628
similar|2629,2636
<EOL>|2637,2638
symptomes|2638,2647
last|2648,2652
year|2653,2657
.|2657,2658
She|2659,2662
was|2663,2666
started|2667,2674
on|2675,2677
IV|2678,2680
fluids|2681,2687
for|2688,2691
<EOL>|2692,2693
rehydration|2693,2704
.|2704,2705
Her|2706,2709
laboratory|2710,2720
values|2721,2727
were|2728,2732
unremarkable|2733,2745
on|2746,2748
<EOL>|2749,2750
admission|2750,2759
and|2760,2763
her|2764,2767
symptoms|2768,2776
gradually|2777,2786
improved|2787,2795
with|2796,2800
anti-emetic|2801,2812
<EOL>|2813,2814
medications|2814,2825
and|2826,2829
IV|2830,2832
fluid|2833,2838
therapy|2839,2846
.|2846,2847
She|2848,2851
was|2852,2855
back|2856,2860
to|2861,2863
her|2864,2867
baseline|2868,2876
<EOL>|2877,2878
clinical|2878,2886
status|2887,2893
after|2894,2899
unfilling|2900,2909
the|2910,2913
band|2914,2918
by|2919,2921
1.5|2922,2925
cc|2925,2927
.|2927,2928
Water|2929,2934
<EOL>|2935,2936
challenge|2936,2945
test|2946,2950
was|2951,2954
done|2955,2959
after|2960,2965
band|2966,2970
adjustment|2971,2981
and|2982,2985
was|2986,2989
negative|2990,2998
<EOL>|2999,3000
for|3000,3003
any|3004,3007
pain|3008,3012
,|3012,3013
nausea|3014,3020
or|3021,3023
vomiting|3024,3032
.|3032,3033
She|3034,3037
was|3038,3041
discharged|3042,3052
in|3053,3055
good|3056,3060
<EOL>|3061,3062
condition|3062,3071
with|3072,3076
instructions|3077,3089
to|3090,3092
follow|3093,3099
up|3100,3102
with|3103,3107
Dr.|3108,3111
_|3112,3113
_|3113,3114
_|3114,3115
<EOL>|3116,3117
_|3117,3118
_|3118,3119
_|3119,3120
after|3121,3126
2|3127,3128
.|3128,3129
<EOL>|3130,3131
<EOL>|3131,3132
<EOL>|3133,3134
Discharge|3134,3143
Medications|3144,3155
:|3155,3156
<EOL>|3156,3157
1.|3157,3159
Lorazepam|3160,3169
0.5|3170,3173
mg|3174,3176
PO|3177,3179
BID|3180,3183
:|3183,3184
PRN|3184,3187
anxiety|3188,3195
<EOL>|3196,3197
2.|3197,3199
BusPIRone|3200,3209
5|3210,3211
mg|3212,3214
PO|3215,3217
TID|3218,3221
<EOL>|3222,3223
<EOL>|3223,3224
<EOL>|3225,3226
Discharge|3226,3235
Disposition|3236,3247
:|3247,3248
<EOL>|3248,3249
Home|3249,3253
<EOL>|3253,3254
<EOL>|3255,3256
Discharge|3256,3265
Diagnosis|3266,3275
:|3275,3276
<EOL>|3276,3277
nausea|3277,3283
and|3284,3287
vomiting|3288,3296
due|3297,3300
to|3301,3303
tight|3304,3309
band|3310,3314
<EOL>|3314,3315
<EOL>|3315,3316
<EOL>|3317,3318
Mental|3339,3345
Status|3346,3352
:|3352,3353
Clear|3354,3359
and|3360,3363
coherent|3364,3372
.|3372,3373
<EOL>|3373,3374
Level|3374,3379
of|3380,3382
Consciousness|3383,3396
:|3396,3397
Alert|3398,3403
and|3404,3407
interactive|3408,3419
.|3419,3420
<EOL>|3420,3421
Activity|3421,3429
Status|3430,3436
:|3436,3437
Ambulatory|3438,3448
-|3449,3450
Independent|3451,3462
.|3462,3463
<EOL>|3463,3464
<EOL>|3464,3465
<EOL>|3466,3467
You|3491,3494
were|3495,3499
admitted|3500,3508
to|3509,3511
_|3512,3513
_|3513,3514
_|3514,3515
for|3516,3519
your|3520,3524
Nausea|3525,3531
and|3532,3535
vomiting|3536,3544
.|3544,3545
Your|3546,3550
<EOL>|3551,3552
band|3552,3556
was|3557,3560
tight|3561,3566
enough|3567,3573
to|3574,3576
cause|3577,3582
your|3583,3587
nausea|3588,3594
and|3595,3598
vomiting|3599,3607
,|3607,3608
1.5|3609,3612
cc|3613,3615
<EOL>|3616,3617
has|3617,3620
been|3621,3625
taken|3626,3631
out|3632,3635
from|3636,3640
your|3641,3645
band|3646,3650
in|3651,3653
which|3654,3659
2.5|3660,3663
cc|3663,3665
total|3666,3671
left|3672,3676
.|3676,3677
you|3678,3681
<EOL>|3682,3683
subsequently|3683,3695
tolerated|3696,3705
a|3706,3707
water|3708,3713
bolus|3714,3719
test|3720,3724
.|3724,3725
You|3726,3729
have|3730,3734
been|3735,3739
deemed|3740,3746
<EOL>|3747,3748
fit|3748,3751
to|3752,3754
be|3755,3757
discharged|3758,3768
from|3769,3773
the|3774,3777
hospital|3778,3786
.|3786,3787
Please|3788,3794
return|3795,3801
if|3802,3804
your|3805,3809
<EOL>|3810,3811
nausea|3811,3817
becomes|3818,3825
untolerable|3826,3837
or|3838,3840
you|3841,3844
start|3845,3850
vomiting|3851,3859
again|3860,3865
.|3865,3866
Please|3867,3873
<EOL>|3874,3875
continue|3875,3883
taking|3884,3890
your|3891,3895
home|3896,3900
medications|3901,3912
.|3912,3913
<EOL>|3913,3914
Thank|3914,3919
you|3920,3923
for|3924,3927
letting|3928,3935
us|3936,3938
participate|3939,3950
in|3951,3953
your|3954,3958
healthcare|3959,3969
.|3969,3970
<EOL>|3971,3972
<EOL>|3972,3973
<EOL>|3974,3975
Followup|3975,3983
Instructions|3984,3996
:|3996,3997
<EOL>|3997,3998
_|3998,3999
_|3999,4000
_|4000,4001
<EOL>|4001,4002

